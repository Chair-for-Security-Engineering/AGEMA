
module AES ( plaintext, key, reset, clk, ciphertext, done );
  (* AGEMA = "secure" *) input [127:0] plaintext;
  (* AGEMA = "secure" *) input [127:0] key;
  (* AGEMA = "clock" *)  input clk;
  (* AGEMA = "reset" *)  input reset;

  output [127:0] ciphertext;
  output done;

  wire   n283, n285, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, RoundReg_Inst_ff_SDE_0_next_state,
         RoundReg_Inst_ff_SDE_0_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_1_next_state,
         RoundReg_Inst_ff_SDE_1_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_2_next_state,
         RoundReg_Inst_ff_SDE_2_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_3_next_state,
         RoundReg_Inst_ff_SDE_3_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_4_next_state,
         RoundReg_Inst_ff_SDE_4_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_5_next_state,
         RoundReg_Inst_ff_SDE_5_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_6_next_state,
         RoundReg_Inst_ff_SDE_6_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_7_next_state,
         RoundReg_Inst_ff_SDE_7_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_8_next_state,
         RoundReg_Inst_ff_SDE_8_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_9_next_state,
         RoundReg_Inst_ff_SDE_9_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_10_next_state,
         RoundReg_Inst_ff_SDE_10_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_11_next_state,
         RoundReg_Inst_ff_SDE_11_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_12_next_state,
         RoundReg_Inst_ff_SDE_12_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_13_next_state,
         RoundReg_Inst_ff_SDE_13_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_14_next_state,
         RoundReg_Inst_ff_SDE_14_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_15_next_state,
         RoundReg_Inst_ff_SDE_15_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_16_next_state,
         RoundReg_Inst_ff_SDE_16_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_17_next_state,
         RoundReg_Inst_ff_SDE_17_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_18_next_state,
         RoundReg_Inst_ff_SDE_18_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_19_next_state,
         RoundReg_Inst_ff_SDE_19_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_20_next_state,
         RoundReg_Inst_ff_SDE_20_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_21_next_state,
         RoundReg_Inst_ff_SDE_21_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_22_next_state,
         RoundReg_Inst_ff_SDE_22_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_23_next_state,
         RoundReg_Inst_ff_SDE_23_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_24_next_state,
         RoundReg_Inst_ff_SDE_24_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_25_next_state,
         RoundReg_Inst_ff_SDE_25_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_26_next_state,
         RoundReg_Inst_ff_SDE_26_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_27_next_state,
         RoundReg_Inst_ff_SDE_27_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_28_next_state,
         RoundReg_Inst_ff_SDE_28_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_29_next_state,
         RoundReg_Inst_ff_SDE_29_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_30_next_state,
         RoundReg_Inst_ff_SDE_30_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_31_next_state,
         RoundReg_Inst_ff_SDE_31_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_32_next_state,
         RoundReg_Inst_ff_SDE_32_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_33_next_state,
         RoundReg_Inst_ff_SDE_33_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_34_next_state,
         RoundReg_Inst_ff_SDE_34_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_35_next_state,
         RoundReg_Inst_ff_SDE_35_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_36_next_state,
         RoundReg_Inst_ff_SDE_36_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_37_next_state,
         RoundReg_Inst_ff_SDE_37_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_38_next_state,
         RoundReg_Inst_ff_SDE_38_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_39_next_state,
         RoundReg_Inst_ff_SDE_39_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_40_next_state,
         RoundReg_Inst_ff_SDE_40_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_41_next_state,
         RoundReg_Inst_ff_SDE_41_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_42_next_state,
         RoundReg_Inst_ff_SDE_42_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_43_next_state,
         RoundReg_Inst_ff_SDE_43_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_44_next_state,
         RoundReg_Inst_ff_SDE_44_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_45_next_state,
         RoundReg_Inst_ff_SDE_45_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_46_next_state,
         RoundReg_Inst_ff_SDE_46_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_47_next_state,
         RoundReg_Inst_ff_SDE_47_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_48_next_state,
         RoundReg_Inst_ff_SDE_48_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_49_next_state,
         RoundReg_Inst_ff_SDE_49_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_50_next_state,
         RoundReg_Inst_ff_SDE_50_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_51_next_state,
         RoundReg_Inst_ff_SDE_51_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_52_next_state,
         RoundReg_Inst_ff_SDE_52_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_53_next_state,
         RoundReg_Inst_ff_SDE_53_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_54_next_state,
         RoundReg_Inst_ff_SDE_54_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_55_next_state,
         RoundReg_Inst_ff_SDE_55_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_56_next_state,
         RoundReg_Inst_ff_SDE_56_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_57_next_state,
         RoundReg_Inst_ff_SDE_57_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_58_next_state,
         RoundReg_Inst_ff_SDE_58_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_59_next_state,
         RoundReg_Inst_ff_SDE_59_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_60_next_state,
         RoundReg_Inst_ff_SDE_60_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_61_next_state,
         RoundReg_Inst_ff_SDE_61_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_62_next_state,
         RoundReg_Inst_ff_SDE_62_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_63_next_state,
         RoundReg_Inst_ff_SDE_63_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_64_next_state,
         RoundReg_Inst_ff_SDE_64_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_65_next_state,
         RoundReg_Inst_ff_SDE_65_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_66_next_state,
         RoundReg_Inst_ff_SDE_66_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_67_next_state,
         RoundReg_Inst_ff_SDE_67_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_68_next_state,
         RoundReg_Inst_ff_SDE_68_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_69_next_state,
         RoundReg_Inst_ff_SDE_69_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_70_next_state,
         RoundReg_Inst_ff_SDE_70_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_71_next_state,
         RoundReg_Inst_ff_SDE_71_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_72_next_state,
         RoundReg_Inst_ff_SDE_72_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_73_next_state,
         RoundReg_Inst_ff_SDE_73_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_74_next_state,
         RoundReg_Inst_ff_SDE_74_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_75_next_state,
         RoundReg_Inst_ff_SDE_75_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_76_next_state,
         RoundReg_Inst_ff_SDE_76_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_77_next_state,
         RoundReg_Inst_ff_SDE_77_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_78_next_state,
         RoundReg_Inst_ff_SDE_78_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_79_next_state,
         RoundReg_Inst_ff_SDE_79_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_80_next_state,
         RoundReg_Inst_ff_SDE_80_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_81_next_state,
         RoundReg_Inst_ff_SDE_81_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_82_next_state,
         RoundReg_Inst_ff_SDE_82_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_83_next_state,
         RoundReg_Inst_ff_SDE_83_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_84_next_state,
         RoundReg_Inst_ff_SDE_84_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_85_next_state,
         RoundReg_Inst_ff_SDE_85_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_86_next_state,
         RoundReg_Inst_ff_SDE_86_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_87_next_state,
         RoundReg_Inst_ff_SDE_87_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_88_next_state,
         RoundReg_Inst_ff_SDE_88_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_89_next_state,
         RoundReg_Inst_ff_SDE_89_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_90_next_state,
         RoundReg_Inst_ff_SDE_90_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_91_next_state,
         RoundReg_Inst_ff_SDE_91_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_92_next_state,
         RoundReg_Inst_ff_SDE_92_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_93_next_state,
         RoundReg_Inst_ff_SDE_93_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_94_next_state,
         RoundReg_Inst_ff_SDE_94_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_95_next_state,
         RoundReg_Inst_ff_SDE_95_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_96_next_state,
         RoundReg_Inst_ff_SDE_96_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_97_next_state,
         RoundReg_Inst_ff_SDE_97_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_98_next_state,
         RoundReg_Inst_ff_SDE_98_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_99_next_state,
         RoundReg_Inst_ff_SDE_99_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_100_next_state,
         RoundReg_Inst_ff_SDE_100_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_101_next_state,
         RoundReg_Inst_ff_SDE_101_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_102_next_state,
         RoundReg_Inst_ff_SDE_102_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_103_next_state,
         RoundReg_Inst_ff_SDE_103_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_104_next_state,
         RoundReg_Inst_ff_SDE_104_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_105_next_state,
         RoundReg_Inst_ff_SDE_105_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_106_next_state,
         RoundReg_Inst_ff_SDE_106_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_107_next_state,
         RoundReg_Inst_ff_SDE_107_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_108_next_state,
         RoundReg_Inst_ff_SDE_108_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_109_next_state,
         RoundReg_Inst_ff_SDE_109_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_110_next_state,
         RoundReg_Inst_ff_SDE_110_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_111_next_state,
         RoundReg_Inst_ff_SDE_111_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_112_next_state,
         RoundReg_Inst_ff_SDE_112_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_113_next_state,
         RoundReg_Inst_ff_SDE_113_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_114_next_state,
         RoundReg_Inst_ff_SDE_114_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_115_next_state,
         RoundReg_Inst_ff_SDE_115_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_116_next_state,
         RoundReg_Inst_ff_SDE_116_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_117_next_state,
         RoundReg_Inst_ff_SDE_117_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_118_next_state,
         RoundReg_Inst_ff_SDE_118_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_119_next_state,
         RoundReg_Inst_ff_SDE_119_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_120_next_state,
         RoundReg_Inst_ff_SDE_120_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_121_next_state,
         RoundReg_Inst_ff_SDE_121_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_122_next_state,
         RoundReg_Inst_ff_SDE_122_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_123_next_state,
         RoundReg_Inst_ff_SDE_123_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_124_next_state,
         RoundReg_Inst_ff_SDE_124_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_125_next_state,
         RoundReg_Inst_ff_SDE_125_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_126_next_state,
         RoundReg_Inst_ff_SDE_126_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_127_next_state,
         RoundReg_Inst_ff_SDE_127_current_state_reg_QN,
         SubBytesIns_Inst_Sbox_0_L29, SubBytesIns_Inst_Sbox_0_L28,
         SubBytesIns_Inst_Sbox_0_L27, SubBytesIns_Inst_Sbox_0_L26,
         SubBytesIns_Inst_Sbox_0_L25, SubBytesIns_Inst_Sbox_0_L24,
         SubBytesIns_Inst_Sbox_0_L23, SubBytesIns_Inst_Sbox_0_L22,
         SubBytesIns_Inst_Sbox_0_L21, SubBytesIns_Inst_Sbox_0_L20,
         SubBytesIns_Inst_Sbox_0_L19, SubBytesIns_Inst_Sbox_0_L18,
         SubBytesIns_Inst_Sbox_0_L17, SubBytesIns_Inst_Sbox_0_L16,
         SubBytesIns_Inst_Sbox_0_L15, SubBytesIns_Inst_Sbox_0_L14,
         SubBytesIns_Inst_Sbox_0_L13, SubBytesIns_Inst_Sbox_0_L12,
         SubBytesIns_Inst_Sbox_0_L11, SubBytesIns_Inst_Sbox_0_L10,
         SubBytesIns_Inst_Sbox_0_L9, SubBytesIns_Inst_Sbox_0_L8,
         SubBytesIns_Inst_Sbox_0_L7, SubBytesIns_Inst_Sbox_0_L6,
         SubBytesIns_Inst_Sbox_0_L5, SubBytesIns_Inst_Sbox_0_L4,
         SubBytesIns_Inst_Sbox_0_L3, SubBytesIns_Inst_Sbox_0_L2,
         SubBytesIns_Inst_Sbox_0_L1, SubBytesIns_Inst_Sbox_0_L0,
         SubBytesIns_Inst_Sbox_0_M63, SubBytesIns_Inst_Sbox_0_M62,
         SubBytesIns_Inst_Sbox_0_M61, SubBytesIns_Inst_Sbox_0_M60,
         SubBytesIns_Inst_Sbox_0_M59, SubBytesIns_Inst_Sbox_0_M58,
         SubBytesIns_Inst_Sbox_0_M57, SubBytesIns_Inst_Sbox_0_M56,
         SubBytesIns_Inst_Sbox_0_M55, SubBytesIns_Inst_Sbox_0_M54,
         SubBytesIns_Inst_Sbox_0_M53, SubBytesIns_Inst_Sbox_0_M52,
         SubBytesIns_Inst_Sbox_0_M51, SubBytesIns_Inst_Sbox_0_M50,
         SubBytesIns_Inst_Sbox_0_M49, SubBytesIns_Inst_Sbox_0_M48,
         SubBytesIns_Inst_Sbox_0_M47, SubBytesIns_Inst_Sbox_0_M46,
         SubBytesIns_Inst_Sbox_0_M45, SubBytesIns_Inst_Sbox_0_M44,
         SubBytesIns_Inst_Sbox_0_M43, SubBytesIns_Inst_Sbox_0_M42,
         SubBytesIns_Inst_Sbox_0_M41, SubBytesIns_Inst_Sbox_0_M40,
         SubBytesIns_Inst_Sbox_0_M39, SubBytesIns_Inst_Sbox_0_M38,
         SubBytesIns_Inst_Sbox_0_M37, SubBytesIns_Inst_Sbox_0_M36,
         SubBytesIns_Inst_Sbox_0_M35, SubBytesIns_Inst_Sbox_0_M34,
         SubBytesIns_Inst_Sbox_0_M33, SubBytesIns_Inst_Sbox_0_M32,
         SubBytesIns_Inst_Sbox_0_M31, SubBytesIns_Inst_Sbox_0_M30,
         SubBytesIns_Inst_Sbox_0_M29, SubBytesIns_Inst_Sbox_0_M28,
         SubBytesIns_Inst_Sbox_0_M27, SubBytesIns_Inst_Sbox_0_M26,
         SubBytesIns_Inst_Sbox_0_M25, SubBytesIns_Inst_Sbox_0_M24,
         SubBytesIns_Inst_Sbox_0_M23, SubBytesIns_Inst_Sbox_0_M22,
         SubBytesIns_Inst_Sbox_0_M21, SubBytesIns_Inst_Sbox_0_M20,
         SubBytesIns_Inst_Sbox_0_M19, SubBytesIns_Inst_Sbox_0_M18,
         SubBytesIns_Inst_Sbox_0_M17, SubBytesIns_Inst_Sbox_0_M16,
         SubBytesIns_Inst_Sbox_0_M15, SubBytesIns_Inst_Sbox_0_M14,
         SubBytesIns_Inst_Sbox_0_M13, SubBytesIns_Inst_Sbox_0_M12,
         SubBytesIns_Inst_Sbox_0_M11, SubBytesIns_Inst_Sbox_0_M10,
         SubBytesIns_Inst_Sbox_0_M9, SubBytesIns_Inst_Sbox_0_M8,
         SubBytesIns_Inst_Sbox_0_M7, SubBytesIns_Inst_Sbox_0_M6,
         SubBytesIns_Inst_Sbox_0_M5, SubBytesIns_Inst_Sbox_0_M4,
         SubBytesIns_Inst_Sbox_0_M3, SubBytesIns_Inst_Sbox_0_M2,
         SubBytesIns_Inst_Sbox_0_M1, SubBytesIns_Inst_Sbox_0_T27,
         SubBytesIns_Inst_Sbox_0_T26, SubBytesIns_Inst_Sbox_0_T25,
         SubBytesIns_Inst_Sbox_0_T24, SubBytesIns_Inst_Sbox_0_T23,
         SubBytesIns_Inst_Sbox_0_T22, SubBytesIns_Inst_Sbox_0_T21,
         SubBytesIns_Inst_Sbox_0_T20, SubBytesIns_Inst_Sbox_0_T19,
         SubBytesIns_Inst_Sbox_0_T18, SubBytesIns_Inst_Sbox_0_T17,
         SubBytesIns_Inst_Sbox_0_T16, SubBytesIns_Inst_Sbox_0_T15,
         SubBytesIns_Inst_Sbox_0_T14, SubBytesIns_Inst_Sbox_0_T13,
         SubBytesIns_Inst_Sbox_0_T12, SubBytesIns_Inst_Sbox_0_T11,
         SubBytesIns_Inst_Sbox_0_T10, SubBytesIns_Inst_Sbox_0_T9,
         SubBytesIns_Inst_Sbox_0_T8, SubBytesIns_Inst_Sbox_0_T7,
         SubBytesIns_Inst_Sbox_0_T6, SubBytesIns_Inst_Sbox_0_T5,
         SubBytesIns_Inst_Sbox_0_T4, SubBytesIns_Inst_Sbox_0_T3,
         SubBytesIns_Inst_Sbox_0_T2, SubBytesIns_Inst_Sbox_0_T1,
         SubBytesIns_Inst_Sbox_1_L29, SubBytesIns_Inst_Sbox_1_L28,
         SubBytesIns_Inst_Sbox_1_L27, SubBytesIns_Inst_Sbox_1_L26,
         SubBytesIns_Inst_Sbox_1_L25, SubBytesIns_Inst_Sbox_1_L24,
         SubBytesIns_Inst_Sbox_1_L23, SubBytesIns_Inst_Sbox_1_L22,
         SubBytesIns_Inst_Sbox_1_L21, SubBytesIns_Inst_Sbox_1_L20,
         SubBytesIns_Inst_Sbox_1_L19, SubBytesIns_Inst_Sbox_1_L18,
         SubBytesIns_Inst_Sbox_1_L17, SubBytesIns_Inst_Sbox_1_L16,
         SubBytesIns_Inst_Sbox_1_L15, SubBytesIns_Inst_Sbox_1_L14,
         SubBytesIns_Inst_Sbox_1_L13, SubBytesIns_Inst_Sbox_1_L12,
         SubBytesIns_Inst_Sbox_1_L11, SubBytesIns_Inst_Sbox_1_L10,
         SubBytesIns_Inst_Sbox_1_L9, SubBytesIns_Inst_Sbox_1_L8,
         SubBytesIns_Inst_Sbox_1_L7, SubBytesIns_Inst_Sbox_1_L6,
         SubBytesIns_Inst_Sbox_1_L5, SubBytesIns_Inst_Sbox_1_L4,
         SubBytesIns_Inst_Sbox_1_L3, SubBytesIns_Inst_Sbox_1_L2,
         SubBytesIns_Inst_Sbox_1_L1, SubBytesIns_Inst_Sbox_1_L0,
         SubBytesIns_Inst_Sbox_1_M63, SubBytesIns_Inst_Sbox_1_M62,
         SubBytesIns_Inst_Sbox_1_M61, SubBytesIns_Inst_Sbox_1_M60,
         SubBytesIns_Inst_Sbox_1_M59, SubBytesIns_Inst_Sbox_1_M58,
         SubBytesIns_Inst_Sbox_1_M57, SubBytesIns_Inst_Sbox_1_M56,
         SubBytesIns_Inst_Sbox_1_M55, SubBytesIns_Inst_Sbox_1_M54,
         SubBytesIns_Inst_Sbox_1_M53, SubBytesIns_Inst_Sbox_1_M52,
         SubBytesIns_Inst_Sbox_1_M51, SubBytesIns_Inst_Sbox_1_M50,
         SubBytesIns_Inst_Sbox_1_M49, SubBytesIns_Inst_Sbox_1_M48,
         SubBytesIns_Inst_Sbox_1_M47, SubBytesIns_Inst_Sbox_1_M46,
         SubBytesIns_Inst_Sbox_1_M45, SubBytesIns_Inst_Sbox_1_M44,
         SubBytesIns_Inst_Sbox_1_M43, SubBytesIns_Inst_Sbox_1_M42,
         SubBytesIns_Inst_Sbox_1_M41, SubBytesIns_Inst_Sbox_1_M40,
         SubBytesIns_Inst_Sbox_1_M39, SubBytesIns_Inst_Sbox_1_M38,
         SubBytesIns_Inst_Sbox_1_M37, SubBytesIns_Inst_Sbox_1_M36,
         SubBytesIns_Inst_Sbox_1_M35, SubBytesIns_Inst_Sbox_1_M34,
         SubBytesIns_Inst_Sbox_1_M33, SubBytesIns_Inst_Sbox_1_M32,
         SubBytesIns_Inst_Sbox_1_M31, SubBytesIns_Inst_Sbox_1_M30,
         SubBytesIns_Inst_Sbox_1_M29, SubBytesIns_Inst_Sbox_1_M28,
         SubBytesIns_Inst_Sbox_1_M27, SubBytesIns_Inst_Sbox_1_M26,
         SubBytesIns_Inst_Sbox_1_M25, SubBytesIns_Inst_Sbox_1_M24,
         SubBytesIns_Inst_Sbox_1_M23, SubBytesIns_Inst_Sbox_1_M22,
         SubBytesIns_Inst_Sbox_1_M21, SubBytesIns_Inst_Sbox_1_M20,
         SubBytesIns_Inst_Sbox_1_M19, SubBytesIns_Inst_Sbox_1_M18,
         SubBytesIns_Inst_Sbox_1_M17, SubBytesIns_Inst_Sbox_1_M16,
         SubBytesIns_Inst_Sbox_1_M15, SubBytesIns_Inst_Sbox_1_M14,
         SubBytesIns_Inst_Sbox_1_M13, SubBytesIns_Inst_Sbox_1_M12,
         SubBytesIns_Inst_Sbox_1_M11, SubBytesIns_Inst_Sbox_1_M10,
         SubBytesIns_Inst_Sbox_1_M9, SubBytesIns_Inst_Sbox_1_M8,
         SubBytesIns_Inst_Sbox_1_M7, SubBytesIns_Inst_Sbox_1_M6,
         SubBytesIns_Inst_Sbox_1_M5, SubBytesIns_Inst_Sbox_1_M4,
         SubBytesIns_Inst_Sbox_1_M3, SubBytesIns_Inst_Sbox_1_M2,
         SubBytesIns_Inst_Sbox_1_M1, SubBytesIns_Inst_Sbox_1_T27,
         SubBytesIns_Inst_Sbox_1_T26, SubBytesIns_Inst_Sbox_1_T25,
         SubBytesIns_Inst_Sbox_1_T24, SubBytesIns_Inst_Sbox_1_T23,
         SubBytesIns_Inst_Sbox_1_T22, SubBytesIns_Inst_Sbox_1_T21,
         SubBytesIns_Inst_Sbox_1_T20, SubBytesIns_Inst_Sbox_1_T19,
         SubBytesIns_Inst_Sbox_1_T18, SubBytesIns_Inst_Sbox_1_T17,
         SubBytesIns_Inst_Sbox_1_T16, SubBytesIns_Inst_Sbox_1_T15,
         SubBytesIns_Inst_Sbox_1_T14, SubBytesIns_Inst_Sbox_1_T13,
         SubBytesIns_Inst_Sbox_1_T12, SubBytesIns_Inst_Sbox_1_T11,
         SubBytesIns_Inst_Sbox_1_T10, SubBytesIns_Inst_Sbox_1_T9,
         SubBytesIns_Inst_Sbox_1_T8, SubBytesIns_Inst_Sbox_1_T7,
         SubBytesIns_Inst_Sbox_1_T6, SubBytesIns_Inst_Sbox_1_T5,
         SubBytesIns_Inst_Sbox_1_T4, SubBytesIns_Inst_Sbox_1_T3,
         SubBytesIns_Inst_Sbox_1_T2, SubBytesIns_Inst_Sbox_1_T1,
         SubBytesIns_Inst_Sbox_2_L29, SubBytesIns_Inst_Sbox_2_L28,
         SubBytesIns_Inst_Sbox_2_L27, SubBytesIns_Inst_Sbox_2_L26,
         SubBytesIns_Inst_Sbox_2_L25, SubBytesIns_Inst_Sbox_2_L24,
         SubBytesIns_Inst_Sbox_2_L23, SubBytesIns_Inst_Sbox_2_L22,
         SubBytesIns_Inst_Sbox_2_L21, SubBytesIns_Inst_Sbox_2_L20,
         SubBytesIns_Inst_Sbox_2_L19, SubBytesIns_Inst_Sbox_2_L18,
         SubBytesIns_Inst_Sbox_2_L17, SubBytesIns_Inst_Sbox_2_L16,
         SubBytesIns_Inst_Sbox_2_L15, SubBytesIns_Inst_Sbox_2_L14,
         SubBytesIns_Inst_Sbox_2_L13, SubBytesIns_Inst_Sbox_2_L12,
         SubBytesIns_Inst_Sbox_2_L11, SubBytesIns_Inst_Sbox_2_L10,
         SubBytesIns_Inst_Sbox_2_L9, SubBytesIns_Inst_Sbox_2_L8,
         SubBytesIns_Inst_Sbox_2_L7, SubBytesIns_Inst_Sbox_2_L6,
         SubBytesIns_Inst_Sbox_2_L5, SubBytesIns_Inst_Sbox_2_L4,
         SubBytesIns_Inst_Sbox_2_L3, SubBytesIns_Inst_Sbox_2_L2,
         SubBytesIns_Inst_Sbox_2_L1, SubBytesIns_Inst_Sbox_2_L0,
         SubBytesIns_Inst_Sbox_2_M63, SubBytesIns_Inst_Sbox_2_M62,
         SubBytesIns_Inst_Sbox_2_M61, SubBytesIns_Inst_Sbox_2_M60,
         SubBytesIns_Inst_Sbox_2_M59, SubBytesIns_Inst_Sbox_2_M58,
         SubBytesIns_Inst_Sbox_2_M57, SubBytesIns_Inst_Sbox_2_M56,
         SubBytesIns_Inst_Sbox_2_M55, SubBytesIns_Inst_Sbox_2_M54,
         SubBytesIns_Inst_Sbox_2_M53, SubBytesIns_Inst_Sbox_2_M52,
         SubBytesIns_Inst_Sbox_2_M51, SubBytesIns_Inst_Sbox_2_M50,
         SubBytesIns_Inst_Sbox_2_M49, SubBytesIns_Inst_Sbox_2_M48,
         SubBytesIns_Inst_Sbox_2_M47, SubBytesIns_Inst_Sbox_2_M46,
         SubBytesIns_Inst_Sbox_2_M45, SubBytesIns_Inst_Sbox_2_M44,
         SubBytesIns_Inst_Sbox_2_M43, SubBytesIns_Inst_Sbox_2_M42,
         SubBytesIns_Inst_Sbox_2_M41, SubBytesIns_Inst_Sbox_2_M40,
         SubBytesIns_Inst_Sbox_2_M39, SubBytesIns_Inst_Sbox_2_M38,
         SubBytesIns_Inst_Sbox_2_M37, SubBytesIns_Inst_Sbox_2_M36,
         SubBytesIns_Inst_Sbox_2_M35, SubBytesIns_Inst_Sbox_2_M34,
         SubBytesIns_Inst_Sbox_2_M33, SubBytesIns_Inst_Sbox_2_M32,
         SubBytesIns_Inst_Sbox_2_M31, SubBytesIns_Inst_Sbox_2_M30,
         SubBytesIns_Inst_Sbox_2_M29, SubBytesIns_Inst_Sbox_2_M28,
         SubBytesIns_Inst_Sbox_2_M27, SubBytesIns_Inst_Sbox_2_M26,
         SubBytesIns_Inst_Sbox_2_M25, SubBytesIns_Inst_Sbox_2_M24,
         SubBytesIns_Inst_Sbox_2_M23, SubBytesIns_Inst_Sbox_2_M22,
         SubBytesIns_Inst_Sbox_2_M21, SubBytesIns_Inst_Sbox_2_M20,
         SubBytesIns_Inst_Sbox_2_M19, SubBytesIns_Inst_Sbox_2_M18,
         SubBytesIns_Inst_Sbox_2_M17, SubBytesIns_Inst_Sbox_2_M16,
         SubBytesIns_Inst_Sbox_2_M15, SubBytesIns_Inst_Sbox_2_M14,
         SubBytesIns_Inst_Sbox_2_M13, SubBytesIns_Inst_Sbox_2_M12,
         SubBytesIns_Inst_Sbox_2_M11, SubBytesIns_Inst_Sbox_2_M10,
         SubBytesIns_Inst_Sbox_2_M9, SubBytesIns_Inst_Sbox_2_M8,
         SubBytesIns_Inst_Sbox_2_M7, SubBytesIns_Inst_Sbox_2_M6,
         SubBytesIns_Inst_Sbox_2_M5, SubBytesIns_Inst_Sbox_2_M4,
         SubBytesIns_Inst_Sbox_2_M3, SubBytesIns_Inst_Sbox_2_M2,
         SubBytesIns_Inst_Sbox_2_M1, SubBytesIns_Inst_Sbox_2_T27,
         SubBytesIns_Inst_Sbox_2_T26, SubBytesIns_Inst_Sbox_2_T25,
         SubBytesIns_Inst_Sbox_2_T24, SubBytesIns_Inst_Sbox_2_T23,
         SubBytesIns_Inst_Sbox_2_T22, SubBytesIns_Inst_Sbox_2_T21,
         SubBytesIns_Inst_Sbox_2_T20, SubBytesIns_Inst_Sbox_2_T19,
         SubBytesIns_Inst_Sbox_2_T18, SubBytesIns_Inst_Sbox_2_T17,
         SubBytesIns_Inst_Sbox_2_T16, SubBytesIns_Inst_Sbox_2_T15,
         SubBytesIns_Inst_Sbox_2_T14, SubBytesIns_Inst_Sbox_2_T13,
         SubBytesIns_Inst_Sbox_2_T12, SubBytesIns_Inst_Sbox_2_T11,
         SubBytesIns_Inst_Sbox_2_T10, SubBytesIns_Inst_Sbox_2_T9,
         SubBytesIns_Inst_Sbox_2_T8, SubBytesIns_Inst_Sbox_2_T7,
         SubBytesIns_Inst_Sbox_2_T6, SubBytesIns_Inst_Sbox_2_T5,
         SubBytesIns_Inst_Sbox_2_T4, SubBytesIns_Inst_Sbox_2_T3,
         SubBytesIns_Inst_Sbox_2_T2, SubBytesIns_Inst_Sbox_2_T1,
         SubBytesIns_Inst_Sbox_3_L29, SubBytesIns_Inst_Sbox_3_L28,
         SubBytesIns_Inst_Sbox_3_L27, SubBytesIns_Inst_Sbox_3_L26,
         SubBytesIns_Inst_Sbox_3_L25, SubBytesIns_Inst_Sbox_3_L24,
         SubBytesIns_Inst_Sbox_3_L23, SubBytesIns_Inst_Sbox_3_L22,
         SubBytesIns_Inst_Sbox_3_L21, SubBytesIns_Inst_Sbox_3_L20,
         SubBytesIns_Inst_Sbox_3_L19, SubBytesIns_Inst_Sbox_3_L18,
         SubBytesIns_Inst_Sbox_3_L17, SubBytesIns_Inst_Sbox_3_L16,
         SubBytesIns_Inst_Sbox_3_L15, SubBytesIns_Inst_Sbox_3_L14,
         SubBytesIns_Inst_Sbox_3_L13, SubBytesIns_Inst_Sbox_3_L12,
         SubBytesIns_Inst_Sbox_3_L11, SubBytesIns_Inst_Sbox_3_L10,
         SubBytesIns_Inst_Sbox_3_L9, SubBytesIns_Inst_Sbox_3_L8,
         SubBytesIns_Inst_Sbox_3_L7, SubBytesIns_Inst_Sbox_3_L6,
         SubBytesIns_Inst_Sbox_3_L5, SubBytesIns_Inst_Sbox_3_L4,
         SubBytesIns_Inst_Sbox_3_L3, SubBytesIns_Inst_Sbox_3_L2,
         SubBytesIns_Inst_Sbox_3_L1, SubBytesIns_Inst_Sbox_3_L0,
         SubBytesIns_Inst_Sbox_3_M63, SubBytesIns_Inst_Sbox_3_M62,
         SubBytesIns_Inst_Sbox_3_M61, SubBytesIns_Inst_Sbox_3_M60,
         SubBytesIns_Inst_Sbox_3_M59, SubBytesIns_Inst_Sbox_3_M58,
         SubBytesIns_Inst_Sbox_3_M57, SubBytesIns_Inst_Sbox_3_M56,
         SubBytesIns_Inst_Sbox_3_M55, SubBytesIns_Inst_Sbox_3_M54,
         SubBytesIns_Inst_Sbox_3_M53, SubBytesIns_Inst_Sbox_3_M52,
         SubBytesIns_Inst_Sbox_3_M51, SubBytesIns_Inst_Sbox_3_M50,
         SubBytesIns_Inst_Sbox_3_M49, SubBytesIns_Inst_Sbox_3_M48,
         SubBytesIns_Inst_Sbox_3_M47, SubBytesIns_Inst_Sbox_3_M46,
         SubBytesIns_Inst_Sbox_3_M45, SubBytesIns_Inst_Sbox_3_M44,
         SubBytesIns_Inst_Sbox_3_M43, SubBytesIns_Inst_Sbox_3_M42,
         SubBytesIns_Inst_Sbox_3_M41, SubBytesIns_Inst_Sbox_3_M40,
         SubBytesIns_Inst_Sbox_3_M39, SubBytesIns_Inst_Sbox_3_M38,
         SubBytesIns_Inst_Sbox_3_M37, SubBytesIns_Inst_Sbox_3_M36,
         SubBytesIns_Inst_Sbox_3_M35, SubBytesIns_Inst_Sbox_3_M34,
         SubBytesIns_Inst_Sbox_3_M33, SubBytesIns_Inst_Sbox_3_M32,
         SubBytesIns_Inst_Sbox_3_M31, SubBytesIns_Inst_Sbox_3_M30,
         SubBytesIns_Inst_Sbox_3_M29, SubBytesIns_Inst_Sbox_3_M28,
         SubBytesIns_Inst_Sbox_3_M27, SubBytesIns_Inst_Sbox_3_M26,
         SubBytesIns_Inst_Sbox_3_M25, SubBytesIns_Inst_Sbox_3_M24,
         SubBytesIns_Inst_Sbox_3_M23, SubBytesIns_Inst_Sbox_3_M22,
         SubBytesIns_Inst_Sbox_3_M21, SubBytesIns_Inst_Sbox_3_M20,
         SubBytesIns_Inst_Sbox_3_M19, SubBytesIns_Inst_Sbox_3_M18,
         SubBytesIns_Inst_Sbox_3_M17, SubBytesIns_Inst_Sbox_3_M16,
         SubBytesIns_Inst_Sbox_3_M15, SubBytesIns_Inst_Sbox_3_M14,
         SubBytesIns_Inst_Sbox_3_M13, SubBytesIns_Inst_Sbox_3_M12,
         SubBytesIns_Inst_Sbox_3_M11, SubBytesIns_Inst_Sbox_3_M10,
         SubBytesIns_Inst_Sbox_3_M9, SubBytesIns_Inst_Sbox_3_M8,
         SubBytesIns_Inst_Sbox_3_M7, SubBytesIns_Inst_Sbox_3_M6,
         SubBytesIns_Inst_Sbox_3_M5, SubBytesIns_Inst_Sbox_3_M4,
         SubBytesIns_Inst_Sbox_3_M3, SubBytesIns_Inst_Sbox_3_M2,
         SubBytesIns_Inst_Sbox_3_M1, SubBytesIns_Inst_Sbox_3_T27,
         SubBytesIns_Inst_Sbox_3_T26, SubBytesIns_Inst_Sbox_3_T25,
         SubBytesIns_Inst_Sbox_3_T24, SubBytesIns_Inst_Sbox_3_T23,
         SubBytesIns_Inst_Sbox_3_T22, SubBytesIns_Inst_Sbox_3_T21,
         SubBytesIns_Inst_Sbox_3_T20, SubBytesIns_Inst_Sbox_3_T19,
         SubBytesIns_Inst_Sbox_3_T18, SubBytesIns_Inst_Sbox_3_T17,
         SubBytesIns_Inst_Sbox_3_T16, SubBytesIns_Inst_Sbox_3_T15,
         SubBytesIns_Inst_Sbox_3_T14, SubBytesIns_Inst_Sbox_3_T13,
         SubBytesIns_Inst_Sbox_3_T12, SubBytesIns_Inst_Sbox_3_T11,
         SubBytesIns_Inst_Sbox_3_T10, SubBytesIns_Inst_Sbox_3_T9,
         SubBytesIns_Inst_Sbox_3_T8, SubBytesIns_Inst_Sbox_3_T7,
         SubBytesIns_Inst_Sbox_3_T6, SubBytesIns_Inst_Sbox_3_T5,
         SubBytesIns_Inst_Sbox_3_T4, SubBytesIns_Inst_Sbox_3_T3,
         SubBytesIns_Inst_Sbox_3_T2, SubBytesIns_Inst_Sbox_3_T1,
         SubBytesIns_Inst_Sbox_4_L29, SubBytesIns_Inst_Sbox_4_L28,
         SubBytesIns_Inst_Sbox_4_L27, SubBytesIns_Inst_Sbox_4_L26,
         SubBytesIns_Inst_Sbox_4_L25, SubBytesIns_Inst_Sbox_4_L24,
         SubBytesIns_Inst_Sbox_4_L23, SubBytesIns_Inst_Sbox_4_L22,
         SubBytesIns_Inst_Sbox_4_L21, SubBytesIns_Inst_Sbox_4_L20,
         SubBytesIns_Inst_Sbox_4_L19, SubBytesIns_Inst_Sbox_4_L18,
         SubBytesIns_Inst_Sbox_4_L17, SubBytesIns_Inst_Sbox_4_L16,
         SubBytesIns_Inst_Sbox_4_L15, SubBytesIns_Inst_Sbox_4_L14,
         SubBytesIns_Inst_Sbox_4_L13, SubBytesIns_Inst_Sbox_4_L12,
         SubBytesIns_Inst_Sbox_4_L11, SubBytesIns_Inst_Sbox_4_L10,
         SubBytesIns_Inst_Sbox_4_L9, SubBytesIns_Inst_Sbox_4_L8,
         SubBytesIns_Inst_Sbox_4_L7, SubBytesIns_Inst_Sbox_4_L6,
         SubBytesIns_Inst_Sbox_4_L5, SubBytesIns_Inst_Sbox_4_L4,
         SubBytesIns_Inst_Sbox_4_L3, SubBytesIns_Inst_Sbox_4_L2,
         SubBytesIns_Inst_Sbox_4_L1, SubBytesIns_Inst_Sbox_4_L0,
         SubBytesIns_Inst_Sbox_4_M63, SubBytesIns_Inst_Sbox_4_M62,
         SubBytesIns_Inst_Sbox_4_M61, SubBytesIns_Inst_Sbox_4_M60,
         SubBytesIns_Inst_Sbox_4_M59, SubBytesIns_Inst_Sbox_4_M58,
         SubBytesIns_Inst_Sbox_4_M57, SubBytesIns_Inst_Sbox_4_M56,
         SubBytesIns_Inst_Sbox_4_M55, SubBytesIns_Inst_Sbox_4_M54,
         SubBytesIns_Inst_Sbox_4_M53, SubBytesIns_Inst_Sbox_4_M52,
         SubBytesIns_Inst_Sbox_4_M51, SubBytesIns_Inst_Sbox_4_M50,
         SubBytesIns_Inst_Sbox_4_M49, SubBytesIns_Inst_Sbox_4_M48,
         SubBytesIns_Inst_Sbox_4_M47, SubBytesIns_Inst_Sbox_4_M46,
         SubBytesIns_Inst_Sbox_4_M45, SubBytesIns_Inst_Sbox_4_M44,
         SubBytesIns_Inst_Sbox_4_M43, SubBytesIns_Inst_Sbox_4_M42,
         SubBytesIns_Inst_Sbox_4_M41, SubBytesIns_Inst_Sbox_4_M40,
         SubBytesIns_Inst_Sbox_4_M39, SubBytesIns_Inst_Sbox_4_M38,
         SubBytesIns_Inst_Sbox_4_M37, SubBytesIns_Inst_Sbox_4_M36,
         SubBytesIns_Inst_Sbox_4_M35, SubBytesIns_Inst_Sbox_4_M34,
         SubBytesIns_Inst_Sbox_4_M33, SubBytesIns_Inst_Sbox_4_M32,
         SubBytesIns_Inst_Sbox_4_M31, SubBytesIns_Inst_Sbox_4_M30,
         SubBytesIns_Inst_Sbox_4_M29, SubBytesIns_Inst_Sbox_4_M28,
         SubBytesIns_Inst_Sbox_4_M27, SubBytesIns_Inst_Sbox_4_M26,
         SubBytesIns_Inst_Sbox_4_M25, SubBytesIns_Inst_Sbox_4_M24,
         SubBytesIns_Inst_Sbox_4_M23, SubBytesIns_Inst_Sbox_4_M22,
         SubBytesIns_Inst_Sbox_4_M21, SubBytesIns_Inst_Sbox_4_M20,
         SubBytesIns_Inst_Sbox_4_M19, SubBytesIns_Inst_Sbox_4_M18,
         SubBytesIns_Inst_Sbox_4_M17, SubBytesIns_Inst_Sbox_4_M16,
         SubBytesIns_Inst_Sbox_4_M15, SubBytesIns_Inst_Sbox_4_M14,
         SubBytesIns_Inst_Sbox_4_M13, SubBytesIns_Inst_Sbox_4_M12,
         SubBytesIns_Inst_Sbox_4_M11, SubBytesIns_Inst_Sbox_4_M10,
         SubBytesIns_Inst_Sbox_4_M9, SubBytesIns_Inst_Sbox_4_M8,
         SubBytesIns_Inst_Sbox_4_M7, SubBytesIns_Inst_Sbox_4_M6,
         SubBytesIns_Inst_Sbox_4_M5, SubBytesIns_Inst_Sbox_4_M4,
         SubBytesIns_Inst_Sbox_4_M3, SubBytesIns_Inst_Sbox_4_M2,
         SubBytesIns_Inst_Sbox_4_M1, SubBytesIns_Inst_Sbox_4_T27,
         SubBytesIns_Inst_Sbox_4_T26, SubBytesIns_Inst_Sbox_4_T25,
         SubBytesIns_Inst_Sbox_4_T24, SubBytesIns_Inst_Sbox_4_T23,
         SubBytesIns_Inst_Sbox_4_T22, SubBytesIns_Inst_Sbox_4_T21,
         SubBytesIns_Inst_Sbox_4_T20, SubBytesIns_Inst_Sbox_4_T19,
         SubBytesIns_Inst_Sbox_4_T18, SubBytesIns_Inst_Sbox_4_T17,
         SubBytesIns_Inst_Sbox_4_T16, SubBytesIns_Inst_Sbox_4_T15,
         SubBytesIns_Inst_Sbox_4_T14, SubBytesIns_Inst_Sbox_4_T13,
         SubBytesIns_Inst_Sbox_4_T12, SubBytesIns_Inst_Sbox_4_T11,
         SubBytesIns_Inst_Sbox_4_T10, SubBytesIns_Inst_Sbox_4_T9,
         SubBytesIns_Inst_Sbox_4_T8, SubBytesIns_Inst_Sbox_4_T7,
         SubBytesIns_Inst_Sbox_4_T6, SubBytesIns_Inst_Sbox_4_T5,
         SubBytesIns_Inst_Sbox_4_T4, SubBytesIns_Inst_Sbox_4_T3,
         SubBytesIns_Inst_Sbox_4_T2, SubBytesIns_Inst_Sbox_4_T1,
         SubBytesIns_Inst_Sbox_5_L29, SubBytesIns_Inst_Sbox_5_L28,
         SubBytesIns_Inst_Sbox_5_L27, SubBytesIns_Inst_Sbox_5_L26,
         SubBytesIns_Inst_Sbox_5_L25, SubBytesIns_Inst_Sbox_5_L24,
         SubBytesIns_Inst_Sbox_5_L23, SubBytesIns_Inst_Sbox_5_L22,
         SubBytesIns_Inst_Sbox_5_L21, SubBytesIns_Inst_Sbox_5_L20,
         SubBytesIns_Inst_Sbox_5_L19, SubBytesIns_Inst_Sbox_5_L18,
         SubBytesIns_Inst_Sbox_5_L17, SubBytesIns_Inst_Sbox_5_L16,
         SubBytesIns_Inst_Sbox_5_L15, SubBytesIns_Inst_Sbox_5_L14,
         SubBytesIns_Inst_Sbox_5_L13, SubBytesIns_Inst_Sbox_5_L12,
         SubBytesIns_Inst_Sbox_5_L11, SubBytesIns_Inst_Sbox_5_L10,
         SubBytesIns_Inst_Sbox_5_L9, SubBytesIns_Inst_Sbox_5_L8,
         SubBytesIns_Inst_Sbox_5_L7, SubBytesIns_Inst_Sbox_5_L6,
         SubBytesIns_Inst_Sbox_5_L5, SubBytesIns_Inst_Sbox_5_L4,
         SubBytesIns_Inst_Sbox_5_L3, SubBytesIns_Inst_Sbox_5_L2,
         SubBytesIns_Inst_Sbox_5_L1, SubBytesIns_Inst_Sbox_5_L0,
         SubBytesIns_Inst_Sbox_5_M63, SubBytesIns_Inst_Sbox_5_M62,
         SubBytesIns_Inst_Sbox_5_M61, SubBytesIns_Inst_Sbox_5_M60,
         SubBytesIns_Inst_Sbox_5_M59, SubBytesIns_Inst_Sbox_5_M58,
         SubBytesIns_Inst_Sbox_5_M57, SubBytesIns_Inst_Sbox_5_M56,
         SubBytesIns_Inst_Sbox_5_M55, SubBytesIns_Inst_Sbox_5_M54,
         SubBytesIns_Inst_Sbox_5_M53, SubBytesIns_Inst_Sbox_5_M52,
         SubBytesIns_Inst_Sbox_5_M51, SubBytesIns_Inst_Sbox_5_M50,
         SubBytesIns_Inst_Sbox_5_M49, SubBytesIns_Inst_Sbox_5_M48,
         SubBytesIns_Inst_Sbox_5_M47, SubBytesIns_Inst_Sbox_5_M46,
         SubBytesIns_Inst_Sbox_5_M45, SubBytesIns_Inst_Sbox_5_M44,
         SubBytesIns_Inst_Sbox_5_M43, SubBytesIns_Inst_Sbox_5_M42,
         SubBytesIns_Inst_Sbox_5_M41, SubBytesIns_Inst_Sbox_5_M40,
         SubBytesIns_Inst_Sbox_5_M39, SubBytesIns_Inst_Sbox_5_M38,
         SubBytesIns_Inst_Sbox_5_M37, SubBytesIns_Inst_Sbox_5_M36,
         SubBytesIns_Inst_Sbox_5_M35, SubBytesIns_Inst_Sbox_5_M34,
         SubBytesIns_Inst_Sbox_5_M33, SubBytesIns_Inst_Sbox_5_M32,
         SubBytesIns_Inst_Sbox_5_M31, SubBytesIns_Inst_Sbox_5_M30,
         SubBytesIns_Inst_Sbox_5_M29, SubBytesIns_Inst_Sbox_5_M28,
         SubBytesIns_Inst_Sbox_5_M27, SubBytesIns_Inst_Sbox_5_M26,
         SubBytesIns_Inst_Sbox_5_M25, SubBytesIns_Inst_Sbox_5_M24,
         SubBytesIns_Inst_Sbox_5_M23, SubBytesIns_Inst_Sbox_5_M22,
         SubBytesIns_Inst_Sbox_5_M21, SubBytesIns_Inst_Sbox_5_M20,
         SubBytesIns_Inst_Sbox_5_M19, SubBytesIns_Inst_Sbox_5_M18,
         SubBytesIns_Inst_Sbox_5_M17, SubBytesIns_Inst_Sbox_5_M16,
         SubBytesIns_Inst_Sbox_5_M15, SubBytesIns_Inst_Sbox_5_M14,
         SubBytesIns_Inst_Sbox_5_M13, SubBytesIns_Inst_Sbox_5_M12,
         SubBytesIns_Inst_Sbox_5_M11, SubBytesIns_Inst_Sbox_5_M10,
         SubBytesIns_Inst_Sbox_5_M9, SubBytesIns_Inst_Sbox_5_M8,
         SubBytesIns_Inst_Sbox_5_M7, SubBytesIns_Inst_Sbox_5_M6,
         SubBytesIns_Inst_Sbox_5_M5, SubBytesIns_Inst_Sbox_5_M4,
         SubBytesIns_Inst_Sbox_5_M3, SubBytesIns_Inst_Sbox_5_M2,
         SubBytesIns_Inst_Sbox_5_M1, SubBytesIns_Inst_Sbox_5_T27,
         SubBytesIns_Inst_Sbox_5_T26, SubBytesIns_Inst_Sbox_5_T25,
         SubBytesIns_Inst_Sbox_5_T24, SubBytesIns_Inst_Sbox_5_T23,
         SubBytesIns_Inst_Sbox_5_T22, SubBytesIns_Inst_Sbox_5_T21,
         SubBytesIns_Inst_Sbox_5_T20, SubBytesIns_Inst_Sbox_5_T19,
         SubBytesIns_Inst_Sbox_5_T18, SubBytesIns_Inst_Sbox_5_T17,
         SubBytesIns_Inst_Sbox_5_T16, SubBytesIns_Inst_Sbox_5_T15,
         SubBytesIns_Inst_Sbox_5_T14, SubBytesIns_Inst_Sbox_5_T13,
         SubBytesIns_Inst_Sbox_5_T12, SubBytesIns_Inst_Sbox_5_T11,
         SubBytesIns_Inst_Sbox_5_T10, SubBytesIns_Inst_Sbox_5_T9,
         SubBytesIns_Inst_Sbox_5_T8, SubBytesIns_Inst_Sbox_5_T7,
         SubBytesIns_Inst_Sbox_5_T6, SubBytesIns_Inst_Sbox_5_T5,
         SubBytesIns_Inst_Sbox_5_T4, SubBytesIns_Inst_Sbox_5_T3,
         SubBytesIns_Inst_Sbox_5_T2, SubBytesIns_Inst_Sbox_5_T1,
         SubBytesIns_Inst_Sbox_6_L29, SubBytesIns_Inst_Sbox_6_L28,
         SubBytesIns_Inst_Sbox_6_L27, SubBytesIns_Inst_Sbox_6_L26,
         SubBytesIns_Inst_Sbox_6_L25, SubBytesIns_Inst_Sbox_6_L24,
         SubBytesIns_Inst_Sbox_6_L23, SubBytesIns_Inst_Sbox_6_L22,
         SubBytesIns_Inst_Sbox_6_L21, SubBytesIns_Inst_Sbox_6_L20,
         SubBytesIns_Inst_Sbox_6_L19, SubBytesIns_Inst_Sbox_6_L18,
         SubBytesIns_Inst_Sbox_6_L17, SubBytesIns_Inst_Sbox_6_L16,
         SubBytesIns_Inst_Sbox_6_L15, SubBytesIns_Inst_Sbox_6_L14,
         SubBytesIns_Inst_Sbox_6_L13, SubBytesIns_Inst_Sbox_6_L12,
         SubBytesIns_Inst_Sbox_6_L11, SubBytesIns_Inst_Sbox_6_L10,
         SubBytesIns_Inst_Sbox_6_L9, SubBytesIns_Inst_Sbox_6_L8,
         SubBytesIns_Inst_Sbox_6_L7, SubBytesIns_Inst_Sbox_6_L6,
         SubBytesIns_Inst_Sbox_6_L5, SubBytesIns_Inst_Sbox_6_L4,
         SubBytesIns_Inst_Sbox_6_L3, SubBytesIns_Inst_Sbox_6_L2,
         SubBytesIns_Inst_Sbox_6_L1, SubBytesIns_Inst_Sbox_6_L0,
         SubBytesIns_Inst_Sbox_6_M63, SubBytesIns_Inst_Sbox_6_M62,
         SubBytesIns_Inst_Sbox_6_M61, SubBytesIns_Inst_Sbox_6_M60,
         SubBytesIns_Inst_Sbox_6_M59, SubBytesIns_Inst_Sbox_6_M58,
         SubBytesIns_Inst_Sbox_6_M57, SubBytesIns_Inst_Sbox_6_M56,
         SubBytesIns_Inst_Sbox_6_M55, SubBytesIns_Inst_Sbox_6_M54,
         SubBytesIns_Inst_Sbox_6_M53, SubBytesIns_Inst_Sbox_6_M52,
         SubBytesIns_Inst_Sbox_6_M51, SubBytesIns_Inst_Sbox_6_M50,
         SubBytesIns_Inst_Sbox_6_M49, SubBytesIns_Inst_Sbox_6_M48,
         SubBytesIns_Inst_Sbox_6_M47, SubBytesIns_Inst_Sbox_6_M46,
         SubBytesIns_Inst_Sbox_6_M45, SubBytesIns_Inst_Sbox_6_M44,
         SubBytesIns_Inst_Sbox_6_M43, SubBytesIns_Inst_Sbox_6_M42,
         SubBytesIns_Inst_Sbox_6_M41, SubBytesIns_Inst_Sbox_6_M40,
         SubBytesIns_Inst_Sbox_6_M39, SubBytesIns_Inst_Sbox_6_M38,
         SubBytesIns_Inst_Sbox_6_M37, SubBytesIns_Inst_Sbox_6_M36,
         SubBytesIns_Inst_Sbox_6_M35, SubBytesIns_Inst_Sbox_6_M34,
         SubBytesIns_Inst_Sbox_6_M33, SubBytesIns_Inst_Sbox_6_M32,
         SubBytesIns_Inst_Sbox_6_M31, SubBytesIns_Inst_Sbox_6_M30,
         SubBytesIns_Inst_Sbox_6_M29, SubBytesIns_Inst_Sbox_6_M28,
         SubBytesIns_Inst_Sbox_6_M27, SubBytesIns_Inst_Sbox_6_M26,
         SubBytesIns_Inst_Sbox_6_M25, SubBytesIns_Inst_Sbox_6_M24,
         SubBytesIns_Inst_Sbox_6_M23, SubBytesIns_Inst_Sbox_6_M22,
         SubBytesIns_Inst_Sbox_6_M21, SubBytesIns_Inst_Sbox_6_M20,
         SubBytesIns_Inst_Sbox_6_M19, SubBytesIns_Inst_Sbox_6_M18,
         SubBytesIns_Inst_Sbox_6_M17, SubBytesIns_Inst_Sbox_6_M16,
         SubBytesIns_Inst_Sbox_6_M15, SubBytesIns_Inst_Sbox_6_M14,
         SubBytesIns_Inst_Sbox_6_M13, SubBytesIns_Inst_Sbox_6_M12,
         SubBytesIns_Inst_Sbox_6_M11, SubBytesIns_Inst_Sbox_6_M10,
         SubBytesIns_Inst_Sbox_6_M9, SubBytesIns_Inst_Sbox_6_M8,
         SubBytesIns_Inst_Sbox_6_M7, SubBytesIns_Inst_Sbox_6_M6,
         SubBytesIns_Inst_Sbox_6_M5, SubBytesIns_Inst_Sbox_6_M4,
         SubBytesIns_Inst_Sbox_6_M3, SubBytesIns_Inst_Sbox_6_M2,
         SubBytesIns_Inst_Sbox_6_M1, SubBytesIns_Inst_Sbox_6_T27,
         SubBytesIns_Inst_Sbox_6_T26, SubBytesIns_Inst_Sbox_6_T25,
         SubBytesIns_Inst_Sbox_6_T24, SubBytesIns_Inst_Sbox_6_T23,
         SubBytesIns_Inst_Sbox_6_T22, SubBytesIns_Inst_Sbox_6_T21,
         SubBytesIns_Inst_Sbox_6_T20, SubBytesIns_Inst_Sbox_6_T19,
         SubBytesIns_Inst_Sbox_6_T18, SubBytesIns_Inst_Sbox_6_T17,
         SubBytesIns_Inst_Sbox_6_T16, SubBytesIns_Inst_Sbox_6_T15,
         SubBytesIns_Inst_Sbox_6_T14, SubBytesIns_Inst_Sbox_6_T13,
         SubBytesIns_Inst_Sbox_6_T12, SubBytesIns_Inst_Sbox_6_T11,
         SubBytesIns_Inst_Sbox_6_T10, SubBytesIns_Inst_Sbox_6_T9,
         SubBytesIns_Inst_Sbox_6_T8, SubBytesIns_Inst_Sbox_6_T7,
         SubBytesIns_Inst_Sbox_6_T6, SubBytesIns_Inst_Sbox_6_T5,
         SubBytesIns_Inst_Sbox_6_T4, SubBytesIns_Inst_Sbox_6_T3,
         SubBytesIns_Inst_Sbox_6_T2, SubBytesIns_Inst_Sbox_6_T1,
         SubBytesIns_Inst_Sbox_7_L29, SubBytesIns_Inst_Sbox_7_L28,
         SubBytesIns_Inst_Sbox_7_L27, SubBytesIns_Inst_Sbox_7_L26,
         SubBytesIns_Inst_Sbox_7_L25, SubBytesIns_Inst_Sbox_7_L24,
         SubBytesIns_Inst_Sbox_7_L23, SubBytesIns_Inst_Sbox_7_L22,
         SubBytesIns_Inst_Sbox_7_L21, SubBytesIns_Inst_Sbox_7_L20,
         SubBytesIns_Inst_Sbox_7_L19, SubBytesIns_Inst_Sbox_7_L18,
         SubBytesIns_Inst_Sbox_7_L17, SubBytesIns_Inst_Sbox_7_L16,
         SubBytesIns_Inst_Sbox_7_L15, SubBytesIns_Inst_Sbox_7_L14,
         SubBytesIns_Inst_Sbox_7_L13, SubBytesIns_Inst_Sbox_7_L12,
         SubBytesIns_Inst_Sbox_7_L11, SubBytesIns_Inst_Sbox_7_L10,
         SubBytesIns_Inst_Sbox_7_L9, SubBytesIns_Inst_Sbox_7_L8,
         SubBytesIns_Inst_Sbox_7_L7, SubBytesIns_Inst_Sbox_7_L6,
         SubBytesIns_Inst_Sbox_7_L5, SubBytesIns_Inst_Sbox_7_L4,
         SubBytesIns_Inst_Sbox_7_L3, SubBytesIns_Inst_Sbox_7_L2,
         SubBytesIns_Inst_Sbox_7_L1, SubBytesIns_Inst_Sbox_7_L0,
         SubBytesIns_Inst_Sbox_7_M63, SubBytesIns_Inst_Sbox_7_M62,
         SubBytesIns_Inst_Sbox_7_M61, SubBytesIns_Inst_Sbox_7_M60,
         SubBytesIns_Inst_Sbox_7_M59, SubBytesIns_Inst_Sbox_7_M58,
         SubBytesIns_Inst_Sbox_7_M57, SubBytesIns_Inst_Sbox_7_M56,
         SubBytesIns_Inst_Sbox_7_M55, SubBytesIns_Inst_Sbox_7_M54,
         SubBytesIns_Inst_Sbox_7_M53, SubBytesIns_Inst_Sbox_7_M52,
         SubBytesIns_Inst_Sbox_7_M51, SubBytesIns_Inst_Sbox_7_M50,
         SubBytesIns_Inst_Sbox_7_M49, SubBytesIns_Inst_Sbox_7_M48,
         SubBytesIns_Inst_Sbox_7_M47, SubBytesIns_Inst_Sbox_7_M46,
         SubBytesIns_Inst_Sbox_7_M45, SubBytesIns_Inst_Sbox_7_M44,
         SubBytesIns_Inst_Sbox_7_M43, SubBytesIns_Inst_Sbox_7_M42,
         SubBytesIns_Inst_Sbox_7_M41, SubBytesIns_Inst_Sbox_7_M40,
         SubBytesIns_Inst_Sbox_7_M39, SubBytesIns_Inst_Sbox_7_M38,
         SubBytesIns_Inst_Sbox_7_M37, SubBytesIns_Inst_Sbox_7_M36,
         SubBytesIns_Inst_Sbox_7_M35, SubBytesIns_Inst_Sbox_7_M34,
         SubBytesIns_Inst_Sbox_7_M33, SubBytesIns_Inst_Sbox_7_M32,
         SubBytesIns_Inst_Sbox_7_M31, SubBytesIns_Inst_Sbox_7_M30,
         SubBytesIns_Inst_Sbox_7_M29, SubBytesIns_Inst_Sbox_7_M28,
         SubBytesIns_Inst_Sbox_7_M27, SubBytesIns_Inst_Sbox_7_M26,
         SubBytesIns_Inst_Sbox_7_M25, SubBytesIns_Inst_Sbox_7_M24,
         SubBytesIns_Inst_Sbox_7_M23, SubBytesIns_Inst_Sbox_7_M22,
         SubBytesIns_Inst_Sbox_7_M21, SubBytesIns_Inst_Sbox_7_M20,
         SubBytesIns_Inst_Sbox_7_M19, SubBytesIns_Inst_Sbox_7_M18,
         SubBytesIns_Inst_Sbox_7_M17, SubBytesIns_Inst_Sbox_7_M16,
         SubBytesIns_Inst_Sbox_7_M15, SubBytesIns_Inst_Sbox_7_M14,
         SubBytesIns_Inst_Sbox_7_M13, SubBytesIns_Inst_Sbox_7_M12,
         SubBytesIns_Inst_Sbox_7_M11, SubBytesIns_Inst_Sbox_7_M10,
         SubBytesIns_Inst_Sbox_7_M9, SubBytesIns_Inst_Sbox_7_M8,
         SubBytesIns_Inst_Sbox_7_M7, SubBytesIns_Inst_Sbox_7_M6,
         SubBytesIns_Inst_Sbox_7_M5, SubBytesIns_Inst_Sbox_7_M4,
         SubBytesIns_Inst_Sbox_7_M3, SubBytesIns_Inst_Sbox_7_M2,
         SubBytesIns_Inst_Sbox_7_M1, SubBytesIns_Inst_Sbox_7_T27,
         SubBytesIns_Inst_Sbox_7_T26, SubBytesIns_Inst_Sbox_7_T25,
         SubBytesIns_Inst_Sbox_7_T24, SubBytesIns_Inst_Sbox_7_T23,
         SubBytesIns_Inst_Sbox_7_T22, SubBytesIns_Inst_Sbox_7_T21,
         SubBytesIns_Inst_Sbox_7_T20, SubBytesIns_Inst_Sbox_7_T19,
         SubBytesIns_Inst_Sbox_7_T18, SubBytesIns_Inst_Sbox_7_T17,
         SubBytesIns_Inst_Sbox_7_T16, SubBytesIns_Inst_Sbox_7_T15,
         SubBytesIns_Inst_Sbox_7_T14, SubBytesIns_Inst_Sbox_7_T13,
         SubBytesIns_Inst_Sbox_7_T12, SubBytesIns_Inst_Sbox_7_T11,
         SubBytesIns_Inst_Sbox_7_T10, SubBytesIns_Inst_Sbox_7_T9,
         SubBytesIns_Inst_Sbox_7_T8, SubBytesIns_Inst_Sbox_7_T7,
         SubBytesIns_Inst_Sbox_7_T6, SubBytesIns_Inst_Sbox_7_T5,
         SubBytesIns_Inst_Sbox_7_T4, SubBytesIns_Inst_Sbox_7_T3,
         SubBytesIns_Inst_Sbox_7_T2, SubBytesIns_Inst_Sbox_7_T1,
         SubBytesIns_Inst_Sbox_8_L29, SubBytesIns_Inst_Sbox_8_L28,
         SubBytesIns_Inst_Sbox_8_L27, SubBytesIns_Inst_Sbox_8_L26,
         SubBytesIns_Inst_Sbox_8_L25, SubBytesIns_Inst_Sbox_8_L24,
         SubBytesIns_Inst_Sbox_8_L23, SubBytesIns_Inst_Sbox_8_L22,
         SubBytesIns_Inst_Sbox_8_L21, SubBytesIns_Inst_Sbox_8_L20,
         SubBytesIns_Inst_Sbox_8_L19, SubBytesIns_Inst_Sbox_8_L18,
         SubBytesIns_Inst_Sbox_8_L17, SubBytesIns_Inst_Sbox_8_L16,
         SubBytesIns_Inst_Sbox_8_L15, SubBytesIns_Inst_Sbox_8_L14,
         SubBytesIns_Inst_Sbox_8_L13, SubBytesIns_Inst_Sbox_8_L12,
         SubBytesIns_Inst_Sbox_8_L11, SubBytesIns_Inst_Sbox_8_L10,
         SubBytesIns_Inst_Sbox_8_L9, SubBytesIns_Inst_Sbox_8_L8,
         SubBytesIns_Inst_Sbox_8_L7, SubBytesIns_Inst_Sbox_8_L6,
         SubBytesIns_Inst_Sbox_8_L5, SubBytesIns_Inst_Sbox_8_L4,
         SubBytesIns_Inst_Sbox_8_L3, SubBytesIns_Inst_Sbox_8_L2,
         SubBytesIns_Inst_Sbox_8_L1, SubBytesIns_Inst_Sbox_8_L0,
         SubBytesIns_Inst_Sbox_8_M63, SubBytesIns_Inst_Sbox_8_M62,
         SubBytesIns_Inst_Sbox_8_M61, SubBytesIns_Inst_Sbox_8_M60,
         SubBytesIns_Inst_Sbox_8_M59, SubBytesIns_Inst_Sbox_8_M58,
         SubBytesIns_Inst_Sbox_8_M57, SubBytesIns_Inst_Sbox_8_M56,
         SubBytesIns_Inst_Sbox_8_M55, SubBytesIns_Inst_Sbox_8_M54,
         SubBytesIns_Inst_Sbox_8_M53, SubBytesIns_Inst_Sbox_8_M52,
         SubBytesIns_Inst_Sbox_8_M51, SubBytesIns_Inst_Sbox_8_M50,
         SubBytesIns_Inst_Sbox_8_M49, SubBytesIns_Inst_Sbox_8_M48,
         SubBytesIns_Inst_Sbox_8_M47, SubBytesIns_Inst_Sbox_8_M46,
         SubBytesIns_Inst_Sbox_8_M45, SubBytesIns_Inst_Sbox_8_M44,
         SubBytesIns_Inst_Sbox_8_M43, SubBytesIns_Inst_Sbox_8_M42,
         SubBytesIns_Inst_Sbox_8_M41, SubBytesIns_Inst_Sbox_8_M40,
         SubBytesIns_Inst_Sbox_8_M39, SubBytesIns_Inst_Sbox_8_M38,
         SubBytesIns_Inst_Sbox_8_M37, SubBytesIns_Inst_Sbox_8_M36,
         SubBytesIns_Inst_Sbox_8_M35, SubBytesIns_Inst_Sbox_8_M34,
         SubBytesIns_Inst_Sbox_8_M33, SubBytesIns_Inst_Sbox_8_M32,
         SubBytesIns_Inst_Sbox_8_M31, SubBytesIns_Inst_Sbox_8_M30,
         SubBytesIns_Inst_Sbox_8_M29, SubBytesIns_Inst_Sbox_8_M28,
         SubBytesIns_Inst_Sbox_8_M27, SubBytesIns_Inst_Sbox_8_M26,
         SubBytesIns_Inst_Sbox_8_M25, SubBytesIns_Inst_Sbox_8_M24,
         SubBytesIns_Inst_Sbox_8_M23, SubBytesIns_Inst_Sbox_8_M22,
         SubBytesIns_Inst_Sbox_8_M21, SubBytesIns_Inst_Sbox_8_M20,
         SubBytesIns_Inst_Sbox_8_M19, SubBytesIns_Inst_Sbox_8_M18,
         SubBytesIns_Inst_Sbox_8_M17, SubBytesIns_Inst_Sbox_8_M16,
         SubBytesIns_Inst_Sbox_8_M15, SubBytesIns_Inst_Sbox_8_M14,
         SubBytesIns_Inst_Sbox_8_M13, SubBytesIns_Inst_Sbox_8_M12,
         SubBytesIns_Inst_Sbox_8_M11, SubBytesIns_Inst_Sbox_8_M10,
         SubBytesIns_Inst_Sbox_8_M9, SubBytesIns_Inst_Sbox_8_M8,
         SubBytesIns_Inst_Sbox_8_M7, SubBytesIns_Inst_Sbox_8_M6,
         SubBytesIns_Inst_Sbox_8_M5, SubBytesIns_Inst_Sbox_8_M4,
         SubBytesIns_Inst_Sbox_8_M3, SubBytesIns_Inst_Sbox_8_M2,
         SubBytesIns_Inst_Sbox_8_M1, SubBytesIns_Inst_Sbox_8_T27,
         SubBytesIns_Inst_Sbox_8_T26, SubBytesIns_Inst_Sbox_8_T25,
         SubBytesIns_Inst_Sbox_8_T24, SubBytesIns_Inst_Sbox_8_T23,
         SubBytesIns_Inst_Sbox_8_T22, SubBytesIns_Inst_Sbox_8_T21,
         SubBytesIns_Inst_Sbox_8_T20, SubBytesIns_Inst_Sbox_8_T19,
         SubBytesIns_Inst_Sbox_8_T18, SubBytesIns_Inst_Sbox_8_T17,
         SubBytesIns_Inst_Sbox_8_T16, SubBytesIns_Inst_Sbox_8_T15,
         SubBytesIns_Inst_Sbox_8_T14, SubBytesIns_Inst_Sbox_8_T13,
         SubBytesIns_Inst_Sbox_8_T12, SubBytesIns_Inst_Sbox_8_T11,
         SubBytesIns_Inst_Sbox_8_T10, SubBytesIns_Inst_Sbox_8_T9,
         SubBytesIns_Inst_Sbox_8_T8, SubBytesIns_Inst_Sbox_8_T7,
         SubBytesIns_Inst_Sbox_8_T6, SubBytesIns_Inst_Sbox_8_T5,
         SubBytesIns_Inst_Sbox_8_T4, SubBytesIns_Inst_Sbox_8_T3,
         SubBytesIns_Inst_Sbox_8_T2, SubBytesIns_Inst_Sbox_8_T1,
         SubBytesIns_Inst_Sbox_9_L29, SubBytesIns_Inst_Sbox_9_L28,
         SubBytesIns_Inst_Sbox_9_L27, SubBytesIns_Inst_Sbox_9_L26,
         SubBytesIns_Inst_Sbox_9_L25, SubBytesIns_Inst_Sbox_9_L24,
         SubBytesIns_Inst_Sbox_9_L23, SubBytesIns_Inst_Sbox_9_L22,
         SubBytesIns_Inst_Sbox_9_L21, SubBytesIns_Inst_Sbox_9_L20,
         SubBytesIns_Inst_Sbox_9_L19, SubBytesIns_Inst_Sbox_9_L18,
         SubBytesIns_Inst_Sbox_9_L17, SubBytesIns_Inst_Sbox_9_L16,
         SubBytesIns_Inst_Sbox_9_L15, SubBytesIns_Inst_Sbox_9_L14,
         SubBytesIns_Inst_Sbox_9_L13, SubBytesIns_Inst_Sbox_9_L12,
         SubBytesIns_Inst_Sbox_9_L11, SubBytesIns_Inst_Sbox_9_L10,
         SubBytesIns_Inst_Sbox_9_L9, SubBytesIns_Inst_Sbox_9_L8,
         SubBytesIns_Inst_Sbox_9_L7, SubBytesIns_Inst_Sbox_9_L6,
         SubBytesIns_Inst_Sbox_9_L5, SubBytesIns_Inst_Sbox_9_L4,
         SubBytesIns_Inst_Sbox_9_L3, SubBytesIns_Inst_Sbox_9_L2,
         SubBytesIns_Inst_Sbox_9_L1, SubBytesIns_Inst_Sbox_9_L0,
         SubBytesIns_Inst_Sbox_9_M63, SubBytesIns_Inst_Sbox_9_M62,
         SubBytesIns_Inst_Sbox_9_M61, SubBytesIns_Inst_Sbox_9_M60,
         SubBytesIns_Inst_Sbox_9_M59, SubBytesIns_Inst_Sbox_9_M58,
         SubBytesIns_Inst_Sbox_9_M57, SubBytesIns_Inst_Sbox_9_M56,
         SubBytesIns_Inst_Sbox_9_M55, SubBytesIns_Inst_Sbox_9_M54,
         SubBytesIns_Inst_Sbox_9_M53, SubBytesIns_Inst_Sbox_9_M52,
         SubBytesIns_Inst_Sbox_9_M51, SubBytesIns_Inst_Sbox_9_M50,
         SubBytesIns_Inst_Sbox_9_M49, SubBytesIns_Inst_Sbox_9_M48,
         SubBytesIns_Inst_Sbox_9_M47, SubBytesIns_Inst_Sbox_9_M46,
         SubBytesIns_Inst_Sbox_9_M45, SubBytesIns_Inst_Sbox_9_M44,
         SubBytesIns_Inst_Sbox_9_M43, SubBytesIns_Inst_Sbox_9_M42,
         SubBytesIns_Inst_Sbox_9_M41, SubBytesIns_Inst_Sbox_9_M40,
         SubBytesIns_Inst_Sbox_9_M39, SubBytesIns_Inst_Sbox_9_M38,
         SubBytesIns_Inst_Sbox_9_M37, SubBytesIns_Inst_Sbox_9_M36,
         SubBytesIns_Inst_Sbox_9_M35, SubBytesIns_Inst_Sbox_9_M34,
         SubBytesIns_Inst_Sbox_9_M33, SubBytesIns_Inst_Sbox_9_M32,
         SubBytesIns_Inst_Sbox_9_M31, SubBytesIns_Inst_Sbox_9_M30,
         SubBytesIns_Inst_Sbox_9_M29, SubBytesIns_Inst_Sbox_9_M28,
         SubBytesIns_Inst_Sbox_9_M27, SubBytesIns_Inst_Sbox_9_M26,
         SubBytesIns_Inst_Sbox_9_M25, SubBytesIns_Inst_Sbox_9_M24,
         SubBytesIns_Inst_Sbox_9_M23, SubBytesIns_Inst_Sbox_9_M22,
         SubBytesIns_Inst_Sbox_9_M21, SubBytesIns_Inst_Sbox_9_M20,
         SubBytesIns_Inst_Sbox_9_M19, SubBytesIns_Inst_Sbox_9_M18,
         SubBytesIns_Inst_Sbox_9_M17, SubBytesIns_Inst_Sbox_9_M16,
         SubBytesIns_Inst_Sbox_9_M15, SubBytesIns_Inst_Sbox_9_M14,
         SubBytesIns_Inst_Sbox_9_M13, SubBytesIns_Inst_Sbox_9_M12,
         SubBytesIns_Inst_Sbox_9_M11, SubBytesIns_Inst_Sbox_9_M10,
         SubBytesIns_Inst_Sbox_9_M9, SubBytesIns_Inst_Sbox_9_M8,
         SubBytesIns_Inst_Sbox_9_M7, SubBytesIns_Inst_Sbox_9_M6,
         SubBytesIns_Inst_Sbox_9_M5, SubBytesIns_Inst_Sbox_9_M4,
         SubBytesIns_Inst_Sbox_9_M3, SubBytesIns_Inst_Sbox_9_M2,
         SubBytesIns_Inst_Sbox_9_M1, SubBytesIns_Inst_Sbox_9_T27,
         SubBytesIns_Inst_Sbox_9_T26, SubBytesIns_Inst_Sbox_9_T25,
         SubBytesIns_Inst_Sbox_9_T24, SubBytesIns_Inst_Sbox_9_T23,
         SubBytesIns_Inst_Sbox_9_T22, SubBytesIns_Inst_Sbox_9_T21,
         SubBytesIns_Inst_Sbox_9_T20, SubBytesIns_Inst_Sbox_9_T19,
         SubBytesIns_Inst_Sbox_9_T18, SubBytesIns_Inst_Sbox_9_T17,
         SubBytesIns_Inst_Sbox_9_T16, SubBytesIns_Inst_Sbox_9_T15,
         SubBytesIns_Inst_Sbox_9_T14, SubBytesIns_Inst_Sbox_9_T13,
         SubBytesIns_Inst_Sbox_9_T12, SubBytesIns_Inst_Sbox_9_T11,
         SubBytesIns_Inst_Sbox_9_T10, SubBytesIns_Inst_Sbox_9_T9,
         SubBytesIns_Inst_Sbox_9_T8, SubBytesIns_Inst_Sbox_9_T7,
         SubBytesIns_Inst_Sbox_9_T6, SubBytesIns_Inst_Sbox_9_T5,
         SubBytesIns_Inst_Sbox_9_T4, SubBytesIns_Inst_Sbox_9_T3,
         SubBytesIns_Inst_Sbox_9_T2, SubBytesIns_Inst_Sbox_9_T1,
         SubBytesIns_Inst_Sbox_10_L29, SubBytesIns_Inst_Sbox_10_L28,
         SubBytesIns_Inst_Sbox_10_L27, SubBytesIns_Inst_Sbox_10_L26,
         SubBytesIns_Inst_Sbox_10_L25, SubBytesIns_Inst_Sbox_10_L24,
         SubBytesIns_Inst_Sbox_10_L23, SubBytesIns_Inst_Sbox_10_L22,
         SubBytesIns_Inst_Sbox_10_L21, SubBytesIns_Inst_Sbox_10_L20,
         SubBytesIns_Inst_Sbox_10_L19, SubBytesIns_Inst_Sbox_10_L18,
         SubBytesIns_Inst_Sbox_10_L17, SubBytesIns_Inst_Sbox_10_L16,
         SubBytesIns_Inst_Sbox_10_L15, SubBytesIns_Inst_Sbox_10_L14,
         SubBytesIns_Inst_Sbox_10_L13, SubBytesIns_Inst_Sbox_10_L12,
         SubBytesIns_Inst_Sbox_10_L11, SubBytesIns_Inst_Sbox_10_L10,
         SubBytesIns_Inst_Sbox_10_L9, SubBytesIns_Inst_Sbox_10_L8,
         SubBytesIns_Inst_Sbox_10_L7, SubBytesIns_Inst_Sbox_10_L6,
         SubBytesIns_Inst_Sbox_10_L5, SubBytesIns_Inst_Sbox_10_L4,
         SubBytesIns_Inst_Sbox_10_L3, SubBytesIns_Inst_Sbox_10_L2,
         SubBytesIns_Inst_Sbox_10_L1, SubBytesIns_Inst_Sbox_10_L0,
         SubBytesIns_Inst_Sbox_10_M63, SubBytesIns_Inst_Sbox_10_M62,
         SubBytesIns_Inst_Sbox_10_M61, SubBytesIns_Inst_Sbox_10_M60,
         SubBytesIns_Inst_Sbox_10_M59, SubBytesIns_Inst_Sbox_10_M58,
         SubBytesIns_Inst_Sbox_10_M57, SubBytesIns_Inst_Sbox_10_M56,
         SubBytesIns_Inst_Sbox_10_M55, SubBytesIns_Inst_Sbox_10_M54,
         SubBytesIns_Inst_Sbox_10_M53, SubBytesIns_Inst_Sbox_10_M52,
         SubBytesIns_Inst_Sbox_10_M51, SubBytesIns_Inst_Sbox_10_M50,
         SubBytesIns_Inst_Sbox_10_M49, SubBytesIns_Inst_Sbox_10_M48,
         SubBytesIns_Inst_Sbox_10_M47, SubBytesIns_Inst_Sbox_10_M46,
         SubBytesIns_Inst_Sbox_10_M45, SubBytesIns_Inst_Sbox_10_M44,
         SubBytesIns_Inst_Sbox_10_M43, SubBytesIns_Inst_Sbox_10_M42,
         SubBytesIns_Inst_Sbox_10_M41, SubBytesIns_Inst_Sbox_10_M40,
         SubBytesIns_Inst_Sbox_10_M39, SubBytesIns_Inst_Sbox_10_M38,
         SubBytesIns_Inst_Sbox_10_M37, SubBytesIns_Inst_Sbox_10_M36,
         SubBytesIns_Inst_Sbox_10_M35, SubBytesIns_Inst_Sbox_10_M34,
         SubBytesIns_Inst_Sbox_10_M33, SubBytesIns_Inst_Sbox_10_M32,
         SubBytesIns_Inst_Sbox_10_M31, SubBytesIns_Inst_Sbox_10_M30,
         SubBytesIns_Inst_Sbox_10_M29, SubBytesIns_Inst_Sbox_10_M28,
         SubBytesIns_Inst_Sbox_10_M27, SubBytesIns_Inst_Sbox_10_M26,
         SubBytesIns_Inst_Sbox_10_M25, SubBytesIns_Inst_Sbox_10_M24,
         SubBytesIns_Inst_Sbox_10_M23, SubBytesIns_Inst_Sbox_10_M22,
         SubBytesIns_Inst_Sbox_10_M21, SubBytesIns_Inst_Sbox_10_M20,
         SubBytesIns_Inst_Sbox_10_M19, SubBytesIns_Inst_Sbox_10_M18,
         SubBytesIns_Inst_Sbox_10_M17, SubBytesIns_Inst_Sbox_10_M16,
         SubBytesIns_Inst_Sbox_10_M15, SubBytesIns_Inst_Sbox_10_M14,
         SubBytesIns_Inst_Sbox_10_M13, SubBytesIns_Inst_Sbox_10_M12,
         SubBytesIns_Inst_Sbox_10_M11, SubBytesIns_Inst_Sbox_10_M10,
         SubBytesIns_Inst_Sbox_10_M9, SubBytesIns_Inst_Sbox_10_M8,
         SubBytesIns_Inst_Sbox_10_M7, SubBytesIns_Inst_Sbox_10_M6,
         SubBytesIns_Inst_Sbox_10_M5, SubBytesIns_Inst_Sbox_10_M4,
         SubBytesIns_Inst_Sbox_10_M3, SubBytesIns_Inst_Sbox_10_M2,
         SubBytesIns_Inst_Sbox_10_M1, SubBytesIns_Inst_Sbox_10_T27,
         SubBytesIns_Inst_Sbox_10_T26, SubBytesIns_Inst_Sbox_10_T25,
         SubBytesIns_Inst_Sbox_10_T24, SubBytesIns_Inst_Sbox_10_T23,
         SubBytesIns_Inst_Sbox_10_T22, SubBytesIns_Inst_Sbox_10_T21,
         SubBytesIns_Inst_Sbox_10_T20, SubBytesIns_Inst_Sbox_10_T19,
         SubBytesIns_Inst_Sbox_10_T18, SubBytesIns_Inst_Sbox_10_T17,
         SubBytesIns_Inst_Sbox_10_T16, SubBytesIns_Inst_Sbox_10_T15,
         SubBytesIns_Inst_Sbox_10_T14, SubBytesIns_Inst_Sbox_10_T13,
         SubBytesIns_Inst_Sbox_10_T12, SubBytesIns_Inst_Sbox_10_T11,
         SubBytesIns_Inst_Sbox_10_T10, SubBytesIns_Inst_Sbox_10_T9,
         SubBytesIns_Inst_Sbox_10_T8, SubBytesIns_Inst_Sbox_10_T7,
         SubBytesIns_Inst_Sbox_10_T6, SubBytesIns_Inst_Sbox_10_T5,
         SubBytesIns_Inst_Sbox_10_T4, SubBytesIns_Inst_Sbox_10_T3,
         SubBytesIns_Inst_Sbox_10_T2, SubBytesIns_Inst_Sbox_10_T1,
         SubBytesIns_Inst_Sbox_11_L29, SubBytesIns_Inst_Sbox_11_L28,
         SubBytesIns_Inst_Sbox_11_L27, SubBytesIns_Inst_Sbox_11_L26,
         SubBytesIns_Inst_Sbox_11_L25, SubBytesIns_Inst_Sbox_11_L24,
         SubBytesIns_Inst_Sbox_11_L23, SubBytesIns_Inst_Sbox_11_L22,
         SubBytesIns_Inst_Sbox_11_L21, SubBytesIns_Inst_Sbox_11_L20,
         SubBytesIns_Inst_Sbox_11_L19, SubBytesIns_Inst_Sbox_11_L18,
         SubBytesIns_Inst_Sbox_11_L17, SubBytesIns_Inst_Sbox_11_L16,
         SubBytesIns_Inst_Sbox_11_L15, SubBytesIns_Inst_Sbox_11_L14,
         SubBytesIns_Inst_Sbox_11_L13, SubBytesIns_Inst_Sbox_11_L12,
         SubBytesIns_Inst_Sbox_11_L11, SubBytesIns_Inst_Sbox_11_L10,
         SubBytesIns_Inst_Sbox_11_L9, SubBytesIns_Inst_Sbox_11_L8,
         SubBytesIns_Inst_Sbox_11_L7, SubBytesIns_Inst_Sbox_11_L6,
         SubBytesIns_Inst_Sbox_11_L5, SubBytesIns_Inst_Sbox_11_L4,
         SubBytesIns_Inst_Sbox_11_L3, SubBytesIns_Inst_Sbox_11_L2,
         SubBytesIns_Inst_Sbox_11_L1, SubBytesIns_Inst_Sbox_11_L0,
         SubBytesIns_Inst_Sbox_11_M63, SubBytesIns_Inst_Sbox_11_M62,
         SubBytesIns_Inst_Sbox_11_M61, SubBytesIns_Inst_Sbox_11_M60,
         SubBytesIns_Inst_Sbox_11_M59, SubBytesIns_Inst_Sbox_11_M58,
         SubBytesIns_Inst_Sbox_11_M57, SubBytesIns_Inst_Sbox_11_M56,
         SubBytesIns_Inst_Sbox_11_M55, SubBytesIns_Inst_Sbox_11_M54,
         SubBytesIns_Inst_Sbox_11_M53, SubBytesIns_Inst_Sbox_11_M52,
         SubBytesIns_Inst_Sbox_11_M51, SubBytesIns_Inst_Sbox_11_M50,
         SubBytesIns_Inst_Sbox_11_M49, SubBytesIns_Inst_Sbox_11_M48,
         SubBytesIns_Inst_Sbox_11_M47, SubBytesIns_Inst_Sbox_11_M46,
         SubBytesIns_Inst_Sbox_11_M45, SubBytesIns_Inst_Sbox_11_M44,
         SubBytesIns_Inst_Sbox_11_M43, SubBytesIns_Inst_Sbox_11_M42,
         SubBytesIns_Inst_Sbox_11_M41, SubBytesIns_Inst_Sbox_11_M40,
         SubBytesIns_Inst_Sbox_11_M39, SubBytesIns_Inst_Sbox_11_M38,
         SubBytesIns_Inst_Sbox_11_M37, SubBytesIns_Inst_Sbox_11_M36,
         SubBytesIns_Inst_Sbox_11_M35, SubBytesIns_Inst_Sbox_11_M34,
         SubBytesIns_Inst_Sbox_11_M33, SubBytesIns_Inst_Sbox_11_M32,
         SubBytesIns_Inst_Sbox_11_M31, SubBytesIns_Inst_Sbox_11_M30,
         SubBytesIns_Inst_Sbox_11_M29, SubBytesIns_Inst_Sbox_11_M28,
         SubBytesIns_Inst_Sbox_11_M27, SubBytesIns_Inst_Sbox_11_M26,
         SubBytesIns_Inst_Sbox_11_M25, SubBytesIns_Inst_Sbox_11_M24,
         SubBytesIns_Inst_Sbox_11_M23, SubBytesIns_Inst_Sbox_11_M22,
         SubBytesIns_Inst_Sbox_11_M21, SubBytesIns_Inst_Sbox_11_M20,
         SubBytesIns_Inst_Sbox_11_M19, SubBytesIns_Inst_Sbox_11_M18,
         SubBytesIns_Inst_Sbox_11_M17, SubBytesIns_Inst_Sbox_11_M16,
         SubBytesIns_Inst_Sbox_11_M15, SubBytesIns_Inst_Sbox_11_M14,
         SubBytesIns_Inst_Sbox_11_M13, SubBytesIns_Inst_Sbox_11_M12,
         SubBytesIns_Inst_Sbox_11_M11, SubBytesIns_Inst_Sbox_11_M10,
         SubBytesIns_Inst_Sbox_11_M9, SubBytesIns_Inst_Sbox_11_M8,
         SubBytesIns_Inst_Sbox_11_M7, SubBytesIns_Inst_Sbox_11_M6,
         SubBytesIns_Inst_Sbox_11_M5, SubBytesIns_Inst_Sbox_11_M4,
         SubBytesIns_Inst_Sbox_11_M3, SubBytesIns_Inst_Sbox_11_M2,
         SubBytesIns_Inst_Sbox_11_M1, SubBytesIns_Inst_Sbox_11_T27,
         SubBytesIns_Inst_Sbox_11_T26, SubBytesIns_Inst_Sbox_11_T25,
         SubBytesIns_Inst_Sbox_11_T24, SubBytesIns_Inst_Sbox_11_T23,
         SubBytesIns_Inst_Sbox_11_T22, SubBytesIns_Inst_Sbox_11_T21,
         SubBytesIns_Inst_Sbox_11_T20, SubBytesIns_Inst_Sbox_11_T19,
         SubBytesIns_Inst_Sbox_11_T18, SubBytesIns_Inst_Sbox_11_T17,
         SubBytesIns_Inst_Sbox_11_T16, SubBytesIns_Inst_Sbox_11_T15,
         SubBytesIns_Inst_Sbox_11_T14, SubBytesIns_Inst_Sbox_11_T13,
         SubBytesIns_Inst_Sbox_11_T12, SubBytesIns_Inst_Sbox_11_T11,
         SubBytesIns_Inst_Sbox_11_T10, SubBytesIns_Inst_Sbox_11_T9,
         SubBytesIns_Inst_Sbox_11_T8, SubBytesIns_Inst_Sbox_11_T7,
         SubBytesIns_Inst_Sbox_11_T6, SubBytesIns_Inst_Sbox_11_T5,
         SubBytesIns_Inst_Sbox_11_T4, SubBytesIns_Inst_Sbox_11_T3,
         SubBytesIns_Inst_Sbox_11_T2, SubBytesIns_Inst_Sbox_11_T1,
         SubBytesIns_Inst_Sbox_12_L29, SubBytesIns_Inst_Sbox_12_L28,
         SubBytesIns_Inst_Sbox_12_L27, SubBytesIns_Inst_Sbox_12_L26,
         SubBytesIns_Inst_Sbox_12_L25, SubBytesIns_Inst_Sbox_12_L24,
         SubBytesIns_Inst_Sbox_12_L23, SubBytesIns_Inst_Sbox_12_L22,
         SubBytesIns_Inst_Sbox_12_L21, SubBytesIns_Inst_Sbox_12_L20,
         SubBytesIns_Inst_Sbox_12_L19, SubBytesIns_Inst_Sbox_12_L18,
         SubBytesIns_Inst_Sbox_12_L17, SubBytesIns_Inst_Sbox_12_L16,
         SubBytesIns_Inst_Sbox_12_L15, SubBytesIns_Inst_Sbox_12_L14,
         SubBytesIns_Inst_Sbox_12_L13, SubBytesIns_Inst_Sbox_12_L12,
         SubBytesIns_Inst_Sbox_12_L11, SubBytesIns_Inst_Sbox_12_L10,
         SubBytesIns_Inst_Sbox_12_L9, SubBytesIns_Inst_Sbox_12_L8,
         SubBytesIns_Inst_Sbox_12_L7, SubBytesIns_Inst_Sbox_12_L6,
         SubBytesIns_Inst_Sbox_12_L5, SubBytesIns_Inst_Sbox_12_L4,
         SubBytesIns_Inst_Sbox_12_L3, SubBytesIns_Inst_Sbox_12_L2,
         SubBytesIns_Inst_Sbox_12_L1, SubBytesIns_Inst_Sbox_12_L0,
         SubBytesIns_Inst_Sbox_12_M63, SubBytesIns_Inst_Sbox_12_M62,
         SubBytesIns_Inst_Sbox_12_M61, SubBytesIns_Inst_Sbox_12_M60,
         SubBytesIns_Inst_Sbox_12_M59, SubBytesIns_Inst_Sbox_12_M58,
         SubBytesIns_Inst_Sbox_12_M57, SubBytesIns_Inst_Sbox_12_M56,
         SubBytesIns_Inst_Sbox_12_M55, SubBytesIns_Inst_Sbox_12_M54,
         SubBytesIns_Inst_Sbox_12_M53, SubBytesIns_Inst_Sbox_12_M52,
         SubBytesIns_Inst_Sbox_12_M51, SubBytesIns_Inst_Sbox_12_M50,
         SubBytesIns_Inst_Sbox_12_M49, SubBytesIns_Inst_Sbox_12_M48,
         SubBytesIns_Inst_Sbox_12_M47, SubBytesIns_Inst_Sbox_12_M46,
         SubBytesIns_Inst_Sbox_12_M45, SubBytesIns_Inst_Sbox_12_M44,
         SubBytesIns_Inst_Sbox_12_M43, SubBytesIns_Inst_Sbox_12_M42,
         SubBytesIns_Inst_Sbox_12_M41, SubBytesIns_Inst_Sbox_12_M40,
         SubBytesIns_Inst_Sbox_12_M39, SubBytesIns_Inst_Sbox_12_M38,
         SubBytesIns_Inst_Sbox_12_M37, SubBytesIns_Inst_Sbox_12_M36,
         SubBytesIns_Inst_Sbox_12_M35, SubBytesIns_Inst_Sbox_12_M34,
         SubBytesIns_Inst_Sbox_12_M33, SubBytesIns_Inst_Sbox_12_M32,
         SubBytesIns_Inst_Sbox_12_M31, SubBytesIns_Inst_Sbox_12_M30,
         SubBytesIns_Inst_Sbox_12_M29, SubBytesIns_Inst_Sbox_12_M28,
         SubBytesIns_Inst_Sbox_12_M27, SubBytesIns_Inst_Sbox_12_M26,
         SubBytesIns_Inst_Sbox_12_M25, SubBytesIns_Inst_Sbox_12_M24,
         SubBytesIns_Inst_Sbox_12_M23, SubBytesIns_Inst_Sbox_12_M22,
         SubBytesIns_Inst_Sbox_12_M21, SubBytesIns_Inst_Sbox_12_M20,
         SubBytesIns_Inst_Sbox_12_M19, SubBytesIns_Inst_Sbox_12_M18,
         SubBytesIns_Inst_Sbox_12_M17, SubBytesIns_Inst_Sbox_12_M16,
         SubBytesIns_Inst_Sbox_12_M15, SubBytesIns_Inst_Sbox_12_M14,
         SubBytesIns_Inst_Sbox_12_M13, SubBytesIns_Inst_Sbox_12_M12,
         SubBytesIns_Inst_Sbox_12_M11, SubBytesIns_Inst_Sbox_12_M10,
         SubBytesIns_Inst_Sbox_12_M9, SubBytesIns_Inst_Sbox_12_M8,
         SubBytesIns_Inst_Sbox_12_M7, SubBytesIns_Inst_Sbox_12_M6,
         SubBytesIns_Inst_Sbox_12_M5, SubBytesIns_Inst_Sbox_12_M4,
         SubBytesIns_Inst_Sbox_12_M3, SubBytesIns_Inst_Sbox_12_M2,
         SubBytesIns_Inst_Sbox_12_M1, SubBytesIns_Inst_Sbox_12_T27,
         SubBytesIns_Inst_Sbox_12_T26, SubBytesIns_Inst_Sbox_12_T25,
         SubBytesIns_Inst_Sbox_12_T24, SubBytesIns_Inst_Sbox_12_T23,
         SubBytesIns_Inst_Sbox_12_T22, SubBytesIns_Inst_Sbox_12_T21,
         SubBytesIns_Inst_Sbox_12_T20, SubBytesIns_Inst_Sbox_12_T19,
         SubBytesIns_Inst_Sbox_12_T18, SubBytesIns_Inst_Sbox_12_T17,
         SubBytesIns_Inst_Sbox_12_T16, SubBytesIns_Inst_Sbox_12_T15,
         SubBytesIns_Inst_Sbox_12_T14, SubBytesIns_Inst_Sbox_12_T13,
         SubBytesIns_Inst_Sbox_12_T12, SubBytesIns_Inst_Sbox_12_T11,
         SubBytesIns_Inst_Sbox_12_T10, SubBytesIns_Inst_Sbox_12_T9,
         SubBytesIns_Inst_Sbox_12_T8, SubBytesIns_Inst_Sbox_12_T7,
         SubBytesIns_Inst_Sbox_12_T6, SubBytesIns_Inst_Sbox_12_T5,
         SubBytesIns_Inst_Sbox_12_T4, SubBytesIns_Inst_Sbox_12_T3,
         SubBytesIns_Inst_Sbox_12_T2, SubBytesIns_Inst_Sbox_12_T1,
         SubBytesIns_Inst_Sbox_13_L29, SubBytesIns_Inst_Sbox_13_L28,
         SubBytesIns_Inst_Sbox_13_L27, SubBytesIns_Inst_Sbox_13_L26,
         SubBytesIns_Inst_Sbox_13_L25, SubBytesIns_Inst_Sbox_13_L24,
         SubBytesIns_Inst_Sbox_13_L23, SubBytesIns_Inst_Sbox_13_L22,
         SubBytesIns_Inst_Sbox_13_L21, SubBytesIns_Inst_Sbox_13_L20,
         SubBytesIns_Inst_Sbox_13_L19, SubBytesIns_Inst_Sbox_13_L18,
         SubBytesIns_Inst_Sbox_13_L17, SubBytesIns_Inst_Sbox_13_L16,
         SubBytesIns_Inst_Sbox_13_L15, SubBytesIns_Inst_Sbox_13_L14,
         SubBytesIns_Inst_Sbox_13_L13, SubBytesIns_Inst_Sbox_13_L12,
         SubBytesIns_Inst_Sbox_13_L11, SubBytesIns_Inst_Sbox_13_L10,
         SubBytesIns_Inst_Sbox_13_L9, SubBytesIns_Inst_Sbox_13_L8,
         SubBytesIns_Inst_Sbox_13_L7, SubBytesIns_Inst_Sbox_13_L6,
         SubBytesIns_Inst_Sbox_13_L5, SubBytesIns_Inst_Sbox_13_L4,
         SubBytesIns_Inst_Sbox_13_L3, SubBytesIns_Inst_Sbox_13_L2,
         SubBytesIns_Inst_Sbox_13_L1, SubBytesIns_Inst_Sbox_13_L0,
         SubBytesIns_Inst_Sbox_13_M63, SubBytesIns_Inst_Sbox_13_M62,
         SubBytesIns_Inst_Sbox_13_M61, SubBytesIns_Inst_Sbox_13_M60,
         SubBytesIns_Inst_Sbox_13_M59, SubBytesIns_Inst_Sbox_13_M58,
         SubBytesIns_Inst_Sbox_13_M57, SubBytesIns_Inst_Sbox_13_M56,
         SubBytesIns_Inst_Sbox_13_M55, SubBytesIns_Inst_Sbox_13_M54,
         SubBytesIns_Inst_Sbox_13_M53, SubBytesIns_Inst_Sbox_13_M52,
         SubBytesIns_Inst_Sbox_13_M51, SubBytesIns_Inst_Sbox_13_M50,
         SubBytesIns_Inst_Sbox_13_M49, SubBytesIns_Inst_Sbox_13_M48,
         SubBytesIns_Inst_Sbox_13_M47, SubBytesIns_Inst_Sbox_13_M46,
         SubBytesIns_Inst_Sbox_13_M45, SubBytesIns_Inst_Sbox_13_M44,
         SubBytesIns_Inst_Sbox_13_M43, SubBytesIns_Inst_Sbox_13_M42,
         SubBytesIns_Inst_Sbox_13_M41, SubBytesIns_Inst_Sbox_13_M40,
         SubBytesIns_Inst_Sbox_13_M39, SubBytesIns_Inst_Sbox_13_M38,
         SubBytesIns_Inst_Sbox_13_M37, SubBytesIns_Inst_Sbox_13_M36,
         SubBytesIns_Inst_Sbox_13_M35, SubBytesIns_Inst_Sbox_13_M34,
         SubBytesIns_Inst_Sbox_13_M33, SubBytesIns_Inst_Sbox_13_M32,
         SubBytesIns_Inst_Sbox_13_M31, SubBytesIns_Inst_Sbox_13_M30,
         SubBytesIns_Inst_Sbox_13_M29, SubBytesIns_Inst_Sbox_13_M28,
         SubBytesIns_Inst_Sbox_13_M27, SubBytesIns_Inst_Sbox_13_M26,
         SubBytesIns_Inst_Sbox_13_M25, SubBytesIns_Inst_Sbox_13_M24,
         SubBytesIns_Inst_Sbox_13_M23, SubBytesIns_Inst_Sbox_13_M22,
         SubBytesIns_Inst_Sbox_13_M21, SubBytesIns_Inst_Sbox_13_M20,
         SubBytesIns_Inst_Sbox_13_M19, SubBytesIns_Inst_Sbox_13_M18,
         SubBytesIns_Inst_Sbox_13_M17, SubBytesIns_Inst_Sbox_13_M16,
         SubBytesIns_Inst_Sbox_13_M15, SubBytesIns_Inst_Sbox_13_M14,
         SubBytesIns_Inst_Sbox_13_M13, SubBytesIns_Inst_Sbox_13_M12,
         SubBytesIns_Inst_Sbox_13_M11, SubBytesIns_Inst_Sbox_13_M10,
         SubBytesIns_Inst_Sbox_13_M9, SubBytesIns_Inst_Sbox_13_M8,
         SubBytesIns_Inst_Sbox_13_M7, SubBytesIns_Inst_Sbox_13_M6,
         SubBytesIns_Inst_Sbox_13_M5, SubBytesIns_Inst_Sbox_13_M4,
         SubBytesIns_Inst_Sbox_13_M3, SubBytesIns_Inst_Sbox_13_M2,
         SubBytesIns_Inst_Sbox_13_M1, SubBytesIns_Inst_Sbox_13_T27,
         SubBytesIns_Inst_Sbox_13_T26, SubBytesIns_Inst_Sbox_13_T25,
         SubBytesIns_Inst_Sbox_13_T24, SubBytesIns_Inst_Sbox_13_T23,
         SubBytesIns_Inst_Sbox_13_T22, SubBytesIns_Inst_Sbox_13_T21,
         SubBytesIns_Inst_Sbox_13_T20, SubBytesIns_Inst_Sbox_13_T19,
         SubBytesIns_Inst_Sbox_13_T18, SubBytesIns_Inst_Sbox_13_T17,
         SubBytesIns_Inst_Sbox_13_T16, SubBytesIns_Inst_Sbox_13_T15,
         SubBytesIns_Inst_Sbox_13_T14, SubBytesIns_Inst_Sbox_13_T13,
         SubBytesIns_Inst_Sbox_13_T12, SubBytesIns_Inst_Sbox_13_T11,
         SubBytesIns_Inst_Sbox_13_T10, SubBytesIns_Inst_Sbox_13_T9,
         SubBytesIns_Inst_Sbox_13_T8, SubBytesIns_Inst_Sbox_13_T7,
         SubBytesIns_Inst_Sbox_13_T6, SubBytesIns_Inst_Sbox_13_T5,
         SubBytesIns_Inst_Sbox_13_T4, SubBytesIns_Inst_Sbox_13_T3,
         SubBytesIns_Inst_Sbox_13_T2, SubBytesIns_Inst_Sbox_13_T1,
         SubBytesIns_Inst_Sbox_14_L29, SubBytesIns_Inst_Sbox_14_L28,
         SubBytesIns_Inst_Sbox_14_L27, SubBytesIns_Inst_Sbox_14_L26,
         SubBytesIns_Inst_Sbox_14_L25, SubBytesIns_Inst_Sbox_14_L24,
         SubBytesIns_Inst_Sbox_14_L23, SubBytesIns_Inst_Sbox_14_L22,
         SubBytesIns_Inst_Sbox_14_L21, SubBytesIns_Inst_Sbox_14_L20,
         SubBytesIns_Inst_Sbox_14_L19, SubBytesIns_Inst_Sbox_14_L18,
         SubBytesIns_Inst_Sbox_14_L17, SubBytesIns_Inst_Sbox_14_L16,
         SubBytesIns_Inst_Sbox_14_L15, SubBytesIns_Inst_Sbox_14_L14,
         SubBytesIns_Inst_Sbox_14_L13, SubBytesIns_Inst_Sbox_14_L12,
         SubBytesIns_Inst_Sbox_14_L11, SubBytesIns_Inst_Sbox_14_L10,
         SubBytesIns_Inst_Sbox_14_L9, SubBytesIns_Inst_Sbox_14_L8,
         SubBytesIns_Inst_Sbox_14_L7, SubBytesIns_Inst_Sbox_14_L6,
         SubBytesIns_Inst_Sbox_14_L5, SubBytesIns_Inst_Sbox_14_L4,
         SubBytesIns_Inst_Sbox_14_L3, SubBytesIns_Inst_Sbox_14_L2,
         SubBytesIns_Inst_Sbox_14_L1, SubBytesIns_Inst_Sbox_14_L0,
         SubBytesIns_Inst_Sbox_14_M63, SubBytesIns_Inst_Sbox_14_M62,
         SubBytesIns_Inst_Sbox_14_M61, SubBytesIns_Inst_Sbox_14_M60,
         SubBytesIns_Inst_Sbox_14_M59, SubBytesIns_Inst_Sbox_14_M58,
         SubBytesIns_Inst_Sbox_14_M57, SubBytesIns_Inst_Sbox_14_M56,
         SubBytesIns_Inst_Sbox_14_M55, SubBytesIns_Inst_Sbox_14_M54,
         SubBytesIns_Inst_Sbox_14_M53, SubBytesIns_Inst_Sbox_14_M52,
         SubBytesIns_Inst_Sbox_14_M51, SubBytesIns_Inst_Sbox_14_M50,
         SubBytesIns_Inst_Sbox_14_M49, SubBytesIns_Inst_Sbox_14_M48,
         SubBytesIns_Inst_Sbox_14_M47, SubBytesIns_Inst_Sbox_14_M46,
         SubBytesIns_Inst_Sbox_14_M45, SubBytesIns_Inst_Sbox_14_M44,
         SubBytesIns_Inst_Sbox_14_M43, SubBytesIns_Inst_Sbox_14_M42,
         SubBytesIns_Inst_Sbox_14_M41, SubBytesIns_Inst_Sbox_14_M40,
         SubBytesIns_Inst_Sbox_14_M39, SubBytesIns_Inst_Sbox_14_M38,
         SubBytesIns_Inst_Sbox_14_M37, SubBytesIns_Inst_Sbox_14_M36,
         SubBytesIns_Inst_Sbox_14_M35, SubBytesIns_Inst_Sbox_14_M34,
         SubBytesIns_Inst_Sbox_14_M33, SubBytesIns_Inst_Sbox_14_M32,
         SubBytesIns_Inst_Sbox_14_M31, SubBytesIns_Inst_Sbox_14_M30,
         SubBytesIns_Inst_Sbox_14_M29, SubBytesIns_Inst_Sbox_14_M28,
         SubBytesIns_Inst_Sbox_14_M27, SubBytesIns_Inst_Sbox_14_M26,
         SubBytesIns_Inst_Sbox_14_M25, SubBytesIns_Inst_Sbox_14_M24,
         SubBytesIns_Inst_Sbox_14_M23, SubBytesIns_Inst_Sbox_14_M22,
         SubBytesIns_Inst_Sbox_14_M21, SubBytesIns_Inst_Sbox_14_M20,
         SubBytesIns_Inst_Sbox_14_M19, SubBytesIns_Inst_Sbox_14_M18,
         SubBytesIns_Inst_Sbox_14_M17, SubBytesIns_Inst_Sbox_14_M16,
         SubBytesIns_Inst_Sbox_14_M15, SubBytesIns_Inst_Sbox_14_M14,
         SubBytesIns_Inst_Sbox_14_M13, SubBytesIns_Inst_Sbox_14_M12,
         SubBytesIns_Inst_Sbox_14_M11, SubBytesIns_Inst_Sbox_14_M10,
         SubBytesIns_Inst_Sbox_14_M9, SubBytesIns_Inst_Sbox_14_M8,
         SubBytesIns_Inst_Sbox_14_M7, SubBytesIns_Inst_Sbox_14_M6,
         SubBytesIns_Inst_Sbox_14_M5, SubBytesIns_Inst_Sbox_14_M4,
         SubBytesIns_Inst_Sbox_14_M3, SubBytesIns_Inst_Sbox_14_M2,
         SubBytesIns_Inst_Sbox_14_M1, SubBytesIns_Inst_Sbox_14_T27,
         SubBytesIns_Inst_Sbox_14_T26, SubBytesIns_Inst_Sbox_14_T25,
         SubBytesIns_Inst_Sbox_14_T24, SubBytesIns_Inst_Sbox_14_T23,
         SubBytesIns_Inst_Sbox_14_T22, SubBytesIns_Inst_Sbox_14_T21,
         SubBytesIns_Inst_Sbox_14_T20, SubBytesIns_Inst_Sbox_14_T19,
         SubBytesIns_Inst_Sbox_14_T18, SubBytesIns_Inst_Sbox_14_T17,
         SubBytesIns_Inst_Sbox_14_T16, SubBytesIns_Inst_Sbox_14_T15,
         SubBytesIns_Inst_Sbox_14_T14, SubBytesIns_Inst_Sbox_14_T13,
         SubBytesIns_Inst_Sbox_14_T12, SubBytesIns_Inst_Sbox_14_T11,
         SubBytesIns_Inst_Sbox_14_T10, SubBytesIns_Inst_Sbox_14_T9,
         SubBytesIns_Inst_Sbox_14_T8, SubBytesIns_Inst_Sbox_14_T7,
         SubBytesIns_Inst_Sbox_14_T6, SubBytesIns_Inst_Sbox_14_T5,
         SubBytesIns_Inst_Sbox_14_T4, SubBytesIns_Inst_Sbox_14_T3,
         SubBytesIns_Inst_Sbox_14_T2, SubBytesIns_Inst_Sbox_14_T1,
         SubBytesIns_Inst_Sbox_15_L29, SubBytesIns_Inst_Sbox_15_L28,
         SubBytesIns_Inst_Sbox_15_L27, SubBytesIns_Inst_Sbox_15_L26,
         SubBytesIns_Inst_Sbox_15_L25, SubBytesIns_Inst_Sbox_15_L24,
         SubBytesIns_Inst_Sbox_15_L23, SubBytesIns_Inst_Sbox_15_L22,
         SubBytesIns_Inst_Sbox_15_L21, SubBytesIns_Inst_Sbox_15_L20,
         SubBytesIns_Inst_Sbox_15_L19, SubBytesIns_Inst_Sbox_15_L18,
         SubBytesIns_Inst_Sbox_15_L17, SubBytesIns_Inst_Sbox_15_L16,
         SubBytesIns_Inst_Sbox_15_L15, SubBytesIns_Inst_Sbox_15_L14,
         SubBytesIns_Inst_Sbox_15_L13, SubBytesIns_Inst_Sbox_15_L12,
         SubBytesIns_Inst_Sbox_15_L11, SubBytesIns_Inst_Sbox_15_L10,
         SubBytesIns_Inst_Sbox_15_L9, SubBytesIns_Inst_Sbox_15_L8,
         SubBytesIns_Inst_Sbox_15_L7, SubBytesIns_Inst_Sbox_15_L6,
         SubBytesIns_Inst_Sbox_15_L5, SubBytesIns_Inst_Sbox_15_L4,
         SubBytesIns_Inst_Sbox_15_L3, SubBytesIns_Inst_Sbox_15_L2,
         SubBytesIns_Inst_Sbox_15_L1, SubBytesIns_Inst_Sbox_15_L0,
         SubBytesIns_Inst_Sbox_15_M63, SubBytesIns_Inst_Sbox_15_M62,
         SubBytesIns_Inst_Sbox_15_M61, SubBytesIns_Inst_Sbox_15_M60,
         SubBytesIns_Inst_Sbox_15_M59, SubBytesIns_Inst_Sbox_15_M58,
         SubBytesIns_Inst_Sbox_15_M57, SubBytesIns_Inst_Sbox_15_M56,
         SubBytesIns_Inst_Sbox_15_M55, SubBytesIns_Inst_Sbox_15_M54,
         SubBytesIns_Inst_Sbox_15_M53, SubBytesIns_Inst_Sbox_15_M52,
         SubBytesIns_Inst_Sbox_15_M51, SubBytesIns_Inst_Sbox_15_M50,
         SubBytesIns_Inst_Sbox_15_M49, SubBytesIns_Inst_Sbox_15_M48,
         SubBytesIns_Inst_Sbox_15_M47, SubBytesIns_Inst_Sbox_15_M46,
         SubBytesIns_Inst_Sbox_15_M45, SubBytesIns_Inst_Sbox_15_M44,
         SubBytesIns_Inst_Sbox_15_M43, SubBytesIns_Inst_Sbox_15_M42,
         SubBytesIns_Inst_Sbox_15_M41, SubBytesIns_Inst_Sbox_15_M40,
         SubBytesIns_Inst_Sbox_15_M39, SubBytesIns_Inst_Sbox_15_M38,
         SubBytesIns_Inst_Sbox_15_M37, SubBytesIns_Inst_Sbox_15_M36,
         SubBytesIns_Inst_Sbox_15_M35, SubBytesIns_Inst_Sbox_15_M34,
         SubBytesIns_Inst_Sbox_15_M33, SubBytesIns_Inst_Sbox_15_M32,
         SubBytesIns_Inst_Sbox_15_M31, SubBytesIns_Inst_Sbox_15_M30,
         SubBytesIns_Inst_Sbox_15_M29, SubBytesIns_Inst_Sbox_15_M28,
         SubBytesIns_Inst_Sbox_15_M27, SubBytesIns_Inst_Sbox_15_M26,
         SubBytesIns_Inst_Sbox_15_M25, SubBytesIns_Inst_Sbox_15_M24,
         SubBytesIns_Inst_Sbox_15_M23, SubBytesIns_Inst_Sbox_15_M22,
         SubBytesIns_Inst_Sbox_15_M21, SubBytesIns_Inst_Sbox_15_M20,
         SubBytesIns_Inst_Sbox_15_M19, SubBytesIns_Inst_Sbox_15_M18,
         SubBytesIns_Inst_Sbox_15_M17, SubBytesIns_Inst_Sbox_15_M16,
         SubBytesIns_Inst_Sbox_15_M15, SubBytesIns_Inst_Sbox_15_M14,
         SubBytesIns_Inst_Sbox_15_M13, SubBytesIns_Inst_Sbox_15_M12,
         SubBytesIns_Inst_Sbox_15_M11, SubBytesIns_Inst_Sbox_15_M10,
         SubBytesIns_Inst_Sbox_15_M9, SubBytesIns_Inst_Sbox_15_M8,
         SubBytesIns_Inst_Sbox_15_M7, SubBytesIns_Inst_Sbox_15_M6,
         SubBytesIns_Inst_Sbox_15_M5, SubBytesIns_Inst_Sbox_15_M4,
         SubBytesIns_Inst_Sbox_15_M3, SubBytesIns_Inst_Sbox_15_M2,
         SubBytesIns_Inst_Sbox_15_M1, SubBytesIns_Inst_Sbox_15_T27,
         SubBytesIns_Inst_Sbox_15_T26, SubBytesIns_Inst_Sbox_15_T25,
         SubBytesIns_Inst_Sbox_15_T24, SubBytesIns_Inst_Sbox_15_T23,
         SubBytesIns_Inst_Sbox_15_T22, SubBytesIns_Inst_Sbox_15_T21,
         SubBytesIns_Inst_Sbox_15_T20, SubBytesIns_Inst_Sbox_15_T19,
         SubBytesIns_Inst_Sbox_15_T18, SubBytesIns_Inst_Sbox_15_T17,
         SubBytesIns_Inst_Sbox_15_T16, SubBytesIns_Inst_Sbox_15_T15,
         SubBytesIns_Inst_Sbox_15_T14, SubBytesIns_Inst_Sbox_15_T13,
         SubBytesIns_Inst_Sbox_15_T12, SubBytesIns_Inst_Sbox_15_T11,
         SubBytesIns_Inst_Sbox_15_T10, SubBytesIns_Inst_Sbox_15_T9,
         SubBytesIns_Inst_Sbox_15_T8, SubBytesIns_Inst_Sbox_15_T7,
         SubBytesIns_Inst_Sbox_15_T6, SubBytesIns_Inst_Sbox_15_T5,
         SubBytesIns_Inst_Sbox_15_T4, SubBytesIns_Inst_Sbox_15_T3,
         SubBytesIns_Inst_Sbox_15_T2, SubBytesIns_Inst_Sbox_15_T1,
         MixColumnsIns_MixOneColumnInst_0_n64,
         MixColumnsIns_MixOneColumnInst_0_n63,
         MixColumnsIns_MixOneColumnInst_0_n62,
         MixColumnsIns_MixOneColumnInst_0_n61,
         MixColumnsIns_MixOneColumnInst_0_n60,
         MixColumnsIns_MixOneColumnInst_0_n59,
         MixColumnsIns_MixOneColumnInst_0_n58,
         MixColumnsIns_MixOneColumnInst_0_n57,
         MixColumnsIns_MixOneColumnInst_0_n56,
         MixColumnsIns_MixOneColumnInst_0_n55,
         MixColumnsIns_MixOneColumnInst_0_n54,
         MixColumnsIns_MixOneColumnInst_0_n53,
         MixColumnsIns_MixOneColumnInst_0_n52,
         MixColumnsIns_MixOneColumnInst_0_n51,
         MixColumnsIns_MixOneColumnInst_0_n50,
         MixColumnsIns_MixOneColumnInst_0_n49,
         MixColumnsIns_MixOneColumnInst_0_n48,
         MixColumnsIns_MixOneColumnInst_0_n47,
         MixColumnsIns_MixOneColumnInst_0_n46,
         MixColumnsIns_MixOneColumnInst_0_n45,
         MixColumnsIns_MixOneColumnInst_0_n44,
         MixColumnsIns_MixOneColumnInst_0_n43,
         MixColumnsIns_MixOneColumnInst_0_n42,
         MixColumnsIns_MixOneColumnInst_0_n41,
         MixColumnsIns_MixOneColumnInst_0_n40,
         MixColumnsIns_MixOneColumnInst_0_n39,
         MixColumnsIns_MixOneColumnInst_0_n38,
         MixColumnsIns_MixOneColumnInst_0_n37,
         MixColumnsIns_MixOneColumnInst_0_n36,
         MixColumnsIns_MixOneColumnInst_0_n35,
         MixColumnsIns_MixOneColumnInst_0_n34,
         MixColumnsIns_MixOneColumnInst_0_n33,
         MixColumnsIns_MixOneColumnInst_0_n32,
         MixColumnsIns_MixOneColumnInst_0_n31,
         MixColumnsIns_MixOneColumnInst_0_n30,
         MixColumnsIns_MixOneColumnInst_0_n29,
         MixColumnsIns_MixOneColumnInst_0_n28,
         MixColumnsIns_MixOneColumnInst_0_n27,
         MixColumnsIns_MixOneColumnInst_0_n26,
         MixColumnsIns_MixOneColumnInst_0_n25,
         MixColumnsIns_MixOneColumnInst_0_n24,
         MixColumnsIns_MixOneColumnInst_0_n23,
         MixColumnsIns_MixOneColumnInst_0_n22,
         MixColumnsIns_MixOneColumnInst_0_n21,
         MixColumnsIns_MixOneColumnInst_0_n20,
         MixColumnsIns_MixOneColumnInst_0_n19,
         MixColumnsIns_MixOneColumnInst_0_n18,
         MixColumnsIns_MixOneColumnInst_0_n17,
         MixColumnsIns_MixOneColumnInst_0_n16,
         MixColumnsIns_MixOneColumnInst_0_n15,
         MixColumnsIns_MixOneColumnInst_0_n14,
         MixColumnsIns_MixOneColumnInst_0_n13,
         MixColumnsIns_MixOneColumnInst_0_n12,
         MixColumnsIns_MixOneColumnInst_0_n11,
         MixColumnsIns_MixOneColumnInst_0_n10,
         MixColumnsIns_MixOneColumnInst_0_n9,
         MixColumnsIns_MixOneColumnInst_0_n8,
         MixColumnsIns_MixOneColumnInst_0_n7,
         MixColumnsIns_MixOneColumnInst_0_n6,
         MixColumnsIns_MixOneColumnInst_0_n5,
         MixColumnsIns_MixOneColumnInst_0_n4,
         MixColumnsIns_MixOneColumnInst_0_n3,
         MixColumnsIns_MixOneColumnInst_0_n2,
         MixColumnsIns_MixOneColumnInst_0_n1,
         MixColumnsIns_MixOneColumnInst_1_n64,
         MixColumnsIns_MixOneColumnInst_1_n63,
         MixColumnsIns_MixOneColumnInst_1_n62,
         MixColumnsIns_MixOneColumnInst_1_n61,
         MixColumnsIns_MixOneColumnInst_1_n60,
         MixColumnsIns_MixOneColumnInst_1_n59,
         MixColumnsIns_MixOneColumnInst_1_n58,
         MixColumnsIns_MixOneColumnInst_1_n57,
         MixColumnsIns_MixOneColumnInst_1_n56,
         MixColumnsIns_MixOneColumnInst_1_n55,
         MixColumnsIns_MixOneColumnInst_1_n54,
         MixColumnsIns_MixOneColumnInst_1_n53,
         MixColumnsIns_MixOneColumnInst_1_n52,
         MixColumnsIns_MixOneColumnInst_1_n51,
         MixColumnsIns_MixOneColumnInst_1_n50,
         MixColumnsIns_MixOneColumnInst_1_n49,
         MixColumnsIns_MixOneColumnInst_1_n48,
         MixColumnsIns_MixOneColumnInst_1_n47,
         MixColumnsIns_MixOneColumnInst_1_n46,
         MixColumnsIns_MixOneColumnInst_1_n45,
         MixColumnsIns_MixOneColumnInst_1_n44,
         MixColumnsIns_MixOneColumnInst_1_n43,
         MixColumnsIns_MixOneColumnInst_1_n42,
         MixColumnsIns_MixOneColumnInst_1_n41,
         MixColumnsIns_MixOneColumnInst_1_n40,
         MixColumnsIns_MixOneColumnInst_1_n39,
         MixColumnsIns_MixOneColumnInst_1_n38,
         MixColumnsIns_MixOneColumnInst_1_n37,
         MixColumnsIns_MixOneColumnInst_1_n36,
         MixColumnsIns_MixOneColumnInst_1_n35,
         MixColumnsIns_MixOneColumnInst_1_n34,
         MixColumnsIns_MixOneColumnInst_1_n33,
         MixColumnsIns_MixOneColumnInst_1_n32,
         MixColumnsIns_MixOneColumnInst_1_n31,
         MixColumnsIns_MixOneColumnInst_1_n30,
         MixColumnsIns_MixOneColumnInst_1_n29,
         MixColumnsIns_MixOneColumnInst_1_n28,
         MixColumnsIns_MixOneColumnInst_1_n27,
         MixColumnsIns_MixOneColumnInst_1_n26,
         MixColumnsIns_MixOneColumnInst_1_n25,
         MixColumnsIns_MixOneColumnInst_1_n24,
         MixColumnsIns_MixOneColumnInst_1_n23,
         MixColumnsIns_MixOneColumnInst_1_n22,
         MixColumnsIns_MixOneColumnInst_1_n21,
         MixColumnsIns_MixOneColumnInst_1_n20,
         MixColumnsIns_MixOneColumnInst_1_n19,
         MixColumnsIns_MixOneColumnInst_1_n18,
         MixColumnsIns_MixOneColumnInst_1_n17,
         MixColumnsIns_MixOneColumnInst_1_n16,
         MixColumnsIns_MixOneColumnInst_1_n15,
         MixColumnsIns_MixOneColumnInst_1_n14,
         MixColumnsIns_MixOneColumnInst_1_n13,
         MixColumnsIns_MixOneColumnInst_1_n12,
         MixColumnsIns_MixOneColumnInst_1_n11,
         MixColumnsIns_MixOneColumnInst_1_n10,
         MixColumnsIns_MixOneColumnInst_1_n9,
         MixColumnsIns_MixOneColumnInst_1_n8,
         MixColumnsIns_MixOneColumnInst_1_n7,
         MixColumnsIns_MixOneColumnInst_1_n6,
         MixColumnsIns_MixOneColumnInst_1_n5,
         MixColumnsIns_MixOneColumnInst_1_n4,
         MixColumnsIns_MixOneColumnInst_1_n3,
         MixColumnsIns_MixOneColumnInst_1_n2,
         MixColumnsIns_MixOneColumnInst_1_n1,
         MixColumnsIns_MixOneColumnInst_2_n64,
         MixColumnsIns_MixOneColumnInst_2_n63,
         MixColumnsIns_MixOneColumnInst_2_n62,
         MixColumnsIns_MixOneColumnInst_2_n61,
         MixColumnsIns_MixOneColumnInst_2_n60,
         MixColumnsIns_MixOneColumnInst_2_n59,
         MixColumnsIns_MixOneColumnInst_2_n58,
         MixColumnsIns_MixOneColumnInst_2_n57,
         MixColumnsIns_MixOneColumnInst_2_n56,
         MixColumnsIns_MixOneColumnInst_2_n55,
         MixColumnsIns_MixOneColumnInst_2_n54,
         MixColumnsIns_MixOneColumnInst_2_n53,
         MixColumnsIns_MixOneColumnInst_2_n52,
         MixColumnsIns_MixOneColumnInst_2_n51,
         MixColumnsIns_MixOneColumnInst_2_n50,
         MixColumnsIns_MixOneColumnInst_2_n49,
         MixColumnsIns_MixOneColumnInst_2_n48,
         MixColumnsIns_MixOneColumnInst_2_n47,
         MixColumnsIns_MixOneColumnInst_2_n46,
         MixColumnsIns_MixOneColumnInst_2_n45,
         MixColumnsIns_MixOneColumnInst_2_n44,
         MixColumnsIns_MixOneColumnInst_2_n43,
         MixColumnsIns_MixOneColumnInst_2_n42,
         MixColumnsIns_MixOneColumnInst_2_n41,
         MixColumnsIns_MixOneColumnInst_2_n40,
         MixColumnsIns_MixOneColumnInst_2_n39,
         MixColumnsIns_MixOneColumnInst_2_n38,
         MixColumnsIns_MixOneColumnInst_2_n37,
         MixColumnsIns_MixOneColumnInst_2_n36,
         MixColumnsIns_MixOneColumnInst_2_n35,
         MixColumnsIns_MixOneColumnInst_2_n34,
         MixColumnsIns_MixOneColumnInst_2_n33,
         MixColumnsIns_MixOneColumnInst_2_n32,
         MixColumnsIns_MixOneColumnInst_2_n31,
         MixColumnsIns_MixOneColumnInst_2_n30,
         MixColumnsIns_MixOneColumnInst_2_n29,
         MixColumnsIns_MixOneColumnInst_2_n28,
         MixColumnsIns_MixOneColumnInst_2_n27,
         MixColumnsIns_MixOneColumnInst_2_n26,
         MixColumnsIns_MixOneColumnInst_2_n25,
         MixColumnsIns_MixOneColumnInst_2_n24,
         MixColumnsIns_MixOneColumnInst_2_n23,
         MixColumnsIns_MixOneColumnInst_2_n22,
         MixColumnsIns_MixOneColumnInst_2_n21,
         MixColumnsIns_MixOneColumnInst_2_n20,
         MixColumnsIns_MixOneColumnInst_2_n19,
         MixColumnsIns_MixOneColumnInst_2_n18,
         MixColumnsIns_MixOneColumnInst_2_n17,
         MixColumnsIns_MixOneColumnInst_2_n16,
         MixColumnsIns_MixOneColumnInst_2_n15,
         MixColumnsIns_MixOneColumnInst_2_n14,
         MixColumnsIns_MixOneColumnInst_2_n13,
         MixColumnsIns_MixOneColumnInst_2_n12,
         MixColumnsIns_MixOneColumnInst_2_n11,
         MixColumnsIns_MixOneColumnInst_2_n10,
         MixColumnsIns_MixOneColumnInst_2_n9,
         MixColumnsIns_MixOneColumnInst_2_n8,
         MixColumnsIns_MixOneColumnInst_2_n7,
         MixColumnsIns_MixOneColumnInst_2_n6,
         MixColumnsIns_MixOneColumnInst_2_n5,
         MixColumnsIns_MixOneColumnInst_2_n4,
         MixColumnsIns_MixOneColumnInst_2_n3,
         MixColumnsIns_MixOneColumnInst_2_n2,
         MixColumnsIns_MixOneColumnInst_2_n1,
         MixColumnsIns_MixOneColumnInst_3_n64,
         MixColumnsIns_MixOneColumnInst_3_n63,
         MixColumnsIns_MixOneColumnInst_3_n62,
         MixColumnsIns_MixOneColumnInst_3_n61,
         MixColumnsIns_MixOneColumnInst_3_n60,
         MixColumnsIns_MixOneColumnInst_3_n59,
         MixColumnsIns_MixOneColumnInst_3_n58,
         MixColumnsIns_MixOneColumnInst_3_n57,
         MixColumnsIns_MixOneColumnInst_3_n56,
         MixColumnsIns_MixOneColumnInst_3_n55,
         MixColumnsIns_MixOneColumnInst_3_n54,
         MixColumnsIns_MixOneColumnInst_3_n53,
         MixColumnsIns_MixOneColumnInst_3_n52,
         MixColumnsIns_MixOneColumnInst_3_n51,
         MixColumnsIns_MixOneColumnInst_3_n50,
         MixColumnsIns_MixOneColumnInst_3_n49,
         MixColumnsIns_MixOneColumnInst_3_n48,
         MixColumnsIns_MixOneColumnInst_3_n47,
         MixColumnsIns_MixOneColumnInst_3_n46,
         MixColumnsIns_MixOneColumnInst_3_n45,
         MixColumnsIns_MixOneColumnInst_3_n44,
         MixColumnsIns_MixOneColumnInst_3_n43,
         MixColumnsIns_MixOneColumnInst_3_n42,
         MixColumnsIns_MixOneColumnInst_3_n41,
         MixColumnsIns_MixOneColumnInst_3_n40,
         MixColumnsIns_MixOneColumnInst_3_n39,
         MixColumnsIns_MixOneColumnInst_3_n38,
         MixColumnsIns_MixOneColumnInst_3_n37,
         MixColumnsIns_MixOneColumnInst_3_n36,
         MixColumnsIns_MixOneColumnInst_3_n35,
         MixColumnsIns_MixOneColumnInst_3_n34,
         MixColumnsIns_MixOneColumnInst_3_n33,
         MixColumnsIns_MixOneColumnInst_3_n32,
         MixColumnsIns_MixOneColumnInst_3_n31,
         MixColumnsIns_MixOneColumnInst_3_n30,
         MixColumnsIns_MixOneColumnInst_3_n29,
         MixColumnsIns_MixOneColumnInst_3_n28,
         MixColumnsIns_MixOneColumnInst_3_n27,
         MixColumnsIns_MixOneColumnInst_3_n26,
         MixColumnsIns_MixOneColumnInst_3_n25,
         MixColumnsIns_MixOneColumnInst_3_n24,
         MixColumnsIns_MixOneColumnInst_3_n23,
         MixColumnsIns_MixOneColumnInst_3_n22,
         MixColumnsIns_MixOneColumnInst_3_n21,
         MixColumnsIns_MixOneColumnInst_3_n20,
         MixColumnsIns_MixOneColumnInst_3_n19,
         MixColumnsIns_MixOneColumnInst_3_n18,
         MixColumnsIns_MixOneColumnInst_3_n17,
         MixColumnsIns_MixOneColumnInst_3_n16,
         MixColumnsIns_MixOneColumnInst_3_n15,
         MixColumnsIns_MixOneColumnInst_3_n14,
         MixColumnsIns_MixOneColumnInst_3_n13,
         MixColumnsIns_MixOneColumnInst_3_n12,
         MixColumnsIns_MixOneColumnInst_3_n11,
         MixColumnsIns_MixOneColumnInst_3_n10,
         MixColumnsIns_MixOneColumnInst_3_n9,
         MixColumnsIns_MixOneColumnInst_3_n8,
         MixColumnsIns_MixOneColumnInst_3_n7,
         MixColumnsIns_MixOneColumnInst_3_n6,
         MixColumnsIns_MixOneColumnInst_3_n5,
         MixColumnsIns_MixOneColumnInst_3_n4,
         MixColumnsIns_MixOneColumnInst_3_n3,
         MixColumnsIns_MixOneColumnInst_3_n2,
         MixColumnsIns_MixOneColumnInst_3_n1, KeyReg_Inst_ff_SDE_0_next_state,
         KeyReg_Inst_ff_SDE_0_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_1_next_state,
         KeyReg_Inst_ff_SDE_1_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_2_next_state,
         KeyReg_Inst_ff_SDE_2_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_3_next_state,
         KeyReg_Inst_ff_SDE_3_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_4_next_state,
         KeyReg_Inst_ff_SDE_4_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_5_next_state,
         KeyReg_Inst_ff_SDE_5_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_6_next_state,
         KeyReg_Inst_ff_SDE_6_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_7_next_state,
         KeyReg_Inst_ff_SDE_7_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_8_next_state,
         KeyReg_Inst_ff_SDE_8_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_9_next_state,
         KeyReg_Inst_ff_SDE_9_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_10_next_state,
         KeyReg_Inst_ff_SDE_10_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_11_next_state,
         KeyReg_Inst_ff_SDE_11_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_12_next_state,
         KeyReg_Inst_ff_SDE_12_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_13_next_state,
         KeyReg_Inst_ff_SDE_13_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_14_next_state,
         KeyReg_Inst_ff_SDE_14_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_15_next_state,
         KeyReg_Inst_ff_SDE_15_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_16_next_state,
         KeyReg_Inst_ff_SDE_16_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_17_next_state,
         KeyReg_Inst_ff_SDE_17_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_18_next_state,
         KeyReg_Inst_ff_SDE_18_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_19_next_state,
         KeyReg_Inst_ff_SDE_19_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_20_next_state,
         KeyReg_Inst_ff_SDE_20_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_21_next_state,
         KeyReg_Inst_ff_SDE_21_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_22_next_state,
         KeyReg_Inst_ff_SDE_22_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_23_next_state,
         KeyReg_Inst_ff_SDE_23_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_24_next_state,
         KeyReg_Inst_ff_SDE_24_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_25_next_state,
         KeyReg_Inst_ff_SDE_25_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_26_next_state,
         KeyReg_Inst_ff_SDE_26_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_27_next_state,
         KeyReg_Inst_ff_SDE_27_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_28_next_state,
         KeyReg_Inst_ff_SDE_28_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_29_next_state,
         KeyReg_Inst_ff_SDE_29_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_30_next_state,
         KeyReg_Inst_ff_SDE_30_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_31_next_state,
         KeyReg_Inst_ff_SDE_31_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_32_next_state,
         KeyReg_Inst_ff_SDE_32_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_33_next_state,
         KeyReg_Inst_ff_SDE_33_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_34_next_state,
         KeyReg_Inst_ff_SDE_34_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_35_next_state,
         KeyReg_Inst_ff_SDE_35_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_36_next_state,
         KeyReg_Inst_ff_SDE_36_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_37_next_state,
         KeyReg_Inst_ff_SDE_37_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_38_next_state,
         KeyReg_Inst_ff_SDE_38_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_39_next_state,
         KeyReg_Inst_ff_SDE_39_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_40_next_state,
         KeyReg_Inst_ff_SDE_40_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_41_next_state,
         KeyReg_Inst_ff_SDE_41_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_42_next_state,
         KeyReg_Inst_ff_SDE_42_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_43_next_state,
         KeyReg_Inst_ff_SDE_43_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_44_next_state,
         KeyReg_Inst_ff_SDE_44_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_45_next_state,
         KeyReg_Inst_ff_SDE_45_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_46_next_state,
         KeyReg_Inst_ff_SDE_46_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_47_next_state,
         KeyReg_Inst_ff_SDE_47_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_48_next_state,
         KeyReg_Inst_ff_SDE_48_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_49_next_state,
         KeyReg_Inst_ff_SDE_49_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_50_next_state,
         KeyReg_Inst_ff_SDE_50_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_51_next_state,
         KeyReg_Inst_ff_SDE_51_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_52_next_state,
         KeyReg_Inst_ff_SDE_52_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_53_next_state,
         KeyReg_Inst_ff_SDE_53_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_54_next_state,
         KeyReg_Inst_ff_SDE_54_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_55_next_state,
         KeyReg_Inst_ff_SDE_55_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_56_next_state,
         KeyReg_Inst_ff_SDE_56_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_57_next_state,
         KeyReg_Inst_ff_SDE_57_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_58_next_state,
         KeyReg_Inst_ff_SDE_58_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_59_next_state,
         KeyReg_Inst_ff_SDE_59_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_60_next_state,
         KeyReg_Inst_ff_SDE_60_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_61_next_state,
         KeyReg_Inst_ff_SDE_61_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_62_next_state,
         KeyReg_Inst_ff_SDE_62_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_63_next_state,
         KeyReg_Inst_ff_SDE_63_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_64_next_state,
         KeyReg_Inst_ff_SDE_64_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_65_next_state,
         KeyReg_Inst_ff_SDE_65_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_66_next_state,
         KeyReg_Inst_ff_SDE_66_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_67_next_state,
         KeyReg_Inst_ff_SDE_67_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_68_next_state,
         KeyReg_Inst_ff_SDE_68_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_69_next_state,
         KeyReg_Inst_ff_SDE_69_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_70_next_state,
         KeyReg_Inst_ff_SDE_70_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_71_next_state,
         KeyReg_Inst_ff_SDE_71_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_72_next_state,
         KeyReg_Inst_ff_SDE_72_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_73_next_state,
         KeyReg_Inst_ff_SDE_73_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_74_next_state,
         KeyReg_Inst_ff_SDE_74_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_75_next_state,
         KeyReg_Inst_ff_SDE_75_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_76_next_state,
         KeyReg_Inst_ff_SDE_76_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_77_next_state,
         KeyReg_Inst_ff_SDE_77_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_78_next_state,
         KeyReg_Inst_ff_SDE_78_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_79_next_state,
         KeyReg_Inst_ff_SDE_79_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_80_next_state,
         KeyReg_Inst_ff_SDE_80_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_81_next_state,
         KeyReg_Inst_ff_SDE_81_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_82_next_state,
         KeyReg_Inst_ff_SDE_82_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_83_next_state,
         KeyReg_Inst_ff_SDE_83_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_84_next_state,
         KeyReg_Inst_ff_SDE_84_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_85_next_state,
         KeyReg_Inst_ff_SDE_85_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_86_next_state,
         KeyReg_Inst_ff_SDE_86_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_87_next_state,
         KeyReg_Inst_ff_SDE_87_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_88_next_state,
         KeyReg_Inst_ff_SDE_88_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_89_next_state,
         KeyReg_Inst_ff_SDE_89_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_90_next_state,
         KeyReg_Inst_ff_SDE_90_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_91_next_state,
         KeyReg_Inst_ff_SDE_91_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_92_next_state,
         KeyReg_Inst_ff_SDE_92_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_93_next_state,
         KeyReg_Inst_ff_SDE_93_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_94_next_state,
         KeyReg_Inst_ff_SDE_94_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_95_next_state,
         KeyReg_Inst_ff_SDE_95_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_96_next_state,
         KeyReg_Inst_ff_SDE_96_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_97_next_state,
         KeyReg_Inst_ff_SDE_97_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_98_next_state,
         KeyReg_Inst_ff_SDE_98_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_99_next_state,
         KeyReg_Inst_ff_SDE_99_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_100_next_state,
         KeyReg_Inst_ff_SDE_100_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_101_next_state,
         KeyReg_Inst_ff_SDE_101_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_102_next_state,
         KeyReg_Inst_ff_SDE_102_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_103_next_state,
         KeyReg_Inst_ff_SDE_103_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_104_next_state,
         KeyReg_Inst_ff_SDE_104_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_105_next_state,
         KeyReg_Inst_ff_SDE_105_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_106_next_state,
         KeyReg_Inst_ff_SDE_106_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_107_next_state,
         KeyReg_Inst_ff_SDE_107_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_108_next_state,
         KeyReg_Inst_ff_SDE_108_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_109_next_state,
         KeyReg_Inst_ff_SDE_109_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_110_next_state,
         KeyReg_Inst_ff_SDE_110_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_111_next_state,
         KeyReg_Inst_ff_SDE_111_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_112_next_state,
         KeyReg_Inst_ff_SDE_112_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_113_next_state,
         KeyReg_Inst_ff_SDE_113_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_114_next_state,
         KeyReg_Inst_ff_SDE_114_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_115_next_state,
         KeyReg_Inst_ff_SDE_115_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_116_next_state,
         KeyReg_Inst_ff_SDE_116_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_117_next_state,
         KeyReg_Inst_ff_SDE_117_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_118_next_state,
         KeyReg_Inst_ff_SDE_118_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_119_next_state,
         KeyReg_Inst_ff_SDE_119_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_120_next_state,
         KeyReg_Inst_ff_SDE_120_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_121_next_state,
         KeyReg_Inst_ff_SDE_121_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_122_next_state,
         KeyReg_Inst_ff_SDE_122_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_123_next_state,
         KeyReg_Inst_ff_SDE_123_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_124_next_state,
         KeyReg_Inst_ff_SDE_124_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_125_next_state,
         KeyReg_Inst_ff_SDE_125_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_126_next_state,
         KeyReg_Inst_ff_SDE_126_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_127_next_state,
         KeyReg_Inst_ff_SDE_127_current_state_reg_QN,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1, RoundCounterIns_n13,
         RoundCounterIns_n12, RoundCounterIns_n11, RoundCounterIns_n10,
         RoundCounterIns_n9, RoundCounterIns_n8, RoundCounterIns_n7,
         RoundCounterIns_n4, RoundCounterIns_n3, RoundCounterIns_n2,
         RoundCounterIns_n1, RoundCounterIns_N10, RoundCounterIns_n5,
         RoundCounterIns_N8, RoundCounterIns_n6, RoundCounterIns_N7,
         RoundCounterIns_count_reg_1__QN, RoundCounterIns_count_reg_3__QN;
  wire   [127:0] RoundOutput;
  wire   [127:0] RoundInput;
  wire   [123:0] MixColumnsInput;
  wire   [127:0] MixColumnsOutput;
  wire   [127:0] KeyExpansionOutput;
  wire   [127:0] RoundKey;
  wire   [5:0] Rcon;
  wire   [3:0] RoundCounter;
  wire   [31:0] MixColumnsIns_MixOneColumnInst_0_DoubleBytes;
  wire   [31:0] MixColumnsIns_MixOneColumnInst_1_DoubleBytes;
  wire   [31:0] MixColumnsIns_MixOneColumnInst_2_DoubleBytes;
  wire   [31:0] MixColumnsIns_MixOneColumnInst_3_DoubleBytes;
  wire   [31:0] KeyExpansionIns_tmp;

  INV_X1 U830 ( .A(n314), .ZN(n319) );
  INV_X1 U831 ( .A(n314), .ZN(n320) );
  INV_X1 U832 ( .A(n314), .ZN(n317) );
  INV_X1 U833 ( .A(n314), .ZN(n315) );
  INV_X1 U834 ( .A(n314), .ZN(n316) );
  INV_X1 U835 ( .A(n314), .ZN(n318) );
  NOR2_X1 U836 ( .A1(n325), .A2(n330), .ZN(n314) );
  INV_X1 U837 ( .A(RoundCounter[0]), .ZN(n325) );
  INV_X1 U838 ( .A(n314), .ZN(n321) );
  NOR2_X1 U839 ( .A1(RoundCounter[2]), .A2(RoundCounter[1]), .ZN(n323) );
  INV_X1 U840 ( .A(n323), .ZN(n322) );
  NOR2_X1 U841 ( .A1(RoundCounter[0]), .A2(n322), .ZN(Rcon[0]) );
  NOR2_X1 U842 ( .A1(RoundCounter[0]), .A2(RoundCounter[3]), .ZN(n337) );
  NOR2_X1 U843 ( .A1(n337), .A2(n322), .ZN(Rcon[1]) );
  NAND2_X1 U844 ( .A1(RoundCounter[3]), .A2(n323), .ZN(n330) );
  INV_X1 U845 ( .A(RoundCounter[2]), .ZN(n328) );
  AND2_X1 U846 ( .A1(n328), .A2(RoundCounter[1]), .ZN(n333) );
  NAND2_X1 U847 ( .A1(n337), .A2(n333), .ZN(n324) );
  NAND2_X1 U848 ( .A1(n321), .A2(n324), .ZN(Rcon[2]) );
  NOR2_X1 U849 ( .A1(RoundCounter[3]), .A2(n325), .ZN(n335) );
  NAND2_X1 U850 ( .A1(n333), .A2(n335), .ZN(n327) );
  NAND2_X1 U851 ( .A1(RoundCounter[3]), .A2(Rcon[0]), .ZN(n326) );
  NAND2_X1 U852 ( .A1(n327), .A2(n326), .ZN(Rcon[3]) );
  NOR2_X1 U853 ( .A1(RoundCounter[1]), .A2(n328), .ZN(n331) );
  NAND2_X1 U854 ( .A1(n337), .A2(n331), .ZN(n329) );
  NAND2_X1 U855 ( .A1(n330), .A2(n329), .ZN(Rcon[4]) );
  NAND2_X1 U856 ( .A1(n335), .A2(n331), .ZN(n332) );
  NAND2_X1 U857 ( .A1(n321), .A2(n332), .ZN(Rcon[5]) );
  MUX2_X1 U858 ( .A(MixColumnsInput[0]), .B(MixColumnsOutput[0]), .S(n321), 
        .Z(RoundOutput[0]) );
  MUX2_X1 U859 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B(
        MixColumnsOutput[100]), .S(n321), .Z(RoundOutput[100]) );
  MUX2_X1 U860 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B(
        MixColumnsOutput[101]), .S(n321), .Z(RoundOutput[101]) );
  MUX2_X1 U861 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B(
        MixColumnsOutput[102]), .S(n321), .Z(RoundOutput[102]) );
  MUX2_X1 U862 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsOutput[103]), .S(n321), .Z(RoundOutput[103]) );
  MUX2_X1 U863 ( .A(MixColumnsInput[104]), .B(MixColumnsOutput[104]), .S(n321), 
        .Z(RoundOutput[104]) );
  MUX2_X1 U864 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .B(
        MixColumnsOutput[105]), .S(n321), .Z(RoundOutput[105]) );
  MUX2_X1 U865 ( .A(MixColumnsInput[106]), .B(MixColumnsOutput[106]), .S(n321), 
        .Z(RoundOutput[106]) );
  MUX2_X1 U866 ( .A(MixColumnsInput[107]), .B(MixColumnsOutput[107]), .S(n315), 
        .Z(RoundOutput[107]) );
  MUX2_X1 U867 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .B(
        MixColumnsOutput[108]), .S(n316), .Z(RoundOutput[108]) );
  MUX2_X1 U868 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .B(
        MixColumnsOutput[109]), .S(n317), .Z(RoundOutput[109]) );
  MUX2_X1 U869 ( .A(MixColumnsInput[10]), .B(MixColumnsOutput[10]), .S(n318), 
        .Z(RoundOutput[10]) );
  MUX2_X1 U870 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .B(
        MixColumnsOutput[110]), .S(n319), .Z(RoundOutput[110]) );
  MUX2_X1 U871 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsOutput[111]), .S(n320), .Z(RoundOutput[111]) );
  MUX2_X1 U872 ( .A(MixColumnsInput[112]), .B(MixColumnsOutput[112]), .S(n319), 
        .Z(RoundOutput[112]) );
  MUX2_X1 U873 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .B(
        MixColumnsOutput[113]), .S(n318), .Z(RoundOutput[113]) );
  MUX2_X1 U874 ( .A(MixColumnsInput[114]), .B(MixColumnsOutput[114]), .S(n318), 
        .Z(RoundOutput[114]) );
  MUX2_X1 U875 ( .A(MixColumnsInput[115]), .B(MixColumnsOutput[115]), .S(n315), 
        .Z(RoundOutput[115]) );
  MUX2_X1 U876 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .B(
        MixColumnsOutput[116]), .S(n316), .Z(RoundOutput[116]) );
  MUX2_X1 U877 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .B(
        MixColumnsOutput[117]), .S(n317), .Z(RoundOutput[117]) );
  MUX2_X1 U878 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .B(
        MixColumnsOutput[118]), .S(n319), .Z(RoundOutput[118]) );
  MUX2_X1 U879 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B(
        MixColumnsOutput[119]), .S(n320), .Z(RoundOutput[119]) );
  MUX2_X1 U880 ( .A(MixColumnsInput[11]), .B(MixColumnsOutput[11]), .S(n320), 
        .Z(RoundOutput[11]) );
  MUX2_X1 U881 ( .A(MixColumnsInput[120]), .B(MixColumnsOutput[120]), .S(n319), 
        .Z(RoundOutput[120]) );
  MUX2_X1 U882 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .B(
        MixColumnsOutput[121]), .S(n318), .Z(RoundOutput[121]) );
  MUX2_X1 U883 ( .A(MixColumnsInput[122]), .B(MixColumnsOutput[122]), .S(n319), 
        .Z(RoundOutput[122]) );
  MUX2_X1 U884 ( .A(MixColumnsInput[123]), .B(MixColumnsOutput[123]), .S(n320), 
        .Z(RoundOutput[123]) );
  MUX2_X1 U885 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .B(
        MixColumnsOutput[124]), .S(n316), .Z(RoundOutput[124]) );
  MUX2_X1 U886 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .B(
        MixColumnsOutput[125]), .S(n320), .Z(RoundOutput[125]) );
  MUX2_X1 U887 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .B(
        MixColumnsOutput[126]), .S(n316), .Z(RoundOutput[126]) );
  MUX2_X1 U888 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B(
        MixColumnsOutput[127]), .S(n317), .Z(RoundOutput[127]) );
  MUX2_X1 U889 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .B(
        MixColumnsOutput[12]), .S(n315), .Z(RoundOutput[12]) );
  MUX2_X1 U890 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .B(
        MixColumnsOutput[13]), .S(n317), .Z(RoundOutput[13]) );
  MUX2_X1 U891 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .B(
        MixColumnsOutput[14]), .S(n316), .Z(RoundOutput[14]) );
  MUX2_X1 U892 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsOutput[15]), .S(n317), .Z(RoundOutput[15]) );
  MUX2_X1 U893 ( .A(MixColumnsInput[16]), .B(MixColumnsOutput[16]), .S(n315), 
        .Z(RoundOutput[16]) );
  MUX2_X1 U894 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .B(
        MixColumnsOutput[17]), .S(n318), .Z(RoundOutput[17]) );
  MUX2_X1 U895 ( .A(MixColumnsInput[18]), .B(MixColumnsOutput[18]), .S(n319), 
        .Z(RoundOutput[18]) );
  MUX2_X1 U896 ( .A(MixColumnsInput[19]), .B(MixColumnsOutput[19]), .S(n320), 
        .Z(RoundOutput[19]) );
  MUX2_X1 U897 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .B(
        MixColumnsOutput[1]), .S(n318), .Z(RoundOutput[1]) );
  MUX2_X1 U898 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .B(
        MixColumnsOutput[20]), .S(n319), .Z(RoundOutput[20]) );
  MUX2_X1 U899 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .B(
        MixColumnsOutput[21]), .S(n316), .Z(RoundOutput[21]) );
  MUX2_X1 U900 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .B(
        MixColumnsOutput[22]), .S(n317), .Z(RoundOutput[22]) );
  MUX2_X1 U901 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B(
        MixColumnsOutput[23]), .S(n315), .Z(RoundOutput[23]) );
  MUX2_X1 U902 ( .A(MixColumnsInput[24]), .B(MixColumnsOutput[24]), .S(n320), 
        .Z(RoundOutput[24]) );
  MUX2_X1 U903 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .B(
        MixColumnsOutput[25]), .S(n318), .Z(RoundOutput[25]) );
  MUX2_X1 U904 ( .A(MixColumnsInput[26]), .B(MixColumnsOutput[26]), .S(n316), 
        .Z(RoundOutput[26]) );
  MUX2_X1 U905 ( .A(MixColumnsInput[27]), .B(MixColumnsOutput[27]), .S(n317), 
        .Z(RoundOutput[27]) );
  MUX2_X1 U906 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .B(
        MixColumnsOutput[28]), .S(n315), .Z(RoundOutput[28]) );
  MUX2_X1 U907 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .B(
        MixColumnsOutput[29]), .S(n319), .Z(RoundOutput[29]) );
  MUX2_X1 U908 ( .A(MixColumnsInput[2]), .B(MixColumnsOutput[2]), .S(n315), 
        .Z(RoundOutput[2]) );
  MUX2_X1 U909 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .B(
        MixColumnsOutput[30]), .S(n320), .Z(RoundOutput[30]) );
  MUX2_X1 U910 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B(
        MixColumnsOutput[31]), .S(n318), .Z(RoundOutput[31]) );
  MUX2_X1 U911 ( .A(MixColumnsInput[32]), .B(MixColumnsOutput[32]), .S(n316), 
        .Z(RoundOutput[32]) );
  MUX2_X1 U912 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .B(
        MixColumnsOutput[33]), .S(n317), .Z(RoundOutput[33]) );
  MUX2_X1 U913 ( .A(MixColumnsInput[34]), .B(MixColumnsOutput[34]), .S(n315), 
        .Z(RoundOutput[34]) );
  MUX2_X1 U914 ( .A(MixColumnsInput[35]), .B(MixColumnsOutput[35]), .S(n320), 
        .Z(RoundOutput[35]) );
  MUX2_X1 U915 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B(
        MixColumnsOutput[36]), .S(n320), .Z(RoundOutput[36]) );
  MUX2_X1 U916 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B(
        MixColumnsOutput[37]), .S(n320), .Z(RoundOutput[37]) );
  MUX2_X1 U917 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B(
        MixColumnsOutput[38]), .S(n320), .Z(RoundOutput[38]) );
  MUX2_X1 U918 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsOutput[39]), .S(n320), .Z(RoundOutput[39]) );
  MUX2_X1 U919 ( .A(MixColumnsInput[3]), .B(MixColumnsOutput[3]), .S(n320), 
        .Z(RoundOutput[3]) );
  MUX2_X1 U920 ( .A(MixColumnsInput[40]), .B(MixColumnsOutput[40]), .S(n320), 
        .Z(RoundOutput[40]) );
  MUX2_X1 U921 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .B(
        MixColumnsOutput[41]), .S(n320), .Z(RoundOutput[41]) );
  MUX2_X1 U922 ( .A(MixColumnsInput[42]), .B(MixColumnsOutput[42]), .S(n320), 
        .Z(RoundOutput[42]) );
  MUX2_X1 U923 ( .A(MixColumnsInput[43]), .B(MixColumnsOutput[43]), .S(n320), 
        .Z(RoundOutput[43]) );
  MUX2_X1 U924 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .B(
        MixColumnsOutput[44]), .S(n320), .Z(RoundOutput[44]) );
  MUX2_X1 U925 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .B(
        MixColumnsOutput[45]), .S(n320), .Z(RoundOutput[45]) );
  MUX2_X1 U926 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .B(
        MixColumnsOutput[46]), .S(n319), .Z(RoundOutput[46]) );
  MUX2_X1 U927 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsOutput[47]), .S(n319), .Z(RoundOutput[47]) );
  MUX2_X1 U928 ( .A(MixColumnsInput[48]), .B(MixColumnsOutput[48]), .S(n319), 
        .Z(RoundOutput[48]) );
  MUX2_X1 U929 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .B(
        MixColumnsOutput[49]), .S(n319), .Z(RoundOutput[49]) );
  MUX2_X1 U930 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B(
        MixColumnsOutput[4]), .S(n319), .Z(RoundOutput[4]) );
  MUX2_X1 U931 ( .A(MixColumnsInput[50]), .B(MixColumnsOutput[50]), .S(n319), 
        .Z(RoundOutput[50]) );
  MUX2_X1 U932 ( .A(MixColumnsInput[51]), .B(MixColumnsOutput[51]), .S(n319), 
        .Z(RoundOutput[51]) );
  MUX2_X1 U933 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .B(
        MixColumnsOutput[52]), .S(n319), .Z(RoundOutput[52]) );
  MUX2_X1 U934 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .B(
        MixColumnsOutput[53]), .S(n319), .Z(RoundOutput[53]) );
  MUX2_X1 U935 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .B(
        MixColumnsOutput[54]), .S(n319), .Z(RoundOutput[54]) );
  MUX2_X1 U936 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B(
        MixColumnsOutput[55]), .S(n319), .Z(RoundOutput[55]) );
  MUX2_X1 U937 ( .A(MixColumnsInput[56]), .B(MixColumnsOutput[56]), .S(n319), 
        .Z(RoundOutput[56]) );
  MUX2_X1 U938 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .B(
        MixColumnsOutput[57]), .S(n318), .Z(RoundOutput[57]) );
  MUX2_X1 U939 ( .A(MixColumnsInput[58]), .B(MixColumnsOutput[58]), .S(n318), 
        .Z(RoundOutput[58]) );
  MUX2_X1 U940 ( .A(MixColumnsInput[59]), .B(MixColumnsOutput[59]), .S(n318), 
        .Z(RoundOutput[59]) );
  MUX2_X1 U941 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B(
        MixColumnsOutput[5]), .S(n318), .Z(RoundOutput[5]) );
  MUX2_X1 U942 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .B(
        MixColumnsOutput[60]), .S(n318), .Z(RoundOutput[60]) );
  MUX2_X1 U943 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .B(
        MixColumnsOutput[61]), .S(n318), .Z(RoundOutput[61]) );
  MUX2_X1 U944 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .B(
        MixColumnsOutput[62]), .S(n318), .Z(RoundOutput[62]) );
  MUX2_X1 U945 ( .A(MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B(
        MixColumnsOutput[63]), .S(n318), .Z(RoundOutput[63]) );
  MUX2_X1 U946 ( .A(MixColumnsInput[64]), .B(MixColumnsOutput[64]), .S(n318), 
        .Z(RoundOutput[64]) );
  MUX2_X1 U947 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .B(
        MixColumnsOutput[65]), .S(n318), .Z(RoundOutput[65]) );
  MUX2_X1 U948 ( .A(MixColumnsInput[66]), .B(MixColumnsOutput[66]), .S(n318), 
        .Z(RoundOutput[66]) );
  MUX2_X1 U949 ( .A(MixColumnsInput[67]), .B(MixColumnsOutput[67]), .S(n318), 
        .Z(RoundOutput[67]) );
  MUX2_X1 U950 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B(
        MixColumnsOutput[68]), .S(n317), .Z(RoundOutput[68]) );
  MUX2_X1 U951 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B(
        MixColumnsOutput[69]), .S(n317), .Z(RoundOutput[69]) );
  MUX2_X1 U952 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B(
        MixColumnsOutput[6]), .S(n317), .Z(RoundOutput[6]) );
  MUX2_X1 U953 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B(
        MixColumnsOutput[70]), .S(n317), .Z(RoundOutput[70]) );
  MUX2_X1 U954 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsOutput[71]), .S(n317), .Z(RoundOutput[71]) );
  MUX2_X1 U955 ( .A(MixColumnsInput[72]), .B(MixColumnsOutput[72]), .S(n317), 
        .Z(RoundOutput[72]) );
  MUX2_X1 U956 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .B(
        MixColumnsOutput[73]), .S(n317), .Z(RoundOutput[73]) );
  MUX2_X1 U957 ( .A(MixColumnsInput[74]), .B(MixColumnsOutput[74]), .S(n317), 
        .Z(RoundOutput[74]) );
  MUX2_X1 U958 ( .A(MixColumnsInput[75]), .B(MixColumnsOutput[75]), .S(n317), 
        .Z(RoundOutput[75]) );
  MUX2_X1 U959 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .B(
        MixColumnsOutput[76]), .S(n317), .Z(RoundOutput[76]) );
  MUX2_X1 U960 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .B(
        MixColumnsOutput[77]), .S(n317), .Z(RoundOutput[77]) );
  MUX2_X1 U961 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .B(
        MixColumnsOutput[78]), .S(n317), .Z(RoundOutput[78]) );
  MUX2_X1 U962 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsOutput[79]), .S(n316), .Z(RoundOutput[79]) );
  MUX2_X1 U963 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsOutput[7]), .S(n316), .Z(RoundOutput[7]) );
  MUX2_X1 U964 ( .A(MixColumnsInput[80]), .B(MixColumnsOutput[80]), .S(n316), 
        .Z(RoundOutput[80]) );
  MUX2_X1 U965 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .B(
        MixColumnsOutput[81]), .S(n316), .Z(RoundOutput[81]) );
  MUX2_X1 U966 ( .A(MixColumnsInput[82]), .B(MixColumnsOutput[82]), .S(n316), 
        .Z(RoundOutput[82]) );
  MUX2_X1 U967 ( .A(MixColumnsInput[83]), .B(MixColumnsOutput[83]), .S(n316), 
        .Z(RoundOutput[83]) );
  MUX2_X1 U968 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .B(
        MixColumnsOutput[84]), .S(n316), .Z(RoundOutput[84]) );
  MUX2_X1 U969 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .B(
        MixColumnsOutput[85]), .S(n316), .Z(RoundOutput[85]) );
  MUX2_X1 U970 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .B(
        MixColumnsOutput[86]), .S(n316), .Z(RoundOutput[86]) );
  MUX2_X1 U971 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B(
        MixColumnsOutput[87]), .S(n316), .Z(RoundOutput[87]) );
  MUX2_X1 U972 ( .A(MixColumnsInput[88]), .B(MixColumnsOutput[88]), .S(n316), 
        .Z(RoundOutput[88]) );
  MUX2_X1 U973 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .B(
        MixColumnsOutput[89]), .S(n316), .Z(RoundOutput[89]) );
  MUX2_X1 U974 ( .A(MixColumnsInput[8]), .B(MixColumnsOutput[8]), .S(n315), 
        .Z(RoundOutput[8]) );
  MUX2_X1 U975 ( .A(MixColumnsInput[90]), .B(MixColumnsOutput[90]), .S(n315), 
        .Z(RoundOutput[90]) );
  MUX2_X1 U976 ( .A(MixColumnsInput[91]), .B(MixColumnsOutput[91]), .S(n315), 
        .Z(RoundOutput[91]) );
  MUX2_X1 U977 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .B(
        MixColumnsOutput[92]), .S(n315), .Z(RoundOutput[92]) );
  MUX2_X1 U978 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .B(
        MixColumnsOutput[93]), .S(n315), .Z(RoundOutput[93]) );
  MUX2_X1 U979 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .B(
        MixColumnsOutput[94]), .S(n315), .Z(RoundOutput[94]) );
  MUX2_X1 U980 ( .A(MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B(
        MixColumnsOutput[95]), .S(n315), .Z(RoundOutput[95]) );
  MUX2_X1 U981 ( .A(MixColumnsInput[96]), .B(MixColumnsOutput[96]), .S(n315), 
        .Z(RoundOutput[96]) );
  MUX2_X1 U982 ( .A(MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .B(
        MixColumnsOutput[97]), .S(n315), .Z(RoundOutput[97]) );
  MUX2_X1 U983 ( .A(MixColumnsInput[98]), .B(MixColumnsOutput[98]), .S(n315), 
        .Z(RoundOutput[98]) );
  MUX2_X1 U984 ( .A(MixColumnsInput[99]), .B(MixColumnsOutput[99]), .S(n315), 
        .Z(RoundOutput[99]) );
  MUX2_X1 U985 ( .A(MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .B(
        MixColumnsOutput[9]), .S(n315), .Z(RoundOutput[9]) );
  XOR2_X1 U986 ( .A(RoundInput[0]), .B(RoundKey[0]), .Z(ciphertext[0]) );
  XOR2_X1 U987 ( .A(RoundInput[100]), .B(RoundKey[100]), .Z(ciphertext[100])
         );
  XOR2_X1 U988 ( .A(RoundInput[101]), .B(RoundKey[101]), .Z(ciphertext[101])
         );
  XOR2_X1 U989 ( .A(RoundInput[102]), .B(RoundKey[102]), .Z(ciphertext[102])
         );
  XOR2_X1 U990 ( .A(RoundInput[103]), .B(RoundKey[103]), .Z(ciphertext[103])
         );
  XOR2_X1 U991 ( .A(RoundInput[104]), .B(RoundKey[104]), .Z(ciphertext[104])
         );
  XOR2_X1 U992 ( .A(RoundInput[105]), .B(RoundKey[105]), .Z(ciphertext[105])
         );
  XOR2_X1 U993 ( .A(RoundInput[106]), .B(RoundKey[106]), .Z(ciphertext[106])
         );
  XOR2_X1 U994 ( .A(RoundInput[107]), .B(RoundKey[107]), .Z(ciphertext[107])
         );
  XOR2_X1 U995 ( .A(RoundInput[108]), .B(RoundKey[108]), .Z(ciphertext[108])
         );
  XOR2_X1 U996 ( .A(RoundInput[109]), .B(RoundKey[109]), .Z(ciphertext[109])
         );
  XOR2_X1 U997 ( .A(RoundInput[10]), .B(RoundKey[10]), .Z(ciphertext[10]) );
  XOR2_X1 U998 ( .A(RoundInput[110]), .B(RoundKey[110]), .Z(ciphertext[110])
         );
  XOR2_X1 U999 ( .A(RoundInput[111]), .B(RoundKey[111]), .Z(ciphertext[111])
         );
  XOR2_X1 U1000 ( .A(RoundInput[112]), .B(RoundKey[112]), .Z(ciphertext[112])
         );
  XOR2_X1 U1001 ( .A(RoundInput[113]), .B(RoundKey[113]), .Z(ciphertext[113])
         );
  XOR2_X1 U1002 ( .A(RoundInput[114]), .B(RoundKey[114]), .Z(ciphertext[114])
         );
  XOR2_X1 U1003 ( .A(RoundInput[115]), .B(RoundKey[115]), .Z(ciphertext[115])
         );
  XOR2_X1 U1004 ( .A(RoundInput[116]), .B(RoundKey[116]), .Z(ciphertext[116])
         );
  XOR2_X1 U1005 ( .A(RoundInput[117]), .B(RoundKey[117]), .Z(ciphertext[117])
         );
  XOR2_X1 U1006 ( .A(RoundInput[118]), .B(RoundKey[118]), .Z(ciphertext[118])
         );
  XOR2_X1 U1007 ( .A(RoundInput[119]), .B(RoundKey[119]), .Z(ciphertext[119])
         );
  XOR2_X1 U1008 ( .A(RoundInput[11]), .B(RoundKey[11]), .Z(ciphertext[11]) );
  XOR2_X1 U1009 ( .A(RoundInput[120]), .B(RoundKey[120]), .Z(ciphertext[120])
         );
  XOR2_X1 U1010 ( .A(RoundInput[121]), .B(RoundKey[121]), .Z(ciphertext[121])
         );
  XOR2_X1 U1011 ( .A(RoundInput[122]), .B(RoundKey[122]), .Z(ciphertext[122])
         );
  XOR2_X1 U1012 ( .A(RoundInput[123]), .B(RoundKey[123]), .Z(ciphertext[123])
         );
  XOR2_X1 U1013 ( .A(RoundInput[124]), .B(RoundKey[124]), .Z(ciphertext[124])
         );
  XOR2_X1 U1014 ( .A(RoundInput[125]), .B(RoundKey[125]), .Z(ciphertext[125])
         );
  XOR2_X1 U1015 ( .A(RoundInput[126]), .B(RoundKey[126]), .Z(ciphertext[126])
         );
  XOR2_X1 U1016 ( .A(RoundInput[127]), .B(RoundKey[127]), .Z(ciphertext[127])
         );
  XOR2_X1 U1017 ( .A(RoundInput[12]), .B(RoundKey[12]), .Z(ciphertext[12]) );
  XOR2_X1 U1018 ( .A(RoundInput[13]), .B(RoundKey[13]), .Z(ciphertext[13]) );
  XOR2_X1 U1019 ( .A(RoundInput[14]), .B(RoundKey[14]), .Z(ciphertext[14]) );
  XOR2_X1 U1020 ( .A(RoundInput[15]), .B(RoundKey[15]), .Z(ciphertext[15]) );
  XOR2_X1 U1021 ( .A(RoundInput[16]), .B(RoundKey[16]), .Z(ciphertext[16]) );
  XOR2_X1 U1022 ( .A(RoundInput[17]), .B(RoundKey[17]), .Z(ciphertext[17]) );
  XOR2_X1 U1023 ( .A(RoundInput[18]), .B(RoundKey[18]), .Z(ciphertext[18]) );
  XOR2_X1 U1024 ( .A(RoundInput[19]), .B(RoundKey[19]), .Z(ciphertext[19]) );
  XOR2_X1 U1025 ( .A(RoundInput[1]), .B(RoundKey[1]), .Z(ciphertext[1]) );
  XOR2_X1 U1026 ( .A(RoundInput[20]), .B(RoundKey[20]), .Z(ciphertext[20]) );
  XOR2_X1 U1027 ( .A(RoundInput[21]), .B(RoundKey[21]), .Z(ciphertext[21]) );
  XOR2_X1 U1028 ( .A(RoundInput[22]), .B(RoundKey[22]), .Z(ciphertext[22]) );
  XOR2_X1 U1029 ( .A(RoundInput[23]), .B(RoundKey[23]), .Z(ciphertext[23]) );
  XOR2_X1 U1030 ( .A(RoundInput[24]), .B(RoundKey[24]), .Z(ciphertext[24]) );
  XOR2_X1 U1031 ( .A(RoundInput[25]), .B(RoundKey[25]), .Z(ciphertext[25]) );
  XOR2_X1 U1032 ( .A(RoundInput[26]), .B(RoundKey[26]), .Z(ciphertext[26]) );
  XOR2_X1 U1033 ( .A(RoundInput[27]), .B(RoundKey[27]), .Z(ciphertext[27]) );
  XOR2_X1 U1034 ( .A(RoundInput[28]), .B(RoundKey[28]), .Z(ciphertext[28]) );
  XOR2_X1 U1035 ( .A(RoundInput[29]), .B(RoundKey[29]), .Z(ciphertext[29]) );
  XOR2_X1 U1036 ( .A(RoundInput[2]), .B(RoundKey[2]), .Z(ciphertext[2]) );
  XOR2_X1 U1037 ( .A(RoundInput[30]), .B(RoundKey[30]), .Z(ciphertext[30]) );
  XOR2_X1 U1038 ( .A(RoundInput[31]), .B(RoundKey[31]), .Z(ciphertext[31]) );
  XOR2_X1 U1039 ( .A(RoundInput[32]), .B(RoundKey[32]), .Z(ciphertext[32]) );
  XOR2_X1 U1040 ( .A(RoundInput[33]), .B(RoundKey[33]), .Z(ciphertext[33]) );
  XOR2_X1 U1041 ( .A(RoundInput[34]), .B(RoundKey[34]), .Z(ciphertext[34]) );
  XOR2_X1 U1042 ( .A(RoundInput[35]), .B(RoundKey[35]), .Z(ciphertext[35]) );
  XOR2_X1 U1043 ( .A(RoundInput[36]), .B(RoundKey[36]), .Z(ciphertext[36]) );
  XOR2_X1 U1044 ( .A(RoundInput[37]), .B(RoundKey[37]), .Z(ciphertext[37]) );
  XOR2_X1 U1045 ( .A(RoundInput[38]), .B(RoundKey[38]), .Z(ciphertext[38]) );
  XOR2_X1 U1046 ( .A(RoundInput[39]), .B(RoundKey[39]), .Z(ciphertext[39]) );
  XOR2_X1 U1047 ( .A(RoundInput[3]), .B(RoundKey[3]), .Z(ciphertext[3]) );
  XOR2_X1 U1048 ( .A(RoundInput[40]), .B(RoundKey[40]), .Z(ciphertext[40]) );
  XOR2_X1 U1049 ( .A(RoundInput[41]), .B(RoundKey[41]), .Z(ciphertext[41]) );
  XOR2_X1 U1050 ( .A(RoundInput[42]), .B(RoundKey[42]), .Z(ciphertext[42]) );
  XOR2_X1 U1051 ( .A(RoundInput[43]), .B(RoundKey[43]), .Z(ciphertext[43]) );
  XOR2_X1 U1052 ( .A(RoundInput[44]), .B(RoundKey[44]), .Z(ciphertext[44]) );
  XOR2_X1 U1053 ( .A(RoundInput[45]), .B(RoundKey[45]), .Z(ciphertext[45]) );
  XOR2_X1 U1054 ( .A(RoundInput[46]), .B(RoundKey[46]), .Z(ciphertext[46]) );
  XOR2_X1 U1055 ( .A(RoundInput[47]), .B(RoundKey[47]), .Z(ciphertext[47]) );
  XOR2_X1 U1056 ( .A(RoundInput[48]), .B(RoundKey[48]), .Z(ciphertext[48]) );
  XOR2_X1 U1057 ( .A(RoundInput[49]), .B(RoundKey[49]), .Z(ciphertext[49]) );
  XOR2_X1 U1058 ( .A(RoundInput[4]), .B(RoundKey[4]), .Z(ciphertext[4]) );
  XOR2_X1 U1059 ( .A(RoundInput[50]), .B(RoundKey[50]), .Z(ciphertext[50]) );
  XOR2_X1 U1060 ( .A(RoundInput[51]), .B(RoundKey[51]), .Z(ciphertext[51]) );
  XOR2_X1 U1061 ( .A(RoundInput[52]), .B(RoundKey[52]), .Z(ciphertext[52]) );
  XOR2_X1 U1062 ( .A(RoundInput[53]), .B(RoundKey[53]), .Z(ciphertext[53]) );
  XOR2_X1 U1063 ( .A(RoundInput[54]), .B(RoundKey[54]), .Z(ciphertext[54]) );
  XOR2_X1 U1064 ( .A(RoundInput[55]), .B(RoundKey[55]), .Z(ciphertext[55]) );
  XOR2_X1 U1065 ( .A(RoundInput[56]), .B(RoundKey[56]), .Z(ciphertext[56]) );
  XOR2_X1 U1066 ( .A(RoundInput[57]), .B(RoundKey[57]), .Z(ciphertext[57]) );
  XOR2_X1 U1067 ( .A(RoundInput[58]), .B(RoundKey[58]), .Z(ciphertext[58]) );
  XOR2_X1 U1068 ( .A(RoundInput[59]), .B(RoundKey[59]), .Z(ciphertext[59]) );
  XOR2_X1 U1069 ( .A(RoundInput[5]), .B(RoundKey[5]), .Z(ciphertext[5]) );
  XOR2_X1 U1070 ( .A(RoundInput[60]), .B(RoundKey[60]), .Z(ciphertext[60]) );
  XOR2_X1 U1071 ( .A(RoundInput[61]), .B(RoundKey[61]), .Z(ciphertext[61]) );
  XOR2_X1 U1072 ( .A(RoundInput[62]), .B(RoundKey[62]), .Z(ciphertext[62]) );
  XOR2_X1 U1073 ( .A(RoundInput[63]), .B(RoundKey[63]), .Z(ciphertext[63]) );
  XOR2_X1 U1074 ( .A(RoundInput[64]), .B(RoundKey[64]), .Z(ciphertext[64]) );
  XOR2_X1 U1075 ( .A(RoundInput[65]), .B(RoundKey[65]), .Z(ciphertext[65]) );
  XOR2_X1 U1076 ( .A(RoundInput[66]), .B(RoundKey[66]), .Z(ciphertext[66]) );
  XOR2_X1 U1077 ( .A(RoundInput[67]), .B(RoundKey[67]), .Z(ciphertext[67]) );
  XOR2_X1 U1078 ( .A(RoundInput[68]), .B(RoundKey[68]), .Z(ciphertext[68]) );
  XOR2_X1 U1079 ( .A(RoundInput[69]), .B(RoundKey[69]), .Z(ciphertext[69]) );
  XOR2_X1 U1080 ( .A(RoundInput[6]), .B(RoundKey[6]), .Z(ciphertext[6]) );
  XOR2_X1 U1081 ( .A(RoundInput[70]), .B(RoundKey[70]), .Z(ciphertext[70]) );
  XOR2_X1 U1082 ( .A(RoundInput[71]), .B(RoundKey[71]), .Z(ciphertext[71]) );
  XOR2_X1 U1083 ( .A(RoundInput[72]), .B(RoundKey[72]), .Z(ciphertext[72]) );
  XOR2_X1 U1084 ( .A(RoundInput[73]), .B(RoundKey[73]), .Z(ciphertext[73]) );
  XOR2_X1 U1085 ( .A(RoundInput[74]), .B(RoundKey[74]), .Z(ciphertext[74]) );
  XOR2_X1 U1086 ( .A(RoundInput[75]), .B(RoundKey[75]), .Z(ciphertext[75]) );
  XOR2_X1 U1087 ( .A(RoundInput[76]), .B(RoundKey[76]), .Z(ciphertext[76]) );
  XOR2_X1 U1088 ( .A(RoundInput[77]), .B(RoundKey[77]), .Z(ciphertext[77]) );
  XOR2_X1 U1089 ( .A(RoundInput[78]), .B(RoundKey[78]), .Z(ciphertext[78]) );
  XOR2_X1 U1090 ( .A(RoundInput[79]), .B(RoundKey[79]), .Z(ciphertext[79]) );
  XOR2_X1 U1091 ( .A(RoundInput[7]), .B(RoundKey[7]), .Z(ciphertext[7]) );
  XOR2_X1 U1092 ( .A(RoundInput[80]), .B(RoundKey[80]), .Z(ciphertext[80]) );
  XOR2_X1 U1093 ( .A(RoundInput[81]), .B(RoundKey[81]), .Z(ciphertext[81]) );
  XOR2_X1 U1094 ( .A(RoundInput[82]), .B(RoundKey[82]), .Z(ciphertext[82]) );
  XOR2_X1 U1095 ( .A(RoundInput[83]), .B(RoundKey[83]), .Z(ciphertext[83]) );
  XOR2_X1 U1096 ( .A(RoundInput[84]), .B(RoundKey[84]), .Z(ciphertext[84]) );
  XOR2_X1 U1097 ( .A(RoundInput[85]), .B(RoundKey[85]), .Z(ciphertext[85]) );
  XOR2_X1 U1098 ( .A(RoundInput[86]), .B(RoundKey[86]), .Z(ciphertext[86]) );
  XOR2_X1 U1099 ( .A(RoundInput[87]), .B(RoundKey[87]), .Z(ciphertext[87]) );
  XOR2_X1 U1100 ( .A(RoundInput[88]), .B(RoundKey[88]), .Z(ciphertext[88]) );
  XOR2_X1 U1101 ( .A(RoundInput[89]), .B(RoundKey[89]), .Z(ciphertext[89]) );
  XOR2_X1 U1102 ( .A(RoundInput[8]), .B(RoundKey[8]), .Z(ciphertext[8]) );
  XOR2_X1 U1103 ( .A(RoundInput[90]), .B(RoundKey[90]), .Z(ciphertext[90]) );
  XOR2_X1 U1104 ( .A(RoundInput[91]), .B(RoundKey[91]), .Z(ciphertext[91]) );
  XOR2_X1 U1105 ( .A(RoundInput[92]), .B(RoundKey[92]), .Z(ciphertext[92]) );
  XOR2_X1 U1106 ( .A(RoundInput[93]), .B(RoundKey[93]), .Z(ciphertext[93]) );
  XOR2_X1 U1107 ( .A(RoundInput[94]), .B(RoundKey[94]), .Z(ciphertext[94]) );
  XOR2_X1 U1108 ( .A(RoundInput[95]), .B(RoundKey[95]), .Z(ciphertext[95]) );
  XOR2_X1 U1109 ( .A(RoundInput[96]), .B(RoundKey[96]), .Z(ciphertext[96]) );
  XOR2_X1 U1110 ( .A(RoundInput[97]), .B(RoundKey[97]), .Z(ciphertext[97]) );
  XOR2_X1 U1111 ( .A(RoundInput[98]), .B(RoundKey[98]), .Z(ciphertext[98]) );
  XOR2_X1 U1112 ( .A(RoundInput[99]), .B(RoundKey[99]), .Z(ciphertext[99]) );
  XOR2_X1 U1113 ( .A(RoundInput[9]), .B(RoundKey[9]), .Z(ciphertext[9]) );
  NAND2_X1 U1114 ( .A1(RoundCounter[3]), .A2(n333), .ZN(n334) );
  NOR2_X1 U1115 ( .A1(RoundCounter[0]), .A2(n334), .ZN(done) );
  INV_X1 U1116 ( .A(n335), .ZN(n336) );
  NAND2_X1 U1117 ( .A1(RoundCounter[2]), .A2(RoundCounter[1]), .ZN(n338) );
  NOR2_X1 U1118 ( .A1(n336), .A2(n338), .ZN(n283) );
  INV_X1 U1119 ( .A(n337), .ZN(n339) );
  NOR2_X1 U1120 ( .A1(n339), .A2(n338), .ZN(n285) );
  MUX2_X1 RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .A(RoundOutput[0]), .B(
        plaintext[0]), .S(reset), .Z(RoundReg_Inst_ff_SDE_0_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_0_current_state_reg_U1 ( .A(RoundInput[0]), .ZN(
        RoundReg_Inst_ff_SDE_0_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_0_next_state), .CK(clk), .Q(RoundInput[0]), .QN()
         );
  MUX2_X1 RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .A(RoundOutput[1]), .B(
        plaintext[1]), .S(reset), .Z(RoundReg_Inst_ff_SDE_1_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_1_current_state_reg_U1 ( .A(RoundInput[1]), .ZN(
        RoundReg_Inst_ff_SDE_1_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_1_next_state), .CK(clk), .Q(RoundInput[1]), .QN()
         );
  MUX2_X1 RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .A(RoundOutput[2]), .B(
        plaintext[2]), .S(reset), .Z(RoundReg_Inst_ff_SDE_2_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_2_current_state_reg_U1 ( .A(RoundInput[2]), .ZN(
        RoundReg_Inst_ff_SDE_2_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_2_next_state), .CK(clk), .Q(RoundInput[2]), .QN()
         );
  MUX2_X1 RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .A(RoundOutput[3]), .B(
        plaintext[3]), .S(reset), .Z(RoundReg_Inst_ff_SDE_3_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_3_current_state_reg_U1 ( .A(RoundInput[3]), .ZN(
        RoundReg_Inst_ff_SDE_3_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_3_next_state), .CK(clk), .Q(RoundInput[3]), .QN()
         );
  MUX2_X1 RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .A(RoundOutput[4]), .B(
        plaintext[4]), .S(reset), .Z(RoundReg_Inst_ff_SDE_4_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_4_current_state_reg_U1 ( .A(RoundInput[4]), .ZN(
        RoundReg_Inst_ff_SDE_4_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_4_next_state), .CK(clk), .Q(RoundInput[4]), .QN()
         );
  MUX2_X1 RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .A(RoundOutput[5]), .B(
        plaintext[5]), .S(reset), .Z(RoundReg_Inst_ff_SDE_5_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_5_current_state_reg_U1 ( .A(RoundInput[5]), .ZN(
        RoundReg_Inst_ff_SDE_5_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_5_next_state), .CK(clk), .Q(RoundInput[5]), .QN()
         );
  MUX2_X1 RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .A(RoundOutput[6]), .B(
        plaintext[6]), .S(reset), .Z(RoundReg_Inst_ff_SDE_6_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_6_current_state_reg_U1 ( .A(RoundInput[6]), .ZN(
        RoundReg_Inst_ff_SDE_6_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_6_next_state), .CK(clk), .Q(RoundInput[6]), .QN()
         );
  MUX2_X1 RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .A(RoundOutput[7]), .B(
        plaintext[7]), .S(reset), .Z(RoundReg_Inst_ff_SDE_7_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_7_current_state_reg_U1 ( .A(RoundInput[7]), .ZN(
        RoundReg_Inst_ff_SDE_7_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_7_next_state), .CK(clk), .Q(RoundInput[7]), .QN()
         );
  MUX2_X1 RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .A(RoundOutput[8]), .B(
        plaintext[8]), .S(reset), .Z(RoundReg_Inst_ff_SDE_8_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_8_current_state_reg_U1 ( .A(RoundInput[8]), .ZN(
        RoundReg_Inst_ff_SDE_8_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_8_next_state), .CK(clk), .Q(RoundInput[8]), .QN()
         );
  MUX2_X1 RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .A(RoundOutput[9]), .B(
        plaintext[9]), .S(reset), .Z(RoundReg_Inst_ff_SDE_9_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_9_current_state_reg_U1 ( .A(RoundInput[9]), .ZN(
        RoundReg_Inst_ff_SDE_9_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_9_next_state), .CK(clk), .Q(RoundInput[9]), .QN()
         );
  MUX2_X1 RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .A(RoundOutput[10]), .B(
        plaintext[10]), .S(reset), .Z(RoundReg_Inst_ff_SDE_10_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_10_current_state_reg_U1 ( .A(RoundInput[10]), 
        .ZN(RoundReg_Inst_ff_SDE_10_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_10_next_state), .CK(clk), .Q(RoundInput[10]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .A(RoundOutput[11]), .B(
        plaintext[11]), .S(reset), .Z(RoundReg_Inst_ff_SDE_11_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_11_current_state_reg_U1 ( .A(RoundInput[11]), 
        .ZN(RoundReg_Inst_ff_SDE_11_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_11_next_state), .CK(clk), .Q(RoundInput[11]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .A(RoundOutput[12]), .B(
        plaintext[12]), .S(reset), .Z(RoundReg_Inst_ff_SDE_12_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_12_current_state_reg_U1 ( .A(RoundInput[12]), 
        .ZN(RoundReg_Inst_ff_SDE_12_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_12_next_state), .CK(clk), .Q(RoundInput[12]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .A(RoundOutput[13]), .B(
        plaintext[13]), .S(reset), .Z(RoundReg_Inst_ff_SDE_13_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_13_current_state_reg_U1 ( .A(RoundInput[13]), 
        .ZN(RoundReg_Inst_ff_SDE_13_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_13_next_state), .CK(clk), .Q(RoundInput[13]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .A(RoundOutput[14]), .B(
        plaintext[14]), .S(reset), .Z(RoundReg_Inst_ff_SDE_14_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_14_current_state_reg_U1 ( .A(RoundInput[14]), 
        .ZN(RoundReg_Inst_ff_SDE_14_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_14_next_state), .CK(clk), .Q(RoundInput[14]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .A(RoundOutput[15]), .B(
        plaintext[15]), .S(reset), .Z(RoundReg_Inst_ff_SDE_15_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_15_current_state_reg_U1 ( .A(RoundInput[15]), 
        .ZN(RoundReg_Inst_ff_SDE_15_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_15_next_state), .CK(clk), .Q(RoundInput[15]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .A(RoundOutput[16]), .B(
        plaintext[16]), .S(reset), .Z(RoundReg_Inst_ff_SDE_16_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_16_current_state_reg_U1 ( .A(RoundInput[16]), 
        .ZN(RoundReg_Inst_ff_SDE_16_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_16_next_state), .CK(clk), .Q(RoundInput[16]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .A(RoundOutput[17]), .B(
        plaintext[17]), .S(reset), .Z(RoundReg_Inst_ff_SDE_17_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_17_current_state_reg_U1 ( .A(RoundInput[17]), 
        .ZN(RoundReg_Inst_ff_SDE_17_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_17_next_state), .CK(clk), .Q(RoundInput[17]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .A(RoundOutput[18]), .B(
        plaintext[18]), .S(reset), .Z(RoundReg_Inst_ff_SDE_18_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_18_current_state_reg_U1 ( .A(RoundInput[18]), 
        .ZN(RoundReg_Inst_ff_SDE_18_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_18_next_state), .CK(clk), .Q(RoundInput[18]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .A(RoundOutput[19]), .B(
        plaintext[19]), .S(reset), .Z(RoundReg_Inst_ff_SDE_19_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_19_current_state_reg_U1 ( .A(RoundInput[19]), 
        .ZN(RoundReg_Inst_ff_SDE_19_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_19_next_state), .CK(clk), .Q(RoundInput[19]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .A(RoundOutput[20]), .B(
        plaintext[20]), .S(reset), .Z(RoundReg_Inst_ff_SDE_20_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_20_current_state_reg_U1 ( .A(RoundInput[20]), 
        .ZN(RoundReg_Inst_ff_SDE_20_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_20_next_state), .CK(clk), .Q(RoundInput[20]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .A(RoundOutput[21]), .B(
        plaintext[21]), .S(reset), .Z(RoundReg_Inst_ff_SDE_21_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_21_current_state_reg_U1 ( .A(RoundInput[21]), 
        .ZN(RoundReg_Inst_ff_SDE_21_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_21_next_state), .CK(clk), .Q(RoundInput[21]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .A(RoundOutput[22]), .B(
        plaintext[22]), .S(reset), .Z(RoundReg_Inst_ff_SDE_22_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_22_current_state_reg_U1 ( .A(RoundInput[22]), 
        .ZN(RoundReg_Inst_ff_SDE_22_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_22_next_state), .CK(clk), .Q(RoundInput[22]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .A(RoundOutput[23]), .B(
        plaintext[23]), .S(reset), .Z(RoundReg_Inst_ff_SDE_23_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_23_current_state_reg_U1 ( .A(RoundInput[23]), 
        .ZN(RoundReg_Inst_ff_SDE_23_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_23_next_state), .CK(clk), .Q(RoundInput[23]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .A(RoundOutput[24]), .B(
        plaintext[24]), .S(reset), .Z(RoundReg_Inst_ff_SDE_24_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_24_current_state_reg_U1 ( .A(RoundInput[24]), 
        .ZN(RoundReg_Inst_ff_SDE_24_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_24_next_state), .CK(clk), .Q(RoundInput[24]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .A(RoundOutput[25]), .B(
        plaintext[25]), .S(reset), .Z(RoundReg_Inst_ff_SDE_25_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_25_current_state_reg_U1 ( .A(RoundInput[25]), 
        .ZN(RoundReg_Inst_ff_SDE_25_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_25_next_state), .CK(clk), .Q(RoundInput[25]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .A(RoundOutput[26]), .B(
        plaintext[26]), .S(reset), .Z(RoundReg_Inst_ff_SDE_26_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_26_current_state_reg_U1 ( .A(RoundInput[26]), 
        .ZN(RoundReg_Inst_ff_SDE_26_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_26_next_state), .CK(clk), .Q(RoundInput[26]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .A(RoundOutput[27]), .B(
        plaintext[27]), .S(reset), .Z(RoundReg_Inst_ff_SDE_27_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_27_current_state_reg_U1 ( .A(RoundInput[27]), 
        .ZN(RoundReg_Inst_ff_SDE_27_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_27_next_state), .CK(clk), .Q(RoundInput[27]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .A(RoundOutput[28]), .B(
        plaintext[28]), .S(reset), .Z(RoundReg_Inst_ff_SDE_28_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_28_current_state_reg_U1 ( .A(RoundInput[28]), 
        .ZN(RoundReg_Inst_ff_SDE_28_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_28_next_state), .CK(clk), .Q(RoundInput[28]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .A(RoundOutput[29]), .B(
        plaintext[29]), .S(reset), .Z(RoundReg_Inst_ff_SDE_29_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_29_current_state_reg_U1 ( .A(RoundInput[29]), 
        .ZN(RoundReg_Inst_ff_SDE_29_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_29_next_state), .CK(clk), .Q(RoundInput[29]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .A(RoundOutput[30]), .B(
        plaintext[30]), .S(reset), .Z(RoundReg_Inst_ff_SDE_30_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_30_current_state_reg_U1 ( .A(RoundInput[30]), 
        .ZN(RoundReg_Inst_ff_SDE_30_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_30_next_state), .CK(clk), .Q(RoundInput[30]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .A(RoundOutput[31]), .B(
        plaintext[31]), .S(reset), .Z(RoundReg_Inst_ff_SDE_31_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_31_current_state_reg_U1 ( .A(RoundInput[31]), 
        .ZN(RoundReg_Inst_ff_SDE_31_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_31_next_state), .CK(clk), .Q(RoundInput[31]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .A(RoundOutput[32]), .B(
        plaintext[32]), .S(reset), .Z(RoundReg_Inst_ff_SDE_32_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_32_current_state_reg_U1 ( .A(RoundInput[32]), 
        .ZN(RoundReg_Inst_ff_SDE_32_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_32_next_state), .CK(clk), .Q(RoundInput[32]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .A(RoundOutput[33]), .B(
        plaintext[33]), .S(reset), .Z(RoundReg_Inst_ff_SDE_33_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_33_current_state_reg_U1 ( .A(RoundInput[33]), 
        .ZN(RoundReg_Inst_ff_SDE_33_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_33_next_state), .CK(clk), .Q(RoundInput[33]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .A(RoundOutput[34]), .B(
        plaintext[34]), .S(reset), .Z(RoundReg_Inst_ff_SDE_34_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_34_current_state_reg_U1 ( .A(RoundInput[34]), 
        .ZN(RoundReg_Inst_ff_SDE_34_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_34_next_state), .CK(clk), .Q(RoundInput[34]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .A(RoundOutput[35]), .B(
        plaintext[35]), .S(reset), .Z(RoundReg_Inst_ff_SDE_35_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_35_current_state_reg_U1 ( .A(RoundInput[35]), 
        .ZN(RoundReg_Inst_ff_SDE_35_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_35_next_state), .CK(clk), .Q(RoundInput[35]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .A(RoundOutput[36]), .B(
        plaintext[36]), .S(reset), .Z(RoundReg_Inst_ff_SDE_36_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_36_current_state_reg_U1 ( .A(RoundInput[36]), 
        .ZN(RoundReg_Inst_ff_SDE_36_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_36_next_state), .CK(clk), .Q(RoundInput[36]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .A(RoundOutput[37]), .B(
        plaintext[37]), .S(reset), .Z(RoundReg_Inst_ff_SDE_37_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_37_current_state_reg_U1 ( .A(RoundInput[37]), 
        .ZN(RoundReg_Inst_ff_SDE_37_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_37_next_state), .CK(clk), .Q(RoundInput[37]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .A(RoundOutput[38]), .B(
        plaintext[38]), .S(reset), .Z(RoundReg_Inst_ff_SDE_38_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_38_current_state_reg_U1 ( .A(RoundInput[38]), 
        .ZN(RoundReg_Inst_ff_SDE_38_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_38_next_state), .CK(clk), .Q(RoundInput[38]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .A(RoundOutput[39]), .B(
        plaintext[39]), .S(reset), .Z(RoundReg_Inst_ff_SDE_39_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_39_current_state_reg_U1 ( .A(RoundInput[39]), 
        .ZN(RoundReg_Inst_ff_SDE_39_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_39_next_state), .CK(clk), .Q(RoundInput[39]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .A(RoundOutput[40]), .B(
        plaintext[40]), .S(reset), .Z(RoundReg_Inst_ff_SDE_40_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_40_current_state_reg_U1 ( .A(RoundInput[40]), 
        .ZN(RoundReg_Inst_ff_SDE_40_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_40_next_state), .CK(clk), .Q(RoundInput[40]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .A(RoundOutput[41]), .B(
        plaintext[41]), .S(reset), .Z(RoundReg_Inst_ff_SDE_41_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_41_current_state_reg_U1 ( .A(RoundInput[41]), 
        .ZN(RoundReg_Inst_ff_SDE_41_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_41_next_state), .CK(clk), .Q(RoundInput[41]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .A(RoundOutput[42]), .B(
        plaintext[42]), .S(reset), .Z(RoundReg_Inst_ff_SDE_42_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_42_current_state_reg_U1 ( .A(RoundInput[42]), 
        .ZN(RoundReg_Inst_ff_SDE_42_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_42_next_state), .CK(clk), .Q(RoundInput[42]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .A(RoundOutput[43]), .B(
        plaintext[43]), .S(reset), .Z(RoundReg_Inst_ff_SDE_43_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_43_current_state_reg_U1 ( .A(RoundInput[43]), 
        .ZN(RoundReg_Inst_ff_SDE_43_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_43_next_state), .CK(clk), .Q(RoundInput[43]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .A(RoundOutput[44]), .B(
        plaintext[44]), .S(reset), .Z(RoundReg_Inst_ff_SDE_44_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_44_current_state_reg_U1 ( .A(RoundInput[44]), 
        .ZN(RoundReg_Inst_ff_SDE_44_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_44_next_state), .CK(clk), .Q(RoundInput[44]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .A(RoundOutput[45]), .B(
        plaintext[45]), .S(reset), .Z(RoundReg_Inst_ff_SDE_45_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_45_current_state_reg_U1 ( .A(RoundInput[45]), 
        .ZN(RoundReg_Inst_ff_SDE_45_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_45_next_state), .CK(clk), .Q(RoundInput[45]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .A(RoundOutput[46]), .B(
        plaintext[46]), .S(reset), .Z(RoundReg_Inst_ff_SDE_46_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_46_current_state_reg_U1 ( .A(RoundInput[46]), 
        .ZN(RoundReg_Inst_ff_SDE_46_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_46_next_state), .CK(clk), .Q(RoundInput[46]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .A(RoundOutput[47]), .B(
        plaintext[47]), .S(reset), .Z(RoundReg_Inst_ff_SDE_47_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_47_current_state_reg_U1 ( .A(RoundInput[47]), 
        .ZN(RoundReg_Inst_ff_SDE_47_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_47_next_state), .CK(clk), .Q(RoundInput[47]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .A(RoundOutput[48]), .B(
        plaintext[48]), .S(reset), .Z(RoundReg_Inst_ff_SDE_48_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_48_current_state_reg_U1 ( .A(RoundInput[48]), 
        .ZN(RoundReg_Inst_ff_SDE_48_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_48_next_state), .CK(clk), .Q(RoundInput[48]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .A(RoundOutput[49]), .B(
        plaintext[49]), .S(reset), .Z(RoundReg_Inst_ff_SDE_49_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_49_current_state_reg_U1 ( .A(RoundInput[49]), 
        .ZN(RoundReg_Inst_ff_SDE_49_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_49_next_state), .CK(clk), .Q(RoundInput[49]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .A(RoundOutput[50]), .B(
        plaintext[50]), .S(reset), .Z(RoundReg_Inst_ff_SDE_50_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_50_current_state_reg_U1 ( .A(RoundInput[50]), 
        .ZN(RoundReg_Inst_ff_SDE_50_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_50_next_state), .CK(clk), .Q(RoundInput[50]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .A(RoundOutput[51]), .B(
        plaintext[51]), .S(reset), .Z(RoundReg_Inst_ff_SDE_51_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_51_current_state_reg_U1 ( .A(RoundInput[51]), 
        .ZN(RoundReg_Inst_ff_SDE_51_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_51_next_state), .CK(clk), .Q(RoundInput[51]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .A(RoundOutput[52]), .B(
        plaintext[52]), .S(reset), .Z(RoundReg_Inst_ff_SDE_52_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_52_current_state_reg_U1 ( .A(RoundInput[52]), 
        .ZN(RoundReg_Inst_ff_SDE_52_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_52_next_state), .CK(clk), .Q(RoundInput[52]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .A(RoundOutput[53]), .B(
        plaintext[53]), .S(reset), .Z(RoundReg_Inst_ff_SDE_53_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_53_current_state_reg_U1 ( .A(RoundInput[53]), 
        .ZN(RoundReg_Inst_ff_SDE_53_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_53_next_state), .CK(clk), .Q(RoundInput[53]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .A(RoundOutput[54]), .B(
        plaintext[54]), .S(reset), .Z(RoundReg_Inst_ff_SDE_54_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_54_current_state_reg_U1 ( .A(RoundInput[54]), 
        .ZN(RoundReg_Inst_ff_SDE_54_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_54_next_state), .CK(clk), .Q(RoundInput[54]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .A(RoundOutput[55]), .B(
        plaintext[55]), .S(reset), .Z(RoundReg_Inst_ff_SDE_55_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_55_current_state_reg_U1 ( .A(RoundInput[55]), 
        .ZN(RoundReg_Inst_ff_SDE_55_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_55_next_state), .CK(clk), .Q(RoundInput[55]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .A(RoundOutput[56]), .B(
        plaintext[56]), .S(reset), .Z(RoundReg_Inst_ff_SDE_56_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_56_current_state_reg_U1 ( .A(RoundInput[56]), 
        .ZN(RoundReg_Inst_ff_SDE_56_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_56_next_state), .CK(clk), .Q(RoundInput[56]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .A(RoundOutput[57]), .B(
        plaintext[57]), .S(reset), .Z(RoundReg_Inst_ff_SDE_57_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_57_current_state_reg_U1 ( .A(RoundInput[57]), 
        .ZN(RoundReg_Inst_ff_SDE_57_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_57_next_state), .CK(clk), .Q(RoundInput[57]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .A(RoundOutput[58]), .B(
        plaintext[58]), .S(reset), .Z(RoundReg_Inst_ff_SDE_58_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_58_current_state_reg_U1 ( .A(RoundInput[58]), 
        .ZN(RoundReg_Inst_ff_SDE_58_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_58_next_state), .CK(clk), .Q(RoundInput[58]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .A(RoundOutput[59]), .B(
        plaintext[59]), .S(reset), .Z(RoundReg_Inst_ff_SDE_59_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_59_current_state_reg_U1 ( .A(RoundInput[59]), 
        .ZN(RoundReg_Inst_ff_SDE_59_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_59_next_state), .CK(clk), .Q(RoundInput[59]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .A(RoundOutput[60]), .B(
        plaintext[60]), .S(reset), .Z(RoundReg_Inst_ff_SDE_60_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_60_current_state_reg_U1 ( .A(RoundInput[60]), 
        .ZN(RoundReg_Inst_ff_SDE_60_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_60_next_state), .CK(clk), .Q(RoundInput[60]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .A(RoundOutput[61]), .B(
        plaintext[61]), .S(reset), .Z(RoundReg_Inst_ff_SDE_61_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_61_current_state_reg_U1 ( .A(RoundInput[61]), 
        .ZN(RoundReg_Inst_ff_SDE_61_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_61_next_state), .CK(clk), .Q(RoundInput[61]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .A(RoundOutput[62]), .B(
        plaintext[62]), .S(reset), .Z(RoundReg_Inst_ff_SDE_62_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_62_current_state_reg_U1 ( .A(RoundInput[62]), 
        .ZN(RoundReg_Inst_ff_SDE_62_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_62_next_state), .CK(clk), .Q(RoundInput[62]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .A(RoundOutput[63]), .B(
        plaintext[63]), .S(reset), .Z(RoundReg_Inst_ff_SDE_63_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_63_current_state_reg_U1 ( .A(RoundInput[63]), 
        .ZN(RoundReg_Inst_ff_SDE_63_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_63_next_state), .CK(clk), .Q(RoundInput[63]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .A(RoundOutput[64]), .B(
        plaintext[64]), .S(reset), .Z(RoundReg_Inst_ff_SDE_64_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_64_current_state_reg_U1 ( .A(RoundInput[64]), 
        .ZN(RoundReg_Inst_ff_SDE_64_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_64_next_state), .CK(clk), .Q(RoundInput[64]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .A(RoundOutput[65]), .B(
        plaintext[65]), .S(reset), .Z(RoundReg_Inst_ff_SDE_65_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_65_current_state_reg_U1 ( .A(RoundInput[65]), 
        .ZN(RoundReg_Inst_ff_SDE_65_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_65_next_state), .CK(clk), .Q(RoundInput[65]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .A(RoundOutput[66]), .B(
        plaintext[66]), .S(reset), .Z(RoundReg_Inst_ff_SDE_66_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_66_current_state_reg_U1 ( .A(RoundInput[66]), 
        .ZN(RoundReg_Inst_ff_SDE_66_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_66_next_state), .CK(clk), .Q(RoundInput[66]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .A(RoundOutput[67]), .B(
        plaintext[67]), .S(reset), .Z(RoundReg_Inst_ff_SDE_67_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_67_current_state_reg_U1 ( .A(RoundInput[67]), 
        .ZN(RoundReg_Inst_ff_SDE_67_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_67_next_state), .CK(clk), .Q(RoundInput[67]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .A(RoundOutput[68]), .B(
        plaintext[68]), .S(reset), .Z(RoundReg_Inst_ff_SDE_68_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_68_current_state_reg_U1 ( .A(RoundInput[68]), 
        .ZN(RoundReg_Inst_ff_SDE_68_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_68_next_state), .CK(clk), .Q(RoundInput[68]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .A(RoundOutput[69]), .B(
        plaintext[69]), .S(reset), .Z(RoundReg_Inst_ff_SDE_69_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_69_current_state_reg_U1 ( .A(RoundInput[69]), 
        .ZN(RoundReg_Inst_ff_SDE_69_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_69_next_state), .CK(clk), .Q(RoundInput[69]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .A(RoundOutput[70]), .B(
        plaintext[70]), .S(reset), .Z(RoundReg_Inst_ff_SDE_70_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_70_current_state_reg_U1 ( .A(RoundInput[70]), 
        .ZN(RoundReg_Inst_ff_SDE_70_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_70_next_state), .CK(clk), .Q(RoundInput[70]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .A(RoundOutput[71]), .B(
        plaintext[71]), .S(reset), .Z(RoundReg_Inst_ff_SDE_71_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_71_current_state_reg_U1 ( .A(RoundInput[71]), 
        .ZN(RoundReg_Inst_ff_SDE_71_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_71_next_state), .CK(clk), .Q(RoundInput[71]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .A(RoundOutput[72]), .B(
        plaintext[72]), .S(reset), .Z(RoundReg_Inst_ff_SDE_72_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_72_current_state_reg_U1 ( .A(RoundInput[72]), 
        .ZN(RoundReg_Inst_ff_SDE_72_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_72_next_state), .CK(clk), .Q(RoundInput[72]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .A(RoundOutput[73]), .B(
        plaintext[73]), .S(reset), .Z(RoundReg_Inst_ff_SDE_73_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_73_current_state_reg_U1 ( .A(RoundInput[73]), 
        .ZN(RoundReg_Inst_ff_SDE_73_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_73_next_state), .CK(clk), .Q(RoundInput[73]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .A(RoundOutput[74]), .B(
        plaintext[74]), .S(reset), .Z(RoundReg_Inst_ff_SDE_74_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_74_current_state_reg_U1 ( .A(RoundInput[74]), 
        .ZN(RoundReg_Inst_ff_SDE_74_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_74_next_state), .CK(clk), .Q(RoundInput[74]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .A(RoundOutput[75]), .B(
        plaintext[75]), .S(reset), .Z(RoundReg_Inst_ff_SDE_75_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_75_current_state_reg_U1 ( .A(RoundInput[75]), 
        .ZN(RoundReg_Inst_ff_SDE_75_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_75_next_state), .CK(clk), .Q(RoundInput[75]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .A(RoundOutput[76]), .B(
        plaintext[76]), .S(reset), .Z(RoundReg_Inst_ff_SDE_76_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_76_current_state_reg_U1 ( .A(RoundInput[76]), 
        .ZN(RoundReg_Inst_ff_SDE_76_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_76_next_state), .CK(clk), .Q(RoundInput[76]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .A(RoundOutput[77]), .B(
        plaintext[77]), .S(reset), .Z(RoundReg_Inst_ff_SDE_77_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_77_current_state_reg_U1 ( .A(RoundInput[77]), 
        .ZN(RoundReg_Inst_ff_SDE_77_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_77_next_state), .CK(clk), .Q(RoundInput[77]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .A(RoundOutput[78]), .B(
        plaintext[78]), .S(reset), .Z(RoundReg_Inst_ff_SDE_78_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_78_current_state_reg_U1 ( .A(RoundInput[78]), 
        .ZN(RoundReg_Inst_ff_SDE_78_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_78_next_state), .CK(clk), .Q(RoundInput[78]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .A(RoundOutput[79]), .B(
        plaintext[79]), .S(reset), .Z(RoundReg_Inst_ff_SDE_79_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_79_current_state_reg_U1 ( .A(RoundInput[79]), 
        .ZN(RoundReg_Inst_ff_SDE_79_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_79_next_state), .CK(clk), .Q(RoundInput[79]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .A(RoundOutput[80]), .B(
        plaintext[80]), .S(reset), .Z(RoundReg_Inst_ff_SDE_80_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_80_current_state_reg_U1 ( .A(RoundInput[80]), 
        .ZN(RoundReg_Inst_ff_SDE_80_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_80_next_state), .CK(clk), .Q(RoundInput[80]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .A(RoundOutput[81]), .B(
        plaintext[81]), .S(reset), .Z(RoundReg_Inst_ff_SDE_81_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_81_current_state_reg_U1 ( .A(RoundInput[81]), 
        .ZN(RoundReg_Inst_ff_SDE_81_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_81_next_state), .CK(clk), .Q(RoundInput[81]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .A(RoundOutput[82]), .B(
        plaintext[82]), .S(reset), .Z(RoundReg_Inst_ff_SDE_82_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_82_current_state_reg_U1 ( .A(RoundInput[82]), 
        .ZN(RoundReg_Inst_ff_SDE_82_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_82_next_state), .CK(clk), .Q(RoundInput[82]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .A(RoundOutput[83]), .B(
        plaintext[83]), .S(reset), .Z(RoundReg_Inst_ff_SDE_83_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_83_current_state_reg_U1 ( .A(RoundInput[83]), 
        .ZN(RoundReg_Inst_ff_SDE_83_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_83_next_state), .CK(clk), .Q(RoundInput[83]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .A(RoundOutput[84]), .B(
        plaintext[84]), .S(reset), .Z(RoundReg_Inst_ff_SDE_84_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_84_current_state_reg_U1 ( .A(RoundInput[84]), 
        .ZN(RoundReg_Inst_ff_SDE_84_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_84_next_state), .CK(clk), .Q(RoundInput[84]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .A(RoundOutput[85]), .B(
        plaintext[85]), .S(reset), .Z(RoundReg_Inst_ff_SDE_85_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_85_current_state_reg_U1 ( .A(RoundInput[85]), 
        .ZN(RoundReg_Inst_ff_SDE_85_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_85_next_state), .CK(clk), .Q(RoundInput[85]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .A(RoundOutput[86]), .B(
        plaintext[86]), .S(reset), .Z(RoundReg_Inst_ff_SDE_86_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_86_current_state_reg_U1 ( .A(RoundInput[86]), 
        .ZN(RoundReg_Inst_ff_SDE_86_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_86_next_state), .CK(clk), .Q(RoundInput[86]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .A(RoundOutput[87]), .B(
        plaintext[87]), .S(reset), .Z(RoundReg_Inst_ff_SDE_87_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_87_current_state_reg_U1 ( .A(RoundInput[87]), 
        .ZN(RoundReg_Inst_ff_SDE_87_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_87_next_state), .CK(clk), .Q(RoundInput[87]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .A(RoundOutput[88]), .B(
        plaintext[88]), .S(reset), .Z(RoundReg_Inst_ff_SDE_88_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_88_current_state_reg_U1 ( .A(RoundInput[88]), 
        .ZN(RoundReg_Inst_ff_SDE_88_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_88_next_state), .CK(clk), .Q(RoundInput[88]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .A(RoundOutput[89]), .B(
        plaintext[89]), .S(reset), .Z(RoundReg_Inst_ff_SDE_89_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_89_current_state_reg_U1 ( .A(RoundInput[89]), 
        .ZN(RoundReg_Inst_ff_SDE_89_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_89_next_state), .CK(clk), .Q(RoundInput[89]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .A(RoundOutput[90]), .B(
        plaintext[90]), .S(reset), .Z(RoundReg_Inst_ff_SDE_90_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_90_current_state_reg_U1 ( .A(RoundInput[90]), 
        .ZN(RoundReg_Inst_ff_SDE_90_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_90_next_state), .CK(clk), .Q(RoundInput[90]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .A(RoundOutput[91]), .B(
        plaintext[91]), .S(reset), .Z(RoundReg_Inst_ff_SDE_91_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_91_current_state_reg_U1 ( .A(RoundInput[91]), 
        .ZN(RoundReg_Inst_ff_SDE_91_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_91_next_state), .CK(clk), .Q(RoundInput[91]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .A(RoundOutput[92]), .B(
        plaintext[92]), .S(reset), .Z(RoundReg_Inst_ff_SDE_92_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_92_current_state_reg_U1 ( .A(RoundInput[92]), 
        .ZN(RoundReg_Inst_ff_SDE_92_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_92_next_state), .CK(clk), .Q(RoundInput[92]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .A(RoundOutput[93]), .B(
        plaintext[93]), .S(reset), .Z(RoundReg_Inst_ff_SDE_93_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_93_current_state_reg_U1 ( .A(RoundInput[93]), 
        .ZN(RoundReg_Inst_ff_SDE_93_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_93_next_state), .CK(clk), .Q(RoundInput[93]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .A(RoundOutput[94]), .B(
        plaintext[94]), .S(reset), .Z(RoundReg_Inst_ff_SDE_94_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_94_current_state_reg_U1 ( .A(RoundInput[94]), 
        .ZN(RoundReg_Inst_ff_SDE_94_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_94_next_state), .CK(clk), .Q(RoundInput[94]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .A(RoundOutput[95]), .B(
        plaintext[95]), .S(reset), .Z(RoundReg_Inst_ff_SDE_95_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_95_current_state_reg_U1 ( .A(RoundInput[95]), 
        .ZN(RoundReg_Inst_ff_SDE_95_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_95_next_state), .CK(clk), .Q(RoundInput[95]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .A(RoundOutput[96]), .B(
        plaintext[96]), .S(reset), .Z(RoundReg_Inst_ff_SDE_96_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_96_current_state_reg_U1 ( .A(RoundInput[96]), 
        .ZN(RoundReg_Inst_ff_SDE_96_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_96_next_state), .CK(clk), .Q(RoundInput[96]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .A(RoundOutput[97]), .B(
        plaintext[97]), .S(reset), .Z(RoundReg_Inst_ff_SDE_97_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_97_current_state_reg_U1 ( .A(RoundInput[97]), 
        .ZN(RoundReg_Inst_ff_SDE_97_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_97_next_state), .CK(clk), .Q(RoundInput[97]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .A(RoundOutput[98]), .B(
        plaintext[98]), .S(reset), .Z(RoundReg_Inst_ff_SDE_98_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_98_current_state_reg_U1 ( .A(RoundInput[98]), 
        .ZN(RoundReg_Inst_ff_SDE_98_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_98_next_state), .CK(clk), .Q(RoundInput[98]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .A(RoundOutput[99]), .B(
        plaintext[99]), .S(reset), .Z(RoundReg_Inst_ff_SDE_99_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_99_current_state_reg_U1 ( .A(RoundInput[99]), 
        .ZN(RoundReg_Inst_ff_SDE_99_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_99_next_state), .CK(clk), .Q(RoundInput[99]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .A(RoundOutput[100]), .B(
        plaintext[100]), .S(reset), .Z(RoundReg_Inst_ff_SDE_100_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_100_current_state_reg_U1 ( .A(RoundInput[100]), 
        .ZN(RoundReg_Inst_ff_SDE_100_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_100_next_state), .CK(clk), .Q(RoundInput[100]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .A(RoundOutput[101]), .B(
        plaintext[101]), .S(reset), .Z(RoundReg_Inst_ff_SDE_101_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_101_current_state_reg_U1 ( .A(RoundInput[101]), 
        .ZN(RoundReg_Inst_ff_SDE_101_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_101_next_state), .CK(clk), .Q(RoundInput[101]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .A(RoundOutput[102]), .B(
        plaintext[102]), .S(reset), .Z(RoundReg_Inst_ff_SDE_102_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_102_current_state_reg_U1 ( .A(RoundInput[102]), 
        .ZN(RoundReg_Inst_ff_SDE_102_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_102_next_state), .CK(clk), .Q(RoundInput[102]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .A(RoundOutput[103]), .B(
        plaintext[103]), .S(reset), .Z(RoundReg_Inst_ff_SDE_103_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_103_current_state_reg_U1 ( .A(RoundInput[103]), 
        .ZN(RoundReg_Inst_ff_SDE_103_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_103_next_state), .CK(clk), .Q(RoundInput[103]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .A(RoundOutput[104]), .B(
        plaintext[104]), .S(reset), .Z(RoundReg_Inst_ff_SDE_104_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_104_current_state_reg_U1 ( .A(RoundInput[104]), 
        .ZN(RoundReg_Inst_ff_SDE_104_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_104_next_state), .CK(clk), .Q(RoundInput[104]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .A(RoundOutput[105]), .B(
        plaintext[105]), .S(reset), .Z(RoundReg_Inst_ff_SDE_105_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_105_current_state_reg_U1 ( .A(RoundInput[105]), 
        .ZN(RoundReg_Inst_ff_SDE_105_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_105_next_state), .CK(clk), .Q(RoundInput[105]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .A(RoundOutput[106]), .B(
        plaintext[106]), .S(reset), .Z(RoundReg_Inst_ff_SDE_106_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_106_current_state_reg_U1 ( .A(RoundInput[106]), 
        .ZN(RoundReg_Inst_ff_SDE_106_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_106_next_state), .CK(clk), .Q(RoundInput[106]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .A(RoundOutput[107]), .B(
        plaintext[107]), .S(reset), .Z(RoundReg_Inst_ff_SDE_107_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_107_current_state_reg_U1 ( .A(RoundInput[107]), 
        .ZN(RoundReg_Inst_ff_SDE_107_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_107_next_state), .CK(clk), .Q(RoundInput[107]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .A(RoundOutput[108]), .B(
        plaintext[108]), .S(reset), .Z(RoundReg_Inst_ff_SDE_108_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_108_current_state_reg_U1 ( .A(RoundInput[108]), 
        .ZN(RoundReg_Inst_ff_SDE_108_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_108_next_state), .CK(clk), .Q(RoundInput[108]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .A(RoundOutput[109]), .B(
        plaintext[109]), .S(reset), .Z(RoundReg_Inst_ff_SDE_109_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_109_current_state_reg_U1 ( .A(RoundInput[109]), 
        .ZN(RoundReg_Inst_ff_SDE_109_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_109_next_state), .CK(clk), .Q(RoundInput[109]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .A(RoundOutput[110]), .B(
        plaintext[110]), .S(reset), .Z(RoundReg_Inst_ff_SDE_110_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_110_current_state_reg_U1 ( .A(RoundInput[110]), 
        .ZN(RoundReg_Inst_ff_SDE_110_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_110_next_state), .CK(clk), .Q(RoundInput[110]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .A(RoundOutput[111]), .B(
        plaintext[111]), .S(reset), .Z(RoundReg_Inst_ff_SDE_111_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_111_current_state_reg_U1 ( .A(RoundInput[111]), 
        .ZN(RoundReg_Inst_ff_SDE_111_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_111_next_state), .CK(clk), .Q(RoundInput[111]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .A(RoundOutput[112]), .B(
        plaintext[112]), .S(reset), .Z(RoundReg_Inst_ff_SDE_112_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_112_current_state_reg_U1 ( .A(RoundInput[112]), 
        .ZN(RoundReg_Inst_ff_SDE_112_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_112_next_state), .CK(clk), .Q(RoundInput[112]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .A(RoundOutput[113]), .B(
        plaintext[113]), .S(reset), .Z(RoundReg_Inst_ff_SDE_113_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_113_current_state_reg_U1 ( .A(RoundInput[113]), 
        .ZN(RoundReg_Inst_ff_SDE_113_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_113_next_state), .CK(clk), .Q(RoundInput[113]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .A(RoundOutput[114]), .B(
        plaintext[114]), .S(reset), .Z(RoundReg_Inst_ff_SDE_114_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_114_current_state_reg_U1 ( .A(RoundInput[114]), 
        .ZN(RoundReg_Inst_ff_SDE_114_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_114_next_state), .CK(clk), .Q(RoundInput[114]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .A(RoundOutput[115]), .B(
        plaintext[115]), .S(reset), .Z(RoundReg_Inst_ff_SDE_115_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_115_current_state_reg_U1 ( .A(RoundInput[115]), 
        .ZN(RoundReg_Inst_ff_SDE_115_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_115_next_state), .CK(clk), .Q(RoundInput[115]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .A(RoundOutput[116]), .B(
        plaintext[116]), .S(reset), .Z(RoundReg_Inst_ff_SDE_116_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_116_current_state_reg_U1 ( .A(RoundInput[116]), 
        .ZN(RoundReg_Inst_ff_SDE_116_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_116_next_state), .CK(clk), .Q(RoundInput[116]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .A(RoundOutput[117]), .B(
        plaintext[117]), .S(reset), .Z(RoundReg_Inst_ff_SDE_117_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_117_current_state_reg_U1 ( .A(RoundInput[117]), 
        .ZN(RoundReg_Inst_ff_SDE_117_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_117_next_state), .CK(clk), .Q(RoundInput[117]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .A(RoundOutput[118]), .B(
        plaintext[118]), .S(reset), .Z(RoundReg_Inst_ff_SDE_118_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_118_current_state_reg_U1 ( .A(RoundInput[118]), 
        .ZN(RoundReg_Inst_ff_SDE_118_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_118_next_state), .CK(clk), .Q(RoundInput[118]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .A(RoundOutput[119]), .B(
        plaintext[119]), .S(reset), .Z(RoundReg_Inst_ff_SDE_119_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_119_current_state_reg_U1 ( .A(RoundInput[119]), 
        .ZN(RoundReg_Inst_ff_SDE_119_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_119_next_state), .CK(clk), .Q(RoundInput[119]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .A(RoundOutput[120]), .B(
        plaintext[120]), .S(reset), .Z(RoundReg_Inst_ff_SDE_120_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_120_current_state_reg_U1 ( .A(RoundInput[120]), 
        .ZN(RoundReg_Inst_ff_SDE_120_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_120_next_state), .CK(clk), .Q(RoundInput[120]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .A(RoundOutput[121]), .B(
        plaintext[121]), .S(reset), .Z(RoundReg_Inst_ff_SDE_121_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_121_current_state_reg_U1 ( .A(RoundInput[121]), 
        .ZN(RoundReg_Inst_ff_SDE_121_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_121_next_state), .CK(clk), .Q(RoundInput[121]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .A(RoundOutput[122]), .B(
        plaintext[122]), .S(reset), .Z(RoundReg_Inst_ff_SDE_122_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_122_current_state_reg_U1 ( .A(RoundInput[122]), 
        .ZN(RoundReg_Inst_ff_SDE_122_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_122_next_state), .CK(clk), .Q(RoundInput[122]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .A(RoundOutput[123]), .B(
        plaintext[123]), .S(reset), .Z(RoundReg_Inst_ff_SDE_123_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_123_current_state_reg_U1 ( .A(RoundInput[123]), 
        .ZN(RoundReg_Inst_ff_SDE_123_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_123_next_state), .CK(clk), .Q(RoundInput[123]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .A(RoundOutput[124]), .B(
        plaintext[124]), .S(reset), .Z(RoundReg_Inst_ff_SDE_124_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_124_current_state_reg_U1 ( .A(RoundInput[124]), 
        .ZN(RoundReg_Inst_ff_SDE_124_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_124_next_state), .CK(clk), .Q(RoundInput[124]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .A(RoundOutput[125]), .B(
        plaintext[125]), .S(reset), .Z(RoundReg_Inst_ff_SDE_125_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_125_current_state_reg_U1 ( .A(RoundInput[125]), 
        .ZN(RoundReg_Inst_ff_SDE_125_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_125_next_state), .CK(clk), .Q(RoundInput[125]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .A(RoundOutput[126]), .B(
        plaintext[126]), .S(reset), .Z(RoundReg_Inst_ff_SDE_126_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_126_current_state_reg_U1 ( .A(RoundInput[126]), 
        .ZN(RoundReg_Inst_ff_SDE_126_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_126_next_state), .CK(clk), .Q(RoundInput[126]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .A(RoundOutput[127]), .B(
        plaintext[127]), .S(reset), .Z(RoundReg_Inst_ff_SDE_127_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_127_current_state_reg_U1 ( .A(RoundInput[127]), 
        .ZN(RoundReg_Inst_ff_SDE_127_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_127_next_state), .CK(clk), .Q(RoundInput[127]), 
        .QN() );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .A(ciphertext[7]), .B(
        ciphertext[4]), .Z(SubBytesIns_Inst_Sbox_0_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .A(ciphertext[7]), .B(
        ciphertext[2]), .Z(SubBytesIns_Inst_Sbox_0_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .A(ciphertext[7]), .B(
        ciphertext[1]), .Z(SubBytesIns_Inst_Sbox_0_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .A(ciphertext[4]), .B(
        ciphertext[2]), .Z(SubBytesIns_Inst_Sbox_0_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .A(ciphertext[3]), .B(
        ciphertext[1]), .Z(SubBytesIns_Inst_Sbox_0_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_0_T1), 
        .B(SubBytesIns_Inst_Sbox_0_T5), .Z(SubBytesIns_Inst_Sbox_0_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .A(ciphertext[6]), .B(
        ciphertext[5]), .Z(SubBytesIns_Inst_Sbox_0_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .A(ciphertext[0]), .B(
        SubBytesIns_Inst_Sbox_0_T6), .Z(SubBytesIns_Inst_Sbox_0_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .A(ciphertext[0]), .B(
        SubBytesIns_Inst_Sbox_0_T7), .Z(SubBytesIns_Inst_Sbox_0_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_0_T6), 
        .B(SubBytesIns_Inst_Sbox_0_T7), .Z(SubBytesIns_Inst_Sbox_0_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .A(ciphertext[6]), .B(
        ciphertext[2]), .Z(SubBytesIns_Inst_Sbox_0_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .A(ciphertext[5]), .B(
        ciphertext[2]), .Z(SubBytesIns_Inst_Sbox_0_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_0_T3), 
        .B(SubBytesIns_Inst_Sbox_0_T4), .Z(SubBytesIns_Inst_Sbox_0_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_0_T6), 
        .B(SubBytesIns_Inst_Sbox_0_T11), .Z(SubBytesIns_Inst_Sbox_0_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_0_T5), 
        .B(SubBytesIns_Inst_Sbox_0_T11), .Z(SubBytesIns_Inst_Sbox_0_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_0_T5), 
        .B(SubBytesIns_Inst_Sbox_0_T12), .Z(SubBytesIns_Inst_Sbox_0_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_0_T9), 
        .B(SubBytesIns_Inst_Sbox_0_T16), .Z(SubBytesIns_Inst_Sbox_0_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .A(ciphertext[4]), .B(
        ciphertext[0]), .Z(SubBytesIns_Inst_Sbox_0_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_0_T7), 
        .B(SubBytesIns_Inst_Sbox_0_T18), .Z(SubBytesIns_Inst_Sbox_0_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_0_T1), 
        .B(SubBytesIns_Inst_Sbox_0_T19), .Z(SubBytesIns_Inst_Sbox_0_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .A(ciphertext[1]), .B(
        ciphertext[0]), .Z(SubBytesIns_Inst_Sbox_0_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_0_T7), 
        .B(SubBytesIns_Inst_Sbox_0_T21), .Z(SubBytesIns_Inst_Sbox_0_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_0_T2), 
        .B(SubBytesIns_Inst_Sbox_0_T22), .Z(SubBytesIns_Inst_Sbox_0_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_0_T2), 
        .B(SubBytesIns_Inst_Sbox_0_T10), .Z(SubBytesIns_Inst_Sbox_0_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_0_T20), 
        .B(SubBytesIns_Inst_Sbox_0_T17), .Z(SubBytesIns_Inst_Sbox_0_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_0_T3), 
        .B(SubBytesIns_Inst_Sbox_0_T16), .Z(SubBytesIns_Inst_Sbox_0_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_0_T1), 
        .B(SubBytesIns_Inst_Sbox_0_T12), .Z(SubBytesIns_Inst_Sbox_0_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T13), 
        .A2(SubBytesIns_Inst_Sbox_0_T6), .ZN(SubBytesIns_Inst_Sbox_0_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T23), 
        .A2(SubBytesIns_Inst_Sbox_0_T8), .ZN(SubBytesIns_Inst_Sbox_0_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_0_T14), 
        .B(SubBytesIns_Inst_Sbox_0_M1), .Z(SubBytesIns_Inst_Sbox_0_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T19), 
        .A2(ciphertext[0]), .ZN(SubBytesIns_Inst_Sbox_0_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_0_M4), 
        .B(SubBytesIns_Inst_Sbox_0_M1), .Z(SubBytesIns_Inst_Sbox_0_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T3), 
        .A2(SubBytesIns_Inst_Sbox_0_T16), .ZN(SubBytesIns_Inst_Sbox_0_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T22), 
        .A2(SubBytesIns_Inst_Sbox_0_T9), .ZN(SubBytesIns_Inst_Sbox_0_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_0_T26), 
        .B(SubBytesIns_Inst_Sbox_0_M6), .Z(SubBytesIns_Inst_Sbox_0_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T20), 
        .A2(SubBytesIns_Inst_Sbox_0_T17), .ZN(SubBytesIns_Inst_Sbox_0_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_0_M9), 
        .B(SubBytesIns_Inst_Sbox_0_M6), .Z(SubBytesIns_Inst_Sbox_0_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T1), 
        .A2(SubBytesIns_Inst_Sbox_0_T15), .ZN(SubBytesIns_Inst_Sbox_0_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T4), 
        .A2(SubBytesIns_Inst_Sbox_0_T27), .ZN(SubBytesIns_Inst_Sbox_0_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_0_M12), 
        .B(SubBytesIns_Inst_Sbox_0_M11), .Z(SubBytesIns_Inst_Sbox_0_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T2), 
        .A2(SubBytesIns_Inst_Sbox_0_T10), .ZN(SubBytesIns_Inst_Sbox_0_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_0_M14), 
        .B(SubBytesIns_Inst_Sbox_0_M11), .Z(SubBytesIns_Inst_Sbox_0_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_0_M3), 
        .B(SubBytesIns_Inst_Sbox_0_M2), .Z(SubBytesIns_Inst_Sbox_0_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_0_M5), 
        .B(SubBytesIns_Inst_Sbox_0_T24), .Z(SubBytesIns_Inst_Sbox_0_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_0_M8), 
        .B(SubBytesIns_Inst_Sbox_0_M7), .Z(SubBytesIns_Inst_Sbox_0_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_0_M10), 
        .B(SubBytesIns_Inst_Sbox_0_M15), .Z(SubBytesIns_Inst_Sbox_0_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_0_M16), 
        .B(SubBytesIns_Inst_Sbox_0_M13), .Z(SubBytesIns_Inst_Sbox_0_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_0_M17), 
        .B(SubBytesIns_Inst_Sbox_0_M15), .Z(SubBytesIns_Inst_Sbox_0_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_0_M18), 
        .B(SubBytesIns_Inst_Sbox_0_M13), .Z(SubBytesIns_Inst_Sbox_0_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_0_M19), 
        .B(SubBytesIns_Inst_Sbox_0_T25), .Z(SubBytesIns_Inst_Sbox_0_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_0_M22), 
        .B(SubBytesIns_Inst_Sbox_0_M23), .Z(SubBytesIns_Inst_Sbox_0_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M22), .A2(SubBytesIns_Inst_Sbox_0_M20), .ZN(SubBytesIns_Inst_Sbox_0_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_0_M21), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_0_M20), 
        .B(SubBytesIns_Inst_Sbox_0_M21), .Z(SubBytesIns_Inst_Sbox_0_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_0_M23), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M28), .A2(SubBytesIns_Inst_Sbox_0_M27), .ZN(SubBytesIns_Inst_Sbox_0_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M26), .A2(SubBytesIns_Inst_Sbox_0_M24), .ZN(SubBytesIns_Inst_Sbox_0_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M20), .A2(SubBytesIns_Inst_Sbox_0_M23), .ZN(SubBytesIns_Inst_Sbox_0_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M27), .A2(SubBytesIns_Inst_Sbox_0_M31), .ZN(SubBytesIns_Inst_Sbox_0_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_0_M27), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M21), .A2(SubBytesIns_Inst_Sbox_0_M22), .ZN(SubBytesIns_Inst_Sbox_0_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M24), .A2(SubBytesIns_Inst_Sbox_0_M34), .ZN(SubBytesIns_Inst_Sbox_0_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_0_M24), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_0_M21), 
        .B(SubBytesIns_Inst_Sbox_0_M29), .Z(SubBytesIns_Inst_Sbox_0_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_0_M32), 
        .B(SubBytesIns_Inst_Sbox_0_M33), .Z(SubBytesIns_Inst_Sbox_0_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_0_M23), 
        .B(SubBytesIns_Inst_Sbox_0_M30), .Z(SubBytesIns_Inst_Sbox_0_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_0_M35), 
        .B(SubBytesIns_Inst_Sbox_0_M36), .Z(SubBytesIns_Inst_Sbox_0_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_0_M38), 
        .B(SubBytesIns_Inst_Sbox_0_M40), .Z(SubBytesIns_Inst_Sbox_0_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_0_M37), 
        .B(SubBytesIns_Inst_Sbox_0_M39), .Z(SubBytesIns_Inst_Sbox_0_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_0_M37), 
        .B(SubBytesIns_Inst_Sbox_0_M38), .Z(SubBytesIns_Inst_Sbox_0_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_0_M39), 
        .B(SubBytesIns_Inst_Sbox_0_M40), .Z(SubBytesIns_Inst_Sbox_0_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_0_M42), 
        .B(SubBytesIns_Inst_Sbox_0_M41), .Z(SubBytesIns_Inst_Sbox_0_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M44), .A2(SubBytesIns_Inst_Sbox_0_T6), .ZN(SubBytesIns_Inst_Sbox_0_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M40), .A2(SubBytesIns_Inst_Sbox_0_T8), .ZN(SubBytesIns_Inst_Sbox_0_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M39), .A2(ciphertext[0]), .ZN(SubBytesIns_Inst_Sbox_0_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M43), .A2(SubBytesIns_Inst_Sbox_0_T16), .ZN(SubBytesIns_Inst_Sbox_0_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M38), .A2(SubBytesIns_Inst_Sbox_0_T9), .ZN(SubBytesIns_Inst_Sbox_0_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M37), .A2(SubBytesIns_Inst_Sbox_0_T17), .ZN(SubBytesIns_Inst_Sbox_0_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M42), .A2(SubBytesIns_Inst_Sbox_0_T15), .ZN(SubBytesIns_Inst_Sbox_0_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M45), .A2(SubBytesIns_Inst_Sbox_0_T27), .ZN(SubBytesIns_Inst_Sbox_0_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M41), .A2(SubBytesIns_Inst_Sbox_0_T10), .ZN(SubBytesIns_Inst_Sbox_0_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M44), .A2(SubBytesIns_Inst_Sbox_0_T13), .ZN(SubBytesIns_Inst_Sbox_0_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M40), .A2(SubBytesIns_Inst_Sbox_0_T23), .ZN(SubBytesIns_Inst_Sbox_0_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M39), .A2(SubBytesIns_Inst_Sbox_0_T19), .ZN(SubBytesIns_Inst_Sbox_0_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M43), .A2(SubBytesIns_Inst_Sbox_0_T3), .ZN(SubBytesIns_Inst_Sbox_0_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M38), .A2(SubBytesIns_Inst_Sbox_0_T22), .ZN(SubBytesIns_Inst_Sbox_0_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M37), .A2(SubBytesIns_Inst_Sbox_0_T20), .ZN(SubBytesIns_Inst_Sbox_0_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M42), .A2(SubBytesIns_Inst_Sbox_0_T1), .ZN(SubBytesIns_Inst_Sbox_0_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M45), .A2(SubBytesIns_Inst_Sbox_0_T4), .ZN(SubBytesIns_Inst_Sbox_0_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M41), .A2(SubBytesIns_Inst_Sbox_0_T2), .ZN(SubBytesIns_Inst_Sbox_0_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_0_M61), 
        .B(SubBytesIns_Inst_Sbox_0_M62), .Z(SubBytesIns_Inst_Sbox_0_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_0_M50), 
        .B(SubBytesIns_Inst_Sbox_0_M56), .Z(SubBytesIns_Inst_Sbox_0_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_0_M46), 
        .B(SubBytesIns_Inst_Sbox_0_M48), .Z(SubBytesIns_Inst_Sbox_0_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_0_M47), 
        .B(SubBytesIns_Inst_Sbox_0_M55), .Z(SubBytesIns_Inst_Sbox_0_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_0_M54), 
        .B(SubBytesIns_Inst_Sbox_0_M58), .Z(SubBytesIns_Inst_Sbox_0_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_0_M49), 
        .B(SubBytesIns_Inst_Sbox_0_M61), .Z(SubBytesIns_Inst_Sbox_0_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_0_M62), 
        .B(SubBytesIns_Inst_Sbox_0_L5), .Z(SubBytesIns_Inst_Sbox_0_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_0_M46), 
        .B(SubBytesIns_Inst_Sbox_0_L3), .Z(SubBytesIns_Inst_Sbox_0_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_0_M51), 
        .B(SubBytesIns_Inst_Sbox_0_M59), .Z(SubBytesIns_Inst_Sbox_0_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_0_M52), 
        .B(SubBytesIns_Inst_Sbox_0_M53), .Z(SubBytesIns_Inst_Sbox_0_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_0_M53), 
        .B(SubBytesIns_Inst_Sbox_0_L4), .Z(SubBytesIns_Inst_Sbox_0_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_0_M60), 
        .B(SubBytesIns_Inst_Sbox_0_L2), .Z(SubBytesIns_Inst_Sbox_0_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_0_M48), 
        .B(SubBytesIns_Inst_Sbox_0_M51), .Z(SubBytesIns_Inst_Sbox_0_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_0_M50), 
        .B(SubBytesIns_Inst_Sbox_0_L0), .Z(SubBytesIns_Inst_Sbox_0_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_0_M52), 
        .B(SubBytesIns_Inst_Sbox_0_M61), .Z(SubBytesIns_Inst_Sbox_0_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_0_M55), 
        .B(SubBytesIns_Inst_Sbox_0_L1), .Z(SubBytesIns_Inst_Sbox_0_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_0_M56), 
        .B(SubBytesIns_Inst_Sbox_0_L0), .Z(SubBytesIns_Inst_Sbox_0_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_0_M57), 
        .B(SubBytesIns_Inst_Sbox_0_L1), .Z(SubBytesIns_Inst_Sbox_0_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_0_M58), 
        .B(SubBytesIns_Inst_Sbox_0_L8), .Z(SubBytesIns_Inst_Sbox_0_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_0_M63), 
        .B(SubBytesIns_Inst_Sbox_0_L4), .Z(SubBytesIns_Inst_Sbox_0_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_0_L0), 
        .B(SubBytesIns_Inst_Sbox_0_L1), .Z(SubBytesIns_Inst_Sbox_0_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_0_L1), 
        .B(SubBytesIns_Inst_Sbox_0_L7), .Z(SubBytesIns_Inst_Sbox_0_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_0_L3), 
        .B(SubBytesIns_Inst_Sbox_0_L12), .Z(SubBytesIns_Inst_Sbox_0_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_0_L18), 
        .B(SubBytesIns_Inst_Sbox_0_L2), .Z(SubBytesIns_Inst_Sbox_0_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_0_L15), 
        .B(SubBytesIns_Inst_Sbox_0_L9), .Z(SubBytesIns_Inst_Sbox_0_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L10), .Z(SubBytesIns_Inst_Sbox_0_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_0_L7), 
        .B(SubBytesIns_Inst_Sbox_0_L9), .Z(SubBytesIns_Inst_Sbox_0_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_0_L8), 
        .B(SubBytesIns_Inst_Sbox_0_L10), .Z(SubBytesIns_Inst_Sbox_0_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_0_L11), 
        .B(SubBytesIns_Inst_Sbox_0_L14), .Z(SubBytesIns_Inst_Sbox_0_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_0_L11), 
        .B(SubBytesIns_Inst_Sbox_0_L17), .Z(SubBytesIns_Inst_Sbox_0_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L24), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_0_L16), 
        .B(SubBytesIns_Inst_Sbox_0_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_0_L19), 
        .B(SubBytesIns_Inst_Sbox_0_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L21), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_0_L20), 
        .B(SubBytesIns_Inst_Sbox_0_L22), .Z(MixColumnsInput[99]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_0_L25), 
        .B(SubBytesIns_Inst_Sbox_0_L29), .Z(MixColumnsInput[98]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_0_L13), 
        .B(SubBytesIns_Inst_Sbox_0_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L23), .ZN(MixColumnsInput[96]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .A(ciphertext[15]), .B(
        ciphertext[12]), .Z(SubBytesIns_Inst_Sbox_1_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .A(ciphertext[15]), .B(
        ciphertext[10]), .Z(SubBytesIns_Inst_Sbox_1_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .A(ciphertext[15]), .B(
        ciphertext[9]), .Z(SubBytesIns_Inst_Sbox_1_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .A(ciphertext[12]), .B(
        ciphertext[10]), .Z(SubBytesIns_Inst_Sbox_1_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .A(ciphertext[11]), .B(
        ciphertext[9]), .Z(SubBytesIns_Inst_Sbox_1_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_1_T1), 
        .B(SubBytesIns_Inst_Sbox_1_T5), .Z(SubBytesIns_Inst_Sbox_1_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .A(ciphertext[14]), .B(
        ciphertext[13]), .Z(SubBytesIns_Inst_Sbox_1_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .A(ciphertext[8]), .B(
        SubBytesIns_Inst_Sbox_1_T6), .Z(SubBytesIns_Inst_Sbox_1_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .A(ciphertext[8]), .B(
        SubBytesIns_Inst_Sbox_1_T7), .Z(SubBytesIns_Inst_Sbox_1_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_1_T6), 
        .B(SubBytesIns_Inst_Sbox_1_T7), .Z(SubBytesIns_Inst_Sbox_1_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .A(ciphertext[14]), .B(
        ciphertext[10]), .Z(SubBytesIns_Inst_Sbox_1_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .A(ciphertext[13]), .B(
        ciphertext[10]), .Z(SubBytesIns_Inst_Sbox_1_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_1_T3), 
        .B(SubBytesIns_Inst_Sbox_1_T4), .Z(SubBytesIns_Inst_Sbox_1_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_1_T6), 
        .B(SubBytesIns_Inst_Sbox_1_T11), .Z(SubBytesIns_Inst_Sbox_1_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_1_T5), 
        .B(SubBytesIns_Inst_Sbox_1_T11), .Z(SubBytesIns_Inst_Sbox_1_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_1_T5), 
        .B(SubBytesIns_Inst_Sbox_1_T12), .Z(SubBytesIns_Inst_Sbox_1_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_1_T9), 
        .B(SubBytesIns_Inst_Sbox_1_T16), .Z(SubBytesIns_Inst_Sbox_1_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .A(ciphertext[12]), .B(
        ciphertext[8]), .Z(SubBytesIns_Inst_Sbox_1_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_1_T7), 
        .B(SubBytesIns_Inst_Sbox_1_T18), .Z(SubBytesIns_Inst_Sbox_1_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_1_T1), 
        .B(SubBytesIns_Inst_Sbox_1_T19), .Z(SubBytesIns_Inst_Sbox_1_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .A(ciphertext[9]), .B(
        ciphertext[8]), .Z(SubBytesIns_Inst_Sbox_1_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_1_T7), 
        .B(SubBytesIns_Inst_Sbox_1_T21), .Z(SubBytesIns_Inst_Sbox_1_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_1_T2), 
        .B(SubBytesIns_Inst_Sbox_1_T22), .Z(SubBytesIns_Inst_Sbox_1_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_1_T2), 
        .B(SubBytesIns_Inst_Sbox_1_T10), .Z(SubBytesIns_Inst_Sbox_1_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_1_T20), 
        .B(SubBytesIns_Inst_Sbox_1_T17), .Z(SubBytesIns_Inst_Sbox_1_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_1_T3), 
        .B(SubBytesIns_Inst_Sbox_1_T16), .Z(SubBytesIns_Inst_Sbox_1_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_1_T1), 
        .B(SubBytesIns_Inst_Sbox_1_T12), .Z(SubBytesIns_Inst_Sbox_1_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T13), 
        .A2(SubBytesIns_Inst_Sbox_1_T6), .ZN(SubBytesIns_Inst_Sbox_1_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T23), 
        .A2(SubBytesIns_Inst_Sbox_1_T8), .ZN(SubBytesIns_Inst_Sbox_1_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_1_T14), 
        .B(SubBytesIns_Inst_Sbox_1_M1), .Z(SubBytesIns_Inst_Sbox_1_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T19), 
        .A2(ciphertext[8]), .ZN(SubBytesIns_Inst_Sbox_1_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_1_M4), 
        .B(SubBytesIns_Inst_Sbox_1_M1), .Z(SubBytesIns_Inst_Sbox_1_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T3), 
        .A2(SubBytesIns_Inst_Sbox_1_T16), .ZN(SubBytesIns_Inst_Sbox_1_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T22), 
        .A2(SubBytesIns_Inst_Sbox_1_T9), .ZN(SubBytesIns_Inst_Sbox_1_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_1_T26), 
        .B(SubBytesIns_Inst_Sbox_1_M6), .Z(SubBytesIns_Inst_Sbox_1_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T20), 
        .A2(SubBytesIns_Inst_Sbox_1_T17), .ZN(SubBytesIns_Inst_Sbox_1_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_1_M9), 
        .B(SubBytesIns_Inst_Sbox_1_M6), .Z(SubBytesIns_Inst_Sbox_1_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T1), 
        .A2(SubBytesIns_Inst_Sbox_1_T15), .ZN(SubBytesIns_Inst_Sbox_1_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T4), 
        .A2(SubBytesIns_Inst_Sbox_1_T27), .ZN(SubBytesIns_Inst_Sbox_1_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_1_M12), 
        .B(SubBytesIns_Inst_Sbox_1_M11), .Z(SubBytesIns_Inst_Sbox_1_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T2), 
        .A2(SubBytesIns_Inst_Sbox_1_T10), .ZN(SubBytesIns_Inst_Sbox_1_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_1_M14), 
        .B(SubBytesIns_Inst_Sbox_1_M11), .Z(SubBytesIns_Inst_Sbox_1_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_1_M3), 
        .B(SubBytesIns_Inst_Sbox_1_M2), .Z(SubBytesIns_Inst_Sbox_1_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_1_M5), 
        .B(SubBytesIns_Inst_Sbox_1_T24), .Z(SubBytesIns_Inst_Sbox_1_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_1_M8), 
        .B(SubBytesIns_Inst_Sbox_1_M7), .Z(SubBytesIns_Inst_Sbox_1_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_1_M10), 
        .B(SubBytesIns_Inst_Sbox_1_M15), .Z(SubBytesIns_Inst_Sbox_1_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_1_M16), 
        .B(SubBytesIns_Inst_Sbox_1_M13), .Z(SubBytesIns_Inst_Sbox_1_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_1_M17), 
        .B(SubBytesIns_Inst_Sbox_1_M15), .Z(SubBytesIns_Inst_Sbox_1_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_1_M18), 
        .B(SubBytesIns_Inst_Sbox_1_M13), .Z(SubBytesIns_Inst_Sbox_1_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_1_M19), 
        .B(SubBytesIns_Inst_Sbox_1_T25), .Z(SubBytesIns_Inst_Sbox_1_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_1_M22), 
        .B(SubBytesIns_Inst_Sbox_1_M23), .Z(SubBytesIns_Inst_Sbox_1_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M22), .A2(SubBytesIns_Inst_Sbox_1_M20), .ZN(SubBytesIns_Inst_Sbox_1_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_1_M21), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_1_M20), 
        .B(SubBytesIns_Inst_Sbox_1_M21), .Z(SubBytesIns_Inst_Sbox_1_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_1_M23), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M28), .A2(SubBytesIns_Inst_Sbox_1_M27), .ZN(SubBytesIns_Inst_Sbox_1_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M26), .A2(SubBytesIns_Inst_Sbox_1_M24), .ZN(SubBytesIns_Inst_Sbox_1_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M20), .A2(SubBytesIns_Inst_Sbox_1_M23), .ZN(SubBytesIns_Inst_Sbox_1_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M27), .A2(SubBytesIns_Inst_Sbox_1_M31), .ZN(SubBytesIns_Inst_Sbox_1_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_1_M27), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M21), .A2(SubBytesIns_Inst_Sbox_1_M22), .ZN(SubBytesIns_Inst_Sbox_1_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M24), .A2(SubBytesIns_Inst_Sbox_1_M34), .ZN(SubBytesIns_Inst_Sbox_1_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_1_M24), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_1_M21), 
        .B(SubBytesIns_Inst_Sbox_1_M29), .Z(SubBytesIns_Inst_Sbox_1_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_1_M32), 
        .B(SubBytesIns_Inst_Sbox_1_M33), .Z(SubBytesIns_Inst_Sbox_1_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_1_M23), 
        .B(SubBytesIns_Inst_Sbox_1_M30), .Z(SubBytesIns_Inst_Sbox_1_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_1_M35), 
        .B(SubBytesIns_Inst_Sbox_1_M36), .Z(SubBytesIns_Inst_Sbox_1_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_1_M38), 
        .B(SubBytesIns_Inst_Sbox_1_M40), .Z(SubBytesIns_Inst_Sbox_1_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_1_M37), 
        .B(SubBytesIns_Inst_Sbox_1_M39), .Z(SubBytesIns_Inst_Sbox_1_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_1_M37), 
        .B(SubBytesIns_Inst_Sbox_1_M38), .Z(SubBytesIns_Inst_Sbox_1_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_1_M39), 
        .B(SubBytesIns_Inst_Sbox_1_M40), .Z(SubBytesIns_Inst_Sbox_1_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_1_M42), 
        .B(SubBytesIns_Inst_Sbox_1_M41), .Z(SubBytesIns_Inst_Sbox_1_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M44), .A2(SubBytesIns_Inst_Sbox_1_T6), .ZN(SubBytesIns_Inst_Sbox_1_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M40), .A2(SubBytesIns_Inst_Sbox_1_T8), .ZN(SubBytesIns_Inst_Sbox_1_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M39), .A2(ciphertext[8]), .ZN(SubBytesIns_Inst_Sbox_1_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M43), .A2(SubBytesIns_Inst_Sbox_1_T16), .ZN(SubBytesIns_Inst_Sbox_1_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M38), .A2(SubBytesIns_Inst_Sbox_1_T9), .ZN(SubBytesIns_Inst_Sbox_1_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M37), .A2(SubBytesIns_Inst_Sbox_1_T17), .ZN(SubBytesIns_Inst_Sbox_1_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M42), .A2(SubBytesIns_Inst_Sbox_1_T15), .ZN(SubBytesIns_Inst_Sbox_1_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M45), .A2(SubBytesIns_Inst_Sbox_1_T27), .ZN(SubBytesIns_Inst_Sbox_1_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M41), .A2(SubBytesIns_Inst_Sbox_1_T10), .ZN(SubBytesIns_Inst_Sbox_1_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M44), .A2(SubBytesIns_Inst_Sbox_1_T13), .ZN(SubBytesIns_Inst_Sbox_1_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M40), .A2(SubBytesIns_Inst_Sbox_1_T23), .ZN(SubBytesIns_Inst_Sbox_1_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M39), .A2(SubBytesIns_Inst_Sbox_1_T19), .ZN(SubBytesIns_Inst_Sbox_1_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M43), .A2(SubBytesIns_Inst_Sbox_1_T3), .ZN(SubBytesIns_Inst_Sbox_1_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M38), .A2(SubBytesIns_Inst_Sbox_1_T22), .ZN(SubBytesIns_Inst_Sbox_1_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M37), .A2(SubBytesIns_Inst_Sbox_1_T20), .ZN(SubBytesIns_Inst_Sbox_1_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M42), .A2(SubBytesIns_Inst_Sbox_1_T1), .ZN(SubBytesIns_Inst_Sbox_1_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M45), .A2(SubBytesIns_Inst_Sbox_1_T4), .ZN(SubBytesIns_Inst_Sbox_1_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M41), .A2(SubBytesIns_Inst_Sbox_1_T2), .ZN(SubBytesIns_Inst_Sbox_1_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_1_M61), 
        .B(SubBytesIns_Inst_Sbox_1_M62), .Z(SubBytesIns_Inst_Sbox_1_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_1_M50), 
        .B(SubBytesIns_Inst_Sbox_1_M56), .Z(SubBytesIns_Inst_Sbox_1_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_1_M46), 
        .B(SubBytesIns_Inst_Sbox_1_M48), .Z(SubBytesIns_Inst_Sbox_1_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_1_M47), 
        .B(SubBytesIns_Inst_Sbox_1_M55), .Z(SubBytesIns_Inst_Sbox_1_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_1_M54), 
        .B(SubBytesIns_Inst_Sbox_1_M58), .Z(SubBytesIns_Inst_Sbox_1_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_1_M49), 
        .B(SubBytesIns_Inst_Sbox_1_M61), .Z(SubBytesIns_Inst_Sbox_1_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_1_M62), 
        .B(SubBytesIns_Inst_Sbox_1_L5), .Z(SubBytesIns_Inst_Sbox_1_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_1_M46), 
        .B(SubBytesIns_Inst_Sbox_1_L3), .Z(SubBytesIns_Inst_Sbox_1_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_1_M51), 
        .B(SubBytesIns_Inst_Sbox_1_M59), .Z(SubBytesIns_Inst_Sbox_1_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_1_M52), 
        .B(SubBytesIns_Inst_Sbox_1_M53), .Z(SubBytesIns_Inst_Sbox_1_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_1_M53), 
        .B(SubBytesIns_Inst_Sbox_1_L4), .Z(SubBytesIns_Inst_Sbox_1_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_1_M60), 
        .B(SubBytesIns_Inst_Sbox_1_L2), .Z(SubBytesIns_Inst_Sbox_1_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_1_M48), 
        .B(SubBytesIns_Inst_Sbox_1_M51), .Z(SubBytesIns_Inst_Sbox_1_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_1_M50), 
        .B(SubBytesIns_Inst_Sbox_1_L0), .Z(SubBytesIns_Inst_Sbox_1_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_1_M52), 
        .B(SubBytesIns_Inst_Sbox_1_M61), .Z(SubBytesIns_Inst_Sbox_1_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_1_M55), 
        .B(SubBytesIns_Inst_Sbox_1_L1), .Z(SubBytesIns_Inst_Sbox_1_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_1_M56), 
        .B(SubBytesIns_Inst_Sbox_1_L0), .Z(SubBytesIns_Inst_Sbox_1_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_1_M57), 
        .B(SubBytesIns_Inst_Sbox_1_L1), .Z(SubBytesIns_Inst_Sbox_1_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_1_M58), 
        .B(SubBytesIns_Inst_Sbox_1_L8), .Z(SubBytesIns_Inst_Sbox_1_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_1_M63), 
        .B(SubBytesIns_Inst_Sbox_1_L4), .Z(SubBytesIns_Inst_Sbox_1_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_1_L0), 
        .B(SubBytesIns_Inst_Sbox_1_L1), .Z(SubBytesIns_Inst_Sbox_1_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_1_L1), 
        .B(SubBytesIns_Inst_Sbox_1_L7), .Z(SubBytesIns_Inst_Sbox_1_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_1_L3), 
        .B(SubBytesIns_Inst_Sbox_1_L12), .Z(SubBytesIns_Inst_Sbox_1_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_1_L18), 
        .B(SubBytesIns_Inst_Sbox_1_L2), .Z(SubBytesIns_Inst_Sbox_1_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_1_L15), 
        .B(SubBytesIns_Inst_Sbox_1_L9), .Z(SubBytesIns_Inst_Sbox_1_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L10), .Z(SubBytesIns_Inst_Sbox_1_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_1_L7), 
        .B(SubBytesIns_Inst_Sbox_1_L9), .Z(SubBytesIns_Inst_Sbox_1_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_1_L8), 
        .B(SubBytesIns_Inst_Sbox_1_L10), .Z(SubBytesIns_Inst_Sbox_1_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_1_L11), 
        .B(SubBytesIns_Inst_Sbox_1_L14), .Z(SubBytesIns_Inst_Sbox_1_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_1_L11), 
        .B(SubBytesIns_Inst_Sbox_1_L17), .Z(SubBytesIns_Inst_Sbox_1_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L24), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_1_L16), 
        .B(SubBytesIns_Inst_Sbox_1_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_1_L19), 
        .B(SubBytesIns_Inst_Sbox_1_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L21), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_1_L20), 
        .B(SubBytesIns_Inst_Sbox_1_L22), .Z(MixColumnsInput[75]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_1_L25), 
        .B(SubBytesIns_Inst_Sbox_1_L29), .Z(MixColumnsInput[74]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_1_L13), 
        .B(SubBytesIns_Inst_Sbox_1_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L23), .ZN(MixColumnsInput[72]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .A(ciphertext[23]), .B(
        ciphertext[20]), .Z(SubBytesIns_Inst_Sbox_2_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .A(ciphertext[23]), .B(
        ciphertext[18]), .Z(SubBytesIns_Inst_Sbox_2_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .A(ciphertext[23]), .B(
        ciphertext[17]), .Z(SubBytesIns_Inst_Sbox_2_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .A(ciphertext[20]), .B(
        ciphertext[18]), .Z(SubBytesIns_Inst_Sbox_2_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .A(ciphertext[19]), .B(
        ciphertext[17]), .Z(SubBytesIns_Inst_Sbox_2_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_2_T1), 
        .B(SubBytesIns_Inst_Sbox_2_T5), .Z(SubBytesIns_Inst_Sbox_2_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .A(ciphertext[22]), .B(
        ciphertext[21]), .Z(SubBytesIns_Inst_Sbox_2_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .A(ciphertext[16]), .B(
        SubBytesIns_Inst_Sbox_2_T6), .Z(SubBytesIns_Inst_Sbox_2_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .A(ciphertext[16]), .B(
        SubBytesIns_Inst_Sbox_2_T7), .Z(SubBytesIns_Inst_Sbox_2_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_2_T6), 
        .B(SubBytesIns_Inst_Sbox_2_T7), .Z(SubBytesIns_Inst_Sbox_2_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .A(ciphertext[22]), .B(
        ciphertext[18]), .Z(SubBytesIns_Inst_Sbox_2_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .A(ciphertext[21]), .B(
        ciphertext[18]), .Z(SubBytesIns_Inst_Sbox_2_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_2_T3), 
        .B(SubBytesIns_Inst_Sbox_2_T4), .Z(SubBytesIns_Inst_Sbox_2_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_2_T6), 
        .B(SubBytesIns_Inst_Sbox_2_T11), .Z(SubBytesIns_Inst_Sbox_2_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_2_T5), 
        .B(SubBytesIns_Inst_Sbox_2_T11), .Z(SubBytesIns_Inst_Sbox_2_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_2_T5), 
        .B(SubBytesIns_Inst_Sbox_2_T12), .Z(SubBytesIns_Inst_Sbox_2_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_2_T9), 
        .B(SubBytesIns_Inst_Sbox_2_T16), .Z(SubBytesIns_Inst_Sbox_2_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .A(ciphertext[20]), .B(
        ciphertext[16]), .Z(SubBytesIns_Inst_Sbox_2_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_2_T7), 
        .B(SubBytesIns_Inst_Sbox_2_T18), .Z(SubBytesIns_Inst_Sbox_2_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_2_T1), 
        .B(SubBytesIns_Inst_Sbox_2_T19), .Z(SubBytesIns_Inst_Sbox_2_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .A(ciphertext[17]), .B(
        ciphertext[16]), .Z(SubBytesIns_Inst_Sbox_2_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_2_T7), 
        .B(SubBytesIns_Inst_Sbox_2_T21), .Z(SubBytesIns_Inst_Sbox_2_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_2_T2), 
        .B(SubBytesIns_Inst_Sbox_2_T22), .Z(SubBytesIns_Inst_Sbox_2_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_2_T2), 
        .B(SubBytesIns_Inst_Sbox_2_T10), .Z(SubBytesIns_Inst_Sbox_2_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_2_T20), 
        .B(SubBytesIns_Inst_Sbox_2_T17), .Z(SubBytesIns_Inst_Sbox_2_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_2_T3), 
        .B(SubBytesIns_Inst_Sbox_2_T16), .Z(SubBytesIns_Inst_Sbox_2_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_2_T1), 
        .B(SubBytesIns_Inst_Sbox_2_T12), .Z(SubBytesIns_Inst_Sbox_2_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T13), 
        .A2(SubBytesIns_Inst_Sbox_2_T6), .ZN(SubBytesIns_Inst_Sbox_2_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T23), 
        .A2(SubBytesIns_Inst_Sbox_2_T8), .ZN(SubBytesIns_Inst_Sbox_2_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_2_T14), 
        .B(SubBytesIns_Inst_Sbox_2_M1), .Z(SubBytesIns_Inst_Sbox_2_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T19), 
        .A2(ciphertext[16]), .ZN(SubBytesIns_Inst_Sbox_2_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_2_M4), 
        .B(SubBytesIns_Inst_Sbox_2_M1), .Z(SubBytesIns_Inst_Sbox_2_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T3), 
        .A2(SubBytesIns_Inst_Sbox_2_T16), .ZN(SubBytesIns_Inst_Sbox_2_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T22), 
        .A2(SubBytesIns_Inst_Sbox_2_T9), .ZN(SubBytesIns_Inst_Sbox_2_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_2_T26), 
        .B(SubBytesIns_Inst_Sbox_2_M6), .Z(SubBytesIns_Inst_Sbox_2_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T20), 
        .A2(SubBytesIns_Inst_Sbox_2_T17), .ZN(SubBytesIns_Inst_Sbox_2_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_2_M9), 
        .B(SubBytesIns_Inst_Sbox_2_M6), .Z(SubBytesIns_Inst_Sbox_2_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T1), 
        .A2(SubBytesIns_Inst_Sbox_2_T15), .ZN(SubBytesIns_Inst_Sbox_2_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T4), 
        .A2(SubBytesIns_Inst_Sbox_2_T27), .ZN(SubBytesIns_Inst_Sbox_2_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_2_M12), 
        .B(SubBytesIns_Inst_Sbox_2_M11), .Z(SubBytesIns_Inst_Sbox_2_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T2), 
        .A2(SubBytesIns_Inst_Sbox_2_T10), .ZN(SubBytesIns_Inst_Sbox_2_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_2_M14), 
        .B(SubBytesIns_Inst_Sbox_2_M11), .Z(SubBytesIns_Inst_Sbox_2_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_2_M3), 
        .B(SubBytesIns_Inst_Sbox_2_M2), .Z(SubBytesIns_Inst_Sbox_2_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_2_M5), 
        .B(SubBytesIns_Inst_Sbox_2_T24), .Z(SubBytesIns_Inst_Sbox_2_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_2_M8), 
        .B(SubBytesIns_Inst_Sbox_2_M7), .Z(SubBytesIns_Inst_Sbox_2_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_2_M10), 
        .B(SubBytesIns_Inst_Sbox_2_M15), .Z(SubBytesIns_Inst_Sbox_2_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_2_M16), 
        .B(SubBytesIns_Inst_Sbox_2_M13), .Z(SubBytesIns_Inst_Sbox_2_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_2_M17), 
        .B(SubBytesIns_Inst_Sbox_2_M15), .Z(SubBytesIns_Inst_Sbox_2_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_2_M18), 
        .B(SubBytesIns_Inst_Sbox_2_M13), .Z(SubBytesIns_Inst_Sbox_2_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_2_M19), 
        .B(SubBytesIns_Inst_Sbox_2_T25), .Z(SubBytesIns_Inst_Sbox_2_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_2_M22), 
        .B(SubBytesIns_Inst_Sbox_2_M23), .Z(SubBytesIns_Inst_Sbox_2_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M22), .A2(SubBytesIns_Inst_Sbox_2_M20), .ZN(SubBytesIns_Inst_Sbox_2_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_2_M21), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_2_M20), 
        .B(SubBytesIns_Inst_Sbox_2_M21), .Z(SubBytesIns_Inst_Sbox_2_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_2_M23), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M28), .A2(SubBytesIns_Inst_Sbox_2_M27), .ZN(SubBytesIns_Inst_Sbox_2_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M26), .A2(SubBytesIns_Inst_Sbox_2_M24), .ZN(SubBytesIns_Inst_Sbox_2_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M20), .A2(SubBytesIns_Inst_Sbox_2_M23), .ZN(SubBytesIns_Inst_Sbox_2_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M27), .A2(SubBytesIns_Inst_Sbox_2_M31), .ZN(SubBytesIns_Inst_Sbox_2_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_2_M27), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M21), .A2(SubBytesIns_Inst_Sbox_2_M22), .ZN(SubBytesIns_Inst_Sbox_2_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M24), .A2(SubBytesIns_Inst_Sbox_2_M34), .ZN(SubBytesIns_Inst_Sbox_2_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_2_M24), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_2_M21), 
        .B(SubBytesIns_Inst_Sbox_2_M29), .Z(SubBytesIns_Inst_Sbox_2_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_2_M32), 
        .B(SubBytesIns_Inst_Sbox_2_M33), .Z(SubBytesIns_Inst_Sbox_2_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_2_M23), 
        .B(SubBytesIns_Inst_Sbox_2_M30), .Z(SubBytesIns_Inst_Sbox_2_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_2_M35), 
        .B(SubBytesIns_Inst_Sbox_2_M36), .Z(SubBytesIns_Inst_Sbox_2_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_2_M38), 
        .B(SubBytesIns_Inst_Sbox_2_M40), .Z(SubBytesIns_Inst_Sbox_2_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_2_M37), 
        .B(SubBytesIns_Inst_Sbox_2_M39), .Z(SubBytesIns_Inst_Sbox_2_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_2_M37), 
        .B(SubBytesIns_Inst_Sbox_2_M38), .Z(SubBytesIns_Inst_Sbox_2_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_2_M39), 
        .B(SubBytesIns_Inst_Sbox_2_M40), .Z(SubBytesIns_Inst_Sbox_2_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_2_M42), 
        .B(SubBytesIns_Inst_Sbox_2_M41), .Z(SubBytesIns_Inst_Sbox_2_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M44), .A2(SubBytesIns_Inst_Sbox_2_T6), .ZN(SubBytesIns_Inst_Sbox_2_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M40), .A2(SubBytesIns_Inst_Sbox_2_T8), .ZN(SubBytesIns_Inst_Sbox_2_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M39), .A2(ciphertext[16]), .ZN(SubBytesIns_Inst_Sbox_2_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M43), .A2(SubBytesIns_Inst_Sbox_2_T16), .ZN(SubBytesIns_Inst_Sbox_2_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M38), .A2(SubBytesIns_Inst_Sbox_2_T9), .ZN(SubBytesIns_Inst_Sbox_2_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M37), .A2(SubBytesIns_Inst_Sbox_2_T17), .ZN(SubBytesIns_Inst_Sbox_2_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M42), .A2(SubBytesIns_Inst_Sbox_2_T15), .ZN(SubBytesIns_Inst_Sbox_2_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M45), .A2(SubBytesIns_Inst_Sbox_2_T27), .ZN(SubBytesIns_Inst_Sbox_2_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M41), .A2(SubBytesIns_Inst_Sbox_2_T10), .ZN(SubBytesIns_Inst_Sbox_2_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M44), .A2(SubBytesIns_Inst_Sbox_2_T13), .ZN(SubBytesIns_Inst_Sbox_2_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M40), .A2(SubBytesIns_Inst_Sbox_2_T23), .ZN(SubBytesIns_Inst_Sbox_2_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M39), .A2(SubBytesIns_Inst_Sbox_2_T19), .ZN(SubBytesIns_Inst_Sbox_2_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M43), .A2(SubBytesIns_Inst_Sbox_2_T3), .ZN(SubBytesIns_Inst_Sbox_2_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M38), .A2(SubBytesIns_Inst_Sbox_2_T22), .ZN(SubBytesIns_Inst_Sbox_2_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M37), .A2(SubBytesIns_Inst_Sbox_2_T20), .ZN(SubBytesIns_Inst_Sbox_2_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M42), .A2(SubBytesIns_Inst_Sbox_2_T1), .ZN(SubBytesIns_Inst_Sbox_2_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M45), .A2(SubBytesIns_Inst_Sbox_2_T4), .ZN(SubBytesIns_Inst_Sbox_2_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M41), .A2(SubBytesIns_Inst_Sbox_2_T2), .ZN(SubBytesIns_Inst_Sbox_2_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_2_M61), 
        .B(SubBytesIns_Inst_Sbox_2_M62), .Z(SubBytesIns_Inst_Sbox_2_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_2_M50), 
        .B(SubBytesIns_Inst_Sbox_2_M56), .Z(SubBytesIns_Inst_Sbox_2_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_2_M46), 
        .B(SubBytesIns_Inst_Sbox_2_M48), .Z(SubBytesIns_Inst_Sbox_2_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_2_M47), 
        .B(SubBytesIns_Inst_Sbox_2_M55), .Z(SubBytesIns_Inst_Sbox_2_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_2_M54), 
        .B(SubBytesIns_Inst_Sbox_2_M58), .Z(SubBytesIns_Inst_Sbox_2_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_2_M49), 
        .B(SubBytesIns_Inst_Sbox_2_M61), .Z(SubBytesIns_Inst_Sbox_2_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_2_M62), 
        .B(SubBytesIns_Inst_Sbox_2_L5), .Z(SubBytesIns_Inst_Sbox_2_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_2_M46), 
        .B(SubBytesIns_Inst_Sbox_2_L3), .Z(SubBytesIns_Inst_Sbox_2_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_2_M51), 
        .B(SubBytesIns_Inst_Sbox_2_M59), .Z(SubBytesIns_Inst_Sbox_2_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_2_M52), 
        .B(SubBytesIns_Inst_Sbox_2_M53), .Z(SubBytesIns_Inst_Sbox_2_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_2_M53), 
        .B(SubBytesIns_Inst_Sbox_2_L4), .Z(SubBytesIns_Inst_Sbox_2_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_2_M60), 
        .B(SubBytesIns_Inst_Sbox_2_L2), .Z(SubBytesIns_Inst_Sbox_2_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_2_M48), 
        .B(SubBytesIns_Inst_Sbox_2_M51), .Z(SubBytesIns_Inst_Sbox_2_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_2_M50), 
        .B(SubBytesIns_Inst_Sbox_2_L0), .Z(SubBytesIns_Inst_Sbox_2_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_2_M52), 
        .B(SubBytesIns_Inst_Sbox_2_M61), .Z(SubBytesIns_Inst_Sbox_2_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_2_M55), 
        .B(SubBytesIns_Inst_Sbox_2_L1), .Z(SubBytesIns_Inst_Sbox_2_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_2_M56), 
        .B(SubBytesIns_Inst_Sbox_2_L0), .Z(SubBytesIns_Inst_Sbox_2_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_2_M57), 
        .B(SubBytesIns_Inst_Sbox_2_L1), .Z(SubBytesIns_Inst_Sbox_2_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_2_M58), 
        .B(SubBytesIns_Inst_Sbox_2_L8), .Z(SubBytesIns_Inst_Sbox_2_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_2_M63), 
        .B(SubBytesIns_Inst_Sbox_2_L4), .Z(SubBytesIns_Inst_Sbox_2_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_2_L0), 
        .B(SubBytesIns_Inst_Sbox_2_L1), .Z(SubBytesIns_Inst_Sbox_2_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_2_L1), 
        .B(SubBytesIns_Inst_Sbox_2_L7), .Z(SubBytesIns_Inst_Sbox_2_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_2_L3), 
        .B(SubBytesIns_Inst_Sbox_2_L12), .Z(SubBytesIns_Inst_Sbox_2_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_2_L18), 
        .B(SubBytesIns_Inst_Sbox_2_L2), .Z(SubBytesIns_Inst_Sbox_2_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_2_L15), 
        .B(SubBytesIns_Inst_Sbox_2_L9), .Z(SubBytesIns_Inst_Sbox_2_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L10), .Z(SubBytesIns_Inst_Sbox_2_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_2_L7), 
        .B(SubBytesIns_Inst_Sbox_2_L9), .Z(SubBytesIns_Inst_Sbox_2_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_2_L8), 
        .B(SubBytesIns_Inst_Sbox_2_L10), .Z(SubBytesIns_Inst_Sbox_2_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_2_L11), 
        .B(SubBytesIns_Inst_Sbox_2_L14), .Z(SubBytesIns_Inst_Sbox_2_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_2_L11), 
        .B(SubBytesIns_Inst_Sbox_2_L17), .Z(SubBytesIns_Inst_Sbox_2_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L24), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_2_L16), 
        .B(SubBytesIns_Inst_Sbox_2_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_2_L19), 
        .B(SubBytesIns_Inst_Sbox_2_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L21), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_2_L20), 
        .B(SubBytesIns_Inst_Sbox_2_L22), .Z(MixColumnsInput[51]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_2_L25), 
        .B(SubBytesIns_Inst_Sbox_2_L29), .Z(MixColumnsInput[50]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_2_L13), 
        .B(SubBytesIns_Inst_Sbox_2_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L23), .ZN(MixColumnsInput[48]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .A(ciphertext[31]), .B(
        ciphertext[28]), .Z(SubBytesIns_Inst_Sbox_3_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .A(ciphertext[31]), .B(
        ciphertext[26]), .Z(SubBytesIns_Inst_Sbox_3_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .A(ciphertext[31]), .B(
        ciphertext[25]), .Z(SubBytesIns_Inst_Sbox_3_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .A(ciphertext[28]), .B(
        ciphertext[26]), .Z(SubBytesIns_Inst_Sbox_3_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .A(ciphertext[27]), .B(
        ciphertext[25]), .Z(SubBytesIns_Inst_Sbox_3_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_3_T1), 
        .B(SubBytesIns_Inst_Sbox_3_T5), .Z(SubBytesIns_Inst_Sbox_3_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .A(ciphertext[30]), .B(
        ciphertext[29]), .Z(SubBytesIns_Inst_Sbox_3_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .A(ciphertext[24]), .B(
        SubBytesIns_Inst_Sbox_3_T6), .Z(SubBytesIns_Inst_Sbox_3_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .A(ciphertext[24]), .B(
        SubBytesIns_Inst_Sbox_3_T7), .Z(SubBytesIns_Inst_Sbox_3_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_3_T6), 
        .B(SubBytesIns_Inst_Sbox_3_T7), .Z(SubBytesIns_Inst_Sbox_3_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .A(ciphertext[30]), .B(
        ciphertext[26]), .Z(SubBytesIns_Inst_Sbox_3_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .A(ciphertext[29]), .B(
        ciphertext[26]), .Z(SubBytesIns_Inst_Sbox_3_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_3_T3), 
        .B(SubBytesIns_Inst_Sbox_3_T4), .Z(SubBytesIns_Inst_Sbox_3_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_3_T6), 
        .B(SubBytesIns_Inst_Sbox_3_T11), .Z(SubBytesIns_Inst_Sbox_3_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_3_T5), 
        .B(SubBytesIns_Inst_Sbox_3_T11), .Z(SubBytesIns_Inst_Sbox_3_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_3_T5), 
        .B(SubBytesIns_Inst_Sbox_3_T12), .Z(SubBytesIns_Inst_Sbox_3_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_3_T9), 
        .B(SubBytesIns_Inst_Sbox_3_T16), .Z(SubBytesIns_Inst_Sbox_3_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .A(ciphertext[28]), .B(
        ciphertext[24]), .Z(SubBytesIns_Inst_Sbox_3_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_3_T7), 
        .B(SubBytesIns_Inst_Sbox_3_T18), .Z(SubBytesIns_Inst_Sbox_3_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_3_T1), 
        .B(SubBytesIns_Inst_Sbox_3_T19), .Z(SubBytesIns_Inst_Sbox_3_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .A(ciphertext[25]), .B(
        ciphertext[24]), .Z(SubBytesIns_Inst_Sbox_3_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_3_T7), 
        .B(SubBytesIns_Inst_Sbox_3_T21), .Z(SubBytesIns_Inst_Sbox_3_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_3_T2), 
        .B(SubBytesIns_Inst_Sbox_3_T22), .Z(SubBytesIns_Inst_Sbox_3_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_3_T2), 
        .B(SubBytesIns_Inst_Sbox_3_T10), .Z(SubBytesIns_Inst_Sbox_3_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_3_T20), 
        .B(SubBytesIns_Inst_Sbox_3_T17), .Z(SubBytesIns_Inst_Sbox_3_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_3_T3), 
        .B(SubBytesIns_Inst_Sbox_3_T16), .Z(SubBytesIns_Inst_Sbox_3_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_3_T1), 
        .B(SubBytesIns_Inst_Sbox_3_T12), .Z(SubBytesIns_Inst_Sbox_3_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T13), 
        .A2(SubBytesIns_Inst_Sbox_3_T6), .ZN(SubBytesIns_Inst_Sbox_3_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T23), 
        .A2(SubBytesIns_Inst_Sbox_3_T8), .ZN(SubBytesIns_Inst_Sbox_3_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_3_T14), 
        .B(SubBytesIns_Inst_Sbox_3_M1), .Z(SubBytesIns_Inst_Sbox_3_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T19), 
        .A2(ciphertext[24]), .ZN(SubBytesIns_Inst_Sbox_3_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_3_M4), 
        .B(SubBytesIns_Inst_Sbox_3_M1), .Z(SubBytesIns_Inst_Sbox_3_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T3), 
        .A2(SubBytesIns_Inst_Sbox_3_T16), .ZN(SubBytesIns_Inst_Sbox_3_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T22), 
        .A2(SubBytesIns_Inst_Sbox_3_T9), .ZN(SubBytesIns_Inst_Sbox_3_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_3_T26), 
        .B(SubBytesIns_Inst_Sbox_3_M6), .Z(SubBytesIns_Inst_Sbox_3_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T20), 
        .A2(SubBytesIns_Inst_Sbox_3_T17), .ZN(SubBytesIns_Inst_Sbox_3_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_3_M9), 
        .B(SubBytesIns_Inst_Sbox_3_M6), .Z(SubBytesIns_Inst_Sbox_3_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T1), 
        .A2(SubBytesIns_Inst_Sbox_3_T15), .ZN(SubBytesIns_Inst_Sbox_3_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T4), 
        .A2(SubBytesIns_Inst_Sbox_3_T27), .ZN(SubBytesIns_Inst_Sbox_3_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_3_M12), 
        .B(SubBytesIns_Inst_Sbox_3_M11), .Z(SubBytesIns_Inst_Sbox_3_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T2), 
        .A2(SubBytesIns_Inst_Sbox_3_T10), .ZN(SubBytesIns_Inst_Sbox_3_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_3_M14), 
        .B(SubBytesIns_Inst_Sbox_3_M11), .Z(SubBytesIns_Inst_Sbox_3_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_3_M3), 
        .B(SubBytesIns_Inst_Sbox_3_M2), .Z(SubBytesIns_Inst_Sbox_3_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_3_M5), 
        .B(SubBytesIns_Inst_Sbox_3_T24), .Z(SubBytesIns_Inst_Sbox_3_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_3_M8), 
        .B(SubBytesIns_Inst_Sbox_3_M7), .Z(SubBytesIns_Inst_Sbox_3_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_3_M10), 
        .B(SubBytesIns_Inst_Sbox_3_M15), .Z(SubBytesIns_Inst_Sbox_3_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_3_M16), 
        .B(SubBytesIns_Inst_Sbox_3_M13), .Z(SubBytesIns_Inst_Sbox_3_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_3_M17), 
        .B(SubBytesIns_Inst_Sbox_3_M15), .Z(SubBytesIns_Inst_Sbox_3_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_3_M18), 
        .B(SubBytesIns_Inst_Sbox_3_M13), .Z(SubBytesIns_Inst_Sbox_3_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_3_M19), 
        .B(SubBytesIns_Inst_Sbox_3_T25), .Z(SubBytesIns_Inst_Sbox_3_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_3_M22), 
        .B(SubBytesIns_Inst_Sbox_3_M23), .Z(SubBytesIns_Inst_Sbox_3_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M22), .A2(SubBytesIns_Inst_Sbox_3_M20), .ZN(SubBytesIns_Inst_Sbox_3_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_3_M21), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_3_M20), 
        .B(SubBytesIns_Inst_Sbox_3_M21), .Z(SubBytesIns_Inst_Sbox_3_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_3_M23), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M28), .A2(SubBytesIns_Inst_Sbox_3_M27), .ZN(SubBytesIns_Inst_Sbox_3_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M26), .A2(SubBytesIns_Inst_Sbox_3_M24), .ZN(SubBytesIns_Inst_Sbox_3_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M20), .A2(SubBytesIns_Inst_Sbox_3_M23), .ZN(SubBytesIns_Inst_Sbox_3_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M27), .A2(SubBytesIns_Inst_Sbox_3_M31), .ZN(SubBytesIns_Inst_Sbox_3_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_3_M27), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M21), .A2(SubBytesIns_Inst_Sbox_3_M22), .ZN(SubBytesIns_Inst_Sbox_3_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M24), .A2(SubBytesIns_Inst_Sbox_3_M34), .ZN(SubBytesIns_Inst_Sbox_3_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_3_M24), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_3_M21), 
        .B(SubBytesIns_Inst_Sbox_3_M29), .Z(SubBytesIns_Inst_Sbox_3_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_3_M32), 
        .B(SubBytesIns_Inst_Sbox_3_M33), .Z(SubBytesIns_Inst_Sbox_3_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_3_M23), 
        .B(SubBytesIns_Inst_Sbox_3_M30), .Z(SubBytesIns_Inst_Sbox_3_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_3_M35), 
        .B(SubBytesIns_Inst_Sbox_3_M36), .Z(SubBytesIns_Inst_Sbox_3_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_3_M38), 
        .B(SubBytesIns_Inst_Sbox_3_M40), .Z(SubBytesIns_Inst_Sbox_3_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_3_M37), 
        .B(SubBytesIns_Inst_Sbox_3_M39), .Z(SubBytesIns_Inst_Sbox_3_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_3_M37), 
        .B(SubBytesIns_Inst_Sbox_3_M38), .Z(SubBytesIns_Inst_Sbox_3_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_3_M39), 
        .B(SubBytesIns_Inst_Sbox_3_M40), .Z(SubBytesIns_Inst_Sbox_3_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_3_M42), 
        .B(SubBytesIns_Inst_Sbox_3_M41), .Z(SubBytesIns_Inst_Sbox_3_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M44), .A2(SubBytesIns_Inst_Sbox_3_T6), .ZN(SubBytesIns_Inst_Sbox_3_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M40), .A2(SubBytesIns_Inst_Sbox_3_T8), .ZN(SubBytesIns_Inst_Sbox_3_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M39), .A2(ciphertext[24]), .ZN(SubBytesIns_Inst_Sbox_3_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M43), .A2(SubBytesIns_Inst_Sbox_3_T16), .ZN(SubBytesIns_Inst_Sbox_3_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M38), .A2(SubBytesIns_Inst_Sbox_3_T9), .ZN(SubBytesIns_Inst_Sbox_3_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M37), .A2(SubBytesIns_Inst_Sbox_3_T17), .ZN(SubBytesIns_Inst_Sbox_3_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M42), .A2(SubBytesIns_Inst_Sbox_3_T15), .ZN(SubBytesIns_Inst_Sbox_3_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M45), .A2(SubBytesIns_Inst_Sbox_3_T27), .ZN(SubBytesIns_Inst_Sbox_3_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M41), .A2(SubBytesIns_Inst_Sbox_3_T10), .ZN(SubBytesIns_Inst_Sbox_3_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M44), .A2(SubBytesIns_Inst_Sbox_3_T13), .ZN(SubBytesIns_Inst_Sbox_3_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M40), .A2(SubBytesIns_Inst_Sbox_3_T23), .ZN(SubBytesIns_Inst_Sbox_3_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M39), .A2(SubBytesIns_Inst_Sbox_3_T19), .ZN(SubBytesIns_Inst_Sbox_3_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M43), .A2(SubBytesIns_Inst_Sbox_3_T3), .ZN(SubBytesIns_Inst_Sbox_3_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M38), .A2(SubBytesIns_Inst_Sbox_3_T22), .ZN(SubBytesIns_Inst_Sbox_3_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M37), .A2(SubBytesIns_Inst_Sbox_3_T20), .ZN(SubBytesIns_Inst_Sbox_3_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M42), .A2(SubBytesIns_Inst_Sbox_3_T1), .ZN(SubBytesIns_Inst_Sbox_3_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M45), .A2(SubBytesIns_Inst_Sbox_3_T4), .ZN(SubBytesIns_Inst_Sbox_3_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M41), .A2(SubBytesIns_Inst_Sbox_3_T2), .ZN(SubBytesIns_Inst_Sbox_3_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_3_M61), 
        .B(SubBytesIns_Inst_Sbox_3_M62), .Z(SubBytesIns_Inst_Sbox_3_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_3_M50), 
        .B(SubBytesIns_Inst_Sbox_3_M56), .Z(SubBytesIns_Inst_Sbox_3_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_3_M46), 
        .B(SubBytesIns_Inst_Sbox_3_M48), .Z(SubBytesIns_Inst_Sbox_3_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_3_M47), 
        .B(SubBytesIns_Inst_Sbox_3_M55), .Z(SubBytesIns_Inst_Sbox_3_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_3_M54), 
        .B(SubBytesIns_Inst_Sbox_3_M58), .Z(SubBytesIns_Inst_Sbox_3_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_3_M49), 
        .B(SubBytesIns_Inst_Sbox_3_M61), .Z(SubBytesIns_Inst_Sbox_3_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_3_M62), 
        .B(SubBytesIns_Inst_Sbox_3_L5), .Z(SubBytesIns_Inst_Sbox_3_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_3_M46), 
        .B(SubBytesIns_Inst_Sbox_3_L3), .Z(SubBytesIns_Inst_Sbox_3_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_3_M51), 
        .B(SubBytesIns_Inst_Sbox_3_M59), .Z(SubBytesIns_Inst_Sbox_3_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_3_M52), 
        .B(SubBytesIns_Inst_Sbox_3_M53), .Z(SubBytesIns_Inst_Sbox_3_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_3_M53), 
        .B(SubBytesIns_Inst_Sbox_3_L4), .Z(SubBytesIns_Inst_Sbox_3_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_3_M60), 
        .B(SubBytesIns_Inst_Sbox_3_L2), .Z(SubBytesIns_Inst_Sbox_3_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_3_M48), 
        .B(SubBytesIns_Inst_Sbox_3_M51), .Z(SubBytesIns_Inst_Sbox_3_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_3_M50), 
        .B(SubBytesIns_Inst_Sbox_3_L0), .Z(SubBytesIns_Inst_Sbox_3_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_3_M52), 
        .B(SubBytesIns_Inst_Sbox_3_M61), .Z(SubBytesIns_Inst_Sbox_3_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_3_M55), 
        .B(SubBytesIns_Inst_Sbox_3_L1), .Z(SubBytesIns_Inst_Sbox_3_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_3_M56), 
        .B(SubBytesIns_Inst_Sbox_3_L0), .Z(SubBytesIns_Inst_Sbox_3_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_3_M57), 
        .B(SubBytesIns_Inst_Sbox_3_L1), .Z(SubBytesIns_Inst_Sbox_3_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_3_M58), 
        .B(SubBytesIns_Inst_Sbox_3_L8), .Z(SubBytesIns_Inst_Sbox_3_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_3_M63), 
        .B(SubBytesIns_Inst_Sbox_3_L4), .Z(SubBytesIns_Inst_Sbox_3_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_3_L0), 
        .B(SubBytesIns_Inst_Sbox_3_L1), .Z(SubBytesIns_Inst_Sbox_3_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_3_L1), 
        .B(SubBytesIns_Inst_Sbox_3_L7), .Z(SubBytesIns_Inst_Sbox_3_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_3_L3), 
        .B(SubBytesIns_Inst_Sbox_3_L12), .Z(SubBytesIns_Inst_Sbox_3_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_3_L18), 
        .B(SubBytesIns_Inst_Sbox_3_L2), .Z(SubBytesIns_Inst_Sbox_3_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_3_L15), 
        .B(SubBytesIns_Inst_Sbox_3_L9), .Z(SubBytesIns_Inst_Sbox_3_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L10), .Z(SubBytesIns_Inst_Sbox_3_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_3_L7), 
        .B(SubBytesIns_Inst_Sbox_3_L9), .Z(SubBytesIns_Inst_Sbox_3_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_3_L8), 
        .B(SubBytesIns_Inst_Sbox_3_L10), .Z(SubBytesIns_Inst_Sbox_3_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_3_L11), 
        .B(SubBytesIns_Inst_Sbox_3_L14), .Z(SubBytesIns_Inst_Sbox_3_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_3_L11), 
        .B(SubBytesIns_Inst_Sbox_3_L17), .Z(SubBytesIns_Inst_Sbox_3_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L24), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_3_L16), 
        .B(SubBytesIns_Inst_Sbox_3_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_3_L19), 
        .B(SubBytesIns_Inst_Sbox_3_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L21), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_3_L20), 
        .B(SubBytesIns_Inst_Sbox_3_L22), .Z(MixColumnsInput[27]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_3_L25), 
        .B(SubBytesIns_Inst_Sbox_3_L29), .Z(MixColumnsInput[26]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_3_L13), 
        .B(SubBytesIns_Inst_Sbox_3_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L23), .ZN(MixColumnsInput[24]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T1_U1 ( .A(ciphertext[39]), .B(
        ciphertext[36]), .Z(SubBytesIns_Inst_Sbox_4_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T2_U1 ( .A(ciphertext[39]), .B(
        ciphertext[34]), .Z(SubBytesIns_Inst_Sbox_4_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T3_U1 ( .A(ciphertext[39]), .B(
        ciphertext[33]), .Z(SubBytesIns_Inst_Sbox_4_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T4_U1 ( .A(ciphertext[36]), .B(
        ciphertext[34]), .Z(SubBytesIns_Inst_Sbox_4_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T5_U1 ( .A(ciphertext[35]), .B(
        ciphertext[33]), .Z(SubBytesIns_Inst_Sbox_4_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_4_T1), 
        .B(SubBytesIns_Inst_Sbox_4_T5), .Z(SubBytesIns_Inst_Sbox_4_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T7_U1 ( .A(ciphertext[38]), .B(
        ciphertext[37]), .Z(SubBytesIns_Inst_Sbox_4_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T8_U1 ( .A(ciphertext[32]), .B(
        SubBytesIns_Inst_Sbox_4_T6), .Z(SubBytesIns_Inst_Sbox_4_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T9_U1 ( .A(ciphertext[32]), .B(
        SubBytesIns_Inst_Sbox_4_T7), .Z(SubBytesIns_Inst_Sbox_4_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_4_T6), 
        .B(SubBytesIns_Inst_Sbox_4_T7), .Z(SubBytesIns_Inst_Sbox_4_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T11_U1 ( .A(ciphertext[38]), .B(
        ciphertext[34]), .Z(SubBytesIns_Inst_Sbox_4_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T12_U1 ( .A(ciphertext[37]), .B(
        ciphertext[34]), .Z(SubBytesIns_Inst_Sbox_4_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_4_T3), 
        .B(SubBytesIns_Inst_Sbox_4_T4), .Z(SubBytesIns_Inst_Sbox_4_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_4_T6), 
        .B(SubBytesIns_Inst_Sbox_4_T11), .Z(SubBytesIns_Inst_Sbox_4_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_4_T5), 
        .B(SubBytesIns_Inst_Sbox_4_T11), .Z(SubBytesIns_Inst_Sbox_4_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_4_T5), 
        .B(SubBytesIns_Inst_Sbox_4_T12), .Z(SubBytesIns_Inst_Sbox_4_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_4_T9), 
        .B(SubBytesIns_Inst_Sbox_4_T16), .Z(SubBytesIns_Inst_Sbox_4_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T18_U1 ( .A(ciphertext[36]), .B(
        ciphertext[32]), .Z(SubBytesIns_Inst_Sbox_4_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_4_T7), 
        .B(SubBytesIns_Inst_Sbox_4_T18), .Z(SubBytesIns_Inst_Sbox_4_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_4_T1), 
        .B(SubBytesIns_Inst_Sbox_4_T19), .Z(SubBytesIns_Inst_Sbox_4_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T21_U1 ( .A(ciphertext[33]), .B(
        ciphertext[32]), .Z(SubBytesIns_Inst_Sbox_4_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_4_T7), 
        .B(SubBytesIns_Inst_Sbox_4_T21), .Z(SubBytesIns_Inst_Sbox_4_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_4_T2), 
        .B(SubBytesIns_Inst_Sbox_4_T22), .Z(SubBytesIns_Inst_Sbox_4_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_4_T2), 
        .B(SubBytesIns_Inst_Sbox_4_T10), .Z(SubBytesIns_Inst_Sbox_4_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_4_T20), 
        .B(SubBytesIns_Inst_Sbox_4_T17), .Z(SubBytesIns_Inst_Sbox_4_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_4_T3), 
        .B(SubBytesIns_Inst_Sbox_4_T16), .Z(SubBytesIns_Inst_Sbox_4_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_4_T1), 
        .B(SubBytesIns_Inst_Sbox_4_T12), .Z(SubBytesIns_Inst_Sbox_4_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T13), 
        .A2(SubBytesIns_Inst_Sbox_4_T6), .ZN(SubBytesIns_Inst_Sbox_4_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T23), 
        .A2(SubBytesIns_Inst_Sbox_4_T8), .ZN(SubBytesIns_Inst_Sbox_4_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_4_T14), 
        .B(SubBytesIns_Inst_Sbox_4_M1), .Z(SubBytesIns_Inst_Sbox_4_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T19), 
        .A2(ciphertext[32]), .ZN(SubBytesIns_Inst_Sbox_4_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_4_M4), 
        .B(SubBytesIns_Inst_Sbox_4_M1), .Z(SubBytesIns_Inst_Sbox_4_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T3), 
        .A2(SubBytesIns_Inst_Sbox_4_T16), .ZN(SubBytesIns_Inst_Sbox_4_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T22), 
        .A2(SubBytesIns_Inst_Sbox_4_T9), .ZN(SubBytesIns_Inst_Sbox_4_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_4_T26), 
        .B(SubBytesIns_Inst_Sbox_4_M6), .Z(SubBytesIns_Inst_Sbox_4_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T20), 
        .A2(SubBytesIns_Inst_Sbox_4_T17), .ZN(SubBytesIns_Inst_Sbox_4_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_4_M9), 
        .B(SubBytesIns_Inst_Sbox_4_M6), .Z(SubBytesIns_Inst_Sbox_4_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T1), 
        .A2(SubBytesIns_Inst_Sbox_4_T15), .ZN(SubBytesIns_Inst_Sbox_4_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T4), 
        .A2(SubBytesIns_Inst_Sbox_4_T27), .ZN(SubBytesIns_Inst_Sbox_4_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_4_M12), 
        .B(SubBytesIns_Inst_Sbox_4_M11), .Z(SubBytesIns_Inst_Sbox_4_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T2), 
        .A2(SubBytesIns_Inst_Sbox_4_T10), .ZN(SubBytesIns_Inst_Sbox_4_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_4_M14), 
        .B(SubBytesIns_Inst_Sbox_4_M11), .Z(SubBytesIns_Inst_Sbox_4_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_4_M3), 
        .B(SubBytesIns_Inst_Sbox_4_M2), .Z(SubBytesIns_Inst_Sbox_4_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_4_M5), 
        .B(SubBytesIns_Inst_Sbox_4_T24), .Z(SubBytesIns_Inst_Sbox_4_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_4_M8), 
        .B(SubBytesIns_Inst_Sbox_4_M7), .Z(SubBytesIns_Inst_Sbox_4_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_4_M10), 
        .B(SubBytesIns_Inst_Sbox_4_M15), .Z(SubBytesIns_Inst_Sbox_4_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_4_M16), 
        .B(SubBytesIns_Inst_Sbox_4_M13), .Z(SubBytesIns_Inst_Sbox_4_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_4_M17), 
        .B(SubBytesIns_Inst_Sbox_4_M15), .Z(SubBytesIns_Inst_Sbox_4_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_4_M18), 
        .B(SubBytesIns_Inst_Sbox_4_M13), .Z(SubBytesIns_Inst_Sbox_4_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_4_M19), 
        .B(SubBytesIns_Inst_Sbox_4_T25), .Z(SubBytesIns_Inst_Sbox_4_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_4_M22), 
        .B(SubBytesIns_Inst_Sbox_4_M23), .Z(SubBytesIns_Inst_Sbox_4_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M22), .A2(SubBytesIns_Inst_Sbox_4_M20), .ZN(SubBytesIns_Inst_Sbox_4_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_4_M21), 
        .B(SubBytesIns_Inst_Sbox_4_M25), .Z(SubBytesIns_Inst_Sbox_4_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_4_M20), 
        .B(SubBytesIns_Inst_Sbox_4_M21), .Z(SubBytesIns_Inst_Sbox_4_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_4_M23), 
        .B(SubBytesIns_Inst_Sbox_4_M25), .Z(SubBytesIns_Inst_Sbox_4_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M28), .A2(SubBytesIns_Inst_Sbox_4_M27), .ZN(SubBytesIns_Inst_Sbox_4_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M26), .A2(SubBytesIns_Inst_Sbox_4_M24), .ZN(SubBytesIns_Inst_Sbox_4_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M20), .A2(SubBytesIns_Inst_Sbox_4_M23), .ZN(SubBytesIns_Inst_Sbox_4_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M27), .A2(SubBytesIns_Inst_Sbox_4_M31), .ZN(SubBytesIns_Inst_Sbox_4_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_4_M27), 
        .B(SubBytesIns_Inst_Sbox_4_M25), .Z(SubBytesIns_Inst_Sbox_4_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M21), .A2(SubBytesIns_Inst_Sbox_4_M22), .ZN(SubBytesIns_Inst_Sbox_4_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M24), .A2(SubBytesIns_Inst_Sbox_4_M34), .ZN(SubBytesIns_Inst_Sbox_4_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_4_M24), 
        .B(SubBytesIns_Inst_Sbox_4_M25), .Z(SubBytesIns_Inst_Sbox_4_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_4_M21), 
        .B(SubBytesIns_Inst_Sbox_4_M29), .Z(SubBytesIns_Inst_Sbox_4_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_4_M32), 
        .B(SubBytesIns_Inst_Sbox_4_M33), .Z(SubBytesIns_Inst_Sbox_4_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_4_M23), 
        .B(SubBytesIns_Inst_Sbox_4_M30), .Z(SubBytesIns_Inst_Sbox_4_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_4_M35), 
        .B(SubBytesIns_Inst_Sbox_4_M36), .Z(SubBytesIns_Inst_Sbox_4_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_4_M38), 
        .B(SubBytesIns_Inst_Sbox_4_M40), .Z(SubBytesIns_Inst_Sbox_4_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_4_M37), 
        .B(SubBytesIns_Inst_Sbox_4_M39), .Z(SubBytesIns_Inst_Sbox_4_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_4_M37), 
        .B(SubBytesIns_Inst_Sbox_4_M38), .Z(SubBytesIns_Inst_Sbox_4_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_4_M39), 
        .B(SubBytesIns_Inst_Sbox_4_M40), .Z(SubBytesIns_Inst_Sbox_4_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_4_M42), 
        .B(SubBytesIns_Inst_Sbox_4_M41), .Z(SubBytesIns_Inst_Sbox_4_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M44), .A2(SubBytesIns_Inst_Sbox_4_T6), .ZN(SubBytesIns_Inst_Sbox_4_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M40), .A2(SubBytesIns_Inst_Sbox_4_T8), .ZN(SubBytesIns_Inst_Sbox_4_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M39), .A2(ciphertext[32]), .ZN(SubBytesIns_Inst_Sbox_4_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M43), .A2(SubBytesIns_Inst_Sbox_4_T16), .ZN(SubBytesIns_Inst_Sbox_4_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M38), .A2(SubBytesIns_Inst_Sbox_4_T9), .ZN(SubBytesIns_Inst_Sbox_4_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M37), .A2(SubBytesIns_Inst_Sbox_4_T17), .ZN(SubBytesIns_Inst_Sbox_4_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M42), .A2(SubBytesIns_Inst_Sbox_4_T15), .ZN(SubBytesIns_Inst_Sbox_4_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M45), .A2(SubBytesIns_Inst_Sbox_4_T27), .ZN(SubBytesIns_Inst_Sbox_4_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M41), .A2(SubBytesIns_Inst_Sbox_4_T10), .ZN(SubBytesIns_Inst_Sbox_4_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M44), .A2(SubBytesIns_Inst_Sbox_4_T13), .ZN(SubBytesIns_Inst_Sbox_4_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M40), .A2(SubBytesIns_Inst_Sbox_4_T23), .ZN(SubBytesIns_Inst_Sbox_4_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M39), .A2(SubBytesIns_Inst_Sbox_4_T19), .ZN(SubBytesIns_Inst_Sbox_4_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M43), .A2(SubBytesIns_Inst_Sbox_4_T3), .ZN(SubBytesIns_Inst_Sbox_4_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M38), .A2(SubBytesIns_Inst_Sbox_4_T22), .ZN(SubBytesIns_Inst_Sbox_4_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M37), .A2(SubBytesIns_Inst_Sbox_4_T20), .ZN(SubBytesIns_Inst_Sbox_4_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M42), .A2(SubBytesIns_Inst_Sbox_4_T1), .ZN(SubBytesIns_Inst_Sbox_4_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M45), .A2(SubBytesIns_Inst_Sbox_4_T4), .ZN(SubBytesIns_Inst_Sbox_4_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M41), .A2(SubBytesIns_Inst_Sbox_4_T2), .ZN(SubBytesIns_Inst_Sbox_4_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_4_M61), 
        .B(SubBytesIns_Inst_Sbox_4_M62), .Z(SubBytesIns_Inst_Sbox_4_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_4_M50), 
        .B(SubBytesIns_Inst_Sbox_4_M56), .Z(SubBytesIns_Inst_Sbox_4_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_4_M46), 
        .B(SubBytesIns_Inst_Sbox_4_M48), .Z(SubBytesIns_Inst_Sbox_4_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_4_M47), 
        .B(SubBytesIns_Inst_Sbox_4_M55), .Z(SubBytesIns_Inst_Sbox_4_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_4_M54), 
        .B(SubBytesIns_Inst_Sbox_4_M58), .Z(SubBytesIns_Inst_Sbox_4_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_4_M49), 
        .B(SubBytesIns_Inst_Sbox_4_M61), .Z(SubBytesIns_Inst_Sbox_4_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_4_M62), 
        .B(SubBytesIns_Inst_Sbox_4_L5), .Z(SubBytesIns_Inst_Sbox_4_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_4_M46), 
        .B(SubBytesIns_Inst_Sbox_4_L3), .Z(SubBytesIns_Inst_Sbox_4_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_4_M51), 
        .B(SubBytesIns_Inst_Sbox_4_M59), .Z(SubBytesIns_Inst_Sbox_4_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_4_M52), 
        .B(SubBytesIns_Inst_Sbox_4_M53), .Z(SubBytesIns_Inst_Sbox_4_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_4_M53), 
        .B(SubBytesIns_Inst_Sbox_4_L4), .Z(SubBytesIns_Inst_Sbox_4_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_4_M60), 
        .B(SubBytesIns_Inst_Sbox_4_L2), .Z(SubBytesIns_Inst_Sbox_4_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_4_M48), 
        .B(SubBytesIns_Inst_Sbox_4_M51), .Z(SubBytesIns_Inst_Sbox_4_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_4_M50), 
        .B(SubBytesIns_Inst_Sbox_4_L0), .Z(SubBytesIns_Inst_Sbox_4_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_4_M52), 
        .B(SubBytesIns_Inst_Sbox_4_M61), .Z(SubBytesIns_Inst_Sbox_4_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_4_M55), 
        .B(SubBytesIns_Inst_Sbox_4_L1), .Z(SubBytesIns_Inst_Sbox_4_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_4_M56), 
        .B(SubBytesIns_Inst_Sbox_4_L0), .Z(SubBytesIns_Inst_Sbox_4_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_4_M57), 
        .B(SubBytesIns_Inst_Sbox_4_L1), .Z(SubBytesIns_Inst_Sbox_4_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_4_M58), 
        .B(SubBytesIns_Inst_Sbox_4_L8), .Z(SubBytesIns_Inst_Sbox_4_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_4_M63), 
        .B(SubBytesIns_Inst_Sbox_4_L4), .Z(SubBytesIns_Inst_Sbox_4_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_4_L0), 
        .B(SubBytesIns_Inst_Sbox_4_L1), .Z(SubBytesIns_Inst_Sbox_4_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_4_L1), 
        .B(SubBytesIns_Inst_Sbox_4_L7), .Z(SubBytesIns_Inst_Sbox_4_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_4_L3), 
        .B(SubBytesIns_Inst_Sbox_4_L12), .Z(SubBytesIns_Inst_Sbox_4_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_4_L18), 
        .B(SubBytesIns_Inst_Sbox_4_L2), .Z(SubBytesIns_Inst_Sbox_4_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_4_L15), 
        .B(SubBytesIns_Inst_Sbox_4_L9), .Z(SubBytesIns_Inst_Sbox_4_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_4_L6), 
        .B(SubBytesIns_Inst_Sbox_4_L10), .Z(SubBytesIns_Inst_Sbox_4_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_4_L7), 
        .B(SubBytesIns_Inst_Sbox_4_L9), .Z(SubBytesIns_Inst_Sbox_4_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_4_L8), 
        .B(SubBytesIns_Inst_Sbox_4_L10), .Z(SubBytesIns_Inst_Sbox_4_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_4_L11), 
        .B(SubBytesIns_Inst_Sbox_4_L14), .Z(SubBytesIns_Inst_Sbox_4_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_4_L11), 
        .B(SubBytesIns_Inst_Sbox_4_L17), .Z(SubBytesIns_Inst_Sbox_4_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_4_L6), 
        .B(SubBytesIns_Inst_Sbox_4_L24), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_4_L16), 
        .B(SubBytesIns_Inst_Sbox_4_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_4_L19), 
        .B(SubBytesIns_Inst_Sbox_4_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_4_L6), 
        .B(SubBytesIns_Inst_Sbox_4_L21), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_4_L20), 
        .B(SubBytesIns_Inst_Sbox_4_L22), .Z(MixColumnsInput[3]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_4_L25), 
        .B(SubBytesIns_Inst_Sbox_4_L29), .Z(MixColumnsInput[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_4_L13), 
        .B(SubBytesIns_Inst_Sbox_4_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_4_L6), 
        .B(SubBytesIns_Inst_Sbox_4_L23), .ZN(MixColumnsInput[0]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T1_U1 ( .A(ciphertext[47]), .B(
        ciphertext[44]), .Z(SubBytesIns_Inst_Sbox_5_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T2_U1 ( .A(ciphertext[47]), .B(
        ciphertext[42]), .Z(SubBytesIns_Inst_Sbox_5_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T3_U1 ( .A(ciphertext[47]), .B(
        ciphertext[41]), .Z(SubBytesIns_Inst_Sbox_5_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T4_U1 ( .A(ciphertext[44]), .B(
        ciphertext[42]), .Z(SubBytesIns_Inst_Sbox_5_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T5_U1 ( .A(ciphertext[43]), .B(
        ciphertext[41]), .Z(SubBytesIns_Inst_Sbox_5_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_5_T1), 
        .B(SubBytesIns_Inst_Sbox_5_T5), .Z(SubBytesIns_Inst_Sbox_5_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T7_U1 ( .A(ciphertext[46]), .B(
        ciphertext[45]), .Z(SubBytesIns_Inst_Sbox_5_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T8_U1 ( .A(ciphertext[40]), .B(
        SubBytesIns_Inst_Sbox_5_T6), .Z(SubBytesIns_Inst_Sbox_5_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T9_U1 ( .A(ciphertext[40]), .B(
        SubBytesIns_Inst_Sbox_5_T7), .Z(SubBytesIns_Inst_Sbox_5_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_5_T6), 
        .B(SubBytesIns_Inst_Sbox_5_T7), .Z(SubBytesIns_Inst_Sbox_5_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T11_U1 ( .A(ciphertext[46]), .B(
        ciphertext[42]), .Z(SubBytesIns_Inst_Sbox_5_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T12_U1 ( .A(ciphertext[45]), .B(
        ciphertext[42]), .Z(SubBytesIns_Inst_Sbox_5_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_5_T3), 
        .B(SubBytesIns_Inst_Sbox_5_T4), .Z(SubBytesIns_Inst_Sbox_5_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_5_T6), 
        .B(SubBytesIns_Inst_Sbox_5_T11), .Z(SubBytesIns_Inst_Sbox_5_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_5_T5), 
        .B(SubBytesIns_Inst_Sbox_5_T11), .Z(SubBytesIns_Inst_Sbox_5_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_5_T5), 
        .B(SubBytesIns_Inst_Sbox_5_T12), .Z(SubBytesIns_Inst_Sbox_5_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_5_T9), 
        .B(SubBytesIns_Inst_Sbox_5_T16), .Z(SubBytesIns_Inst_Sbox_5_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T18_U1 ( .A(ciphertext[44]), .B(
        ciphertext[40]), .Z(SubBytesIns_Inst_Sbox_5_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_5_T7), 
        .B(SubBytesIns_Inst_Sbox_5_T18), .Z(SubBytesIns_Inst_Sbox_5_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_5_T1), 
        .B(SubBytesIns_Inst_Sbox_5_T19), .Z(SubBytesIns_Inst_Sbox_5_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T21_U1 ( .A(ciphertext[41]), .B(
        ciphertext[40]), .Z(SubBytesIns_Inst_Sbox_5_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_5_T7), 
        .B(SubBytesIns_Inst_Sbox_5_T21), .Z(SubBytesIns_Inst_Sbox_5_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_5_T2), 
        .B(SubBytesIns_Inst_Sbox_5_T22), .Z(SubBytesIns_Inst_Sbox_5_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_5_T2), 
        .B(SubBytesIns_Inst_Sbox_5_T10), .Z(SubBytesIns_Inst_Sbox_5_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_5_T20), 
        .B(SubBytesIns_Inst_Sbox_5_T17), .Z(SubBytesIns_Inst_Sbox_5_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_5_T3), 
        .B(SubBytesIns_Inst_Sbox_5_T16), .Z(SubBytesIns_Inst_Sbox_5_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_5_T1), 
        .B(SubBytesIns_Inst_Sbox_5_T12), .Z(SubBytesIns_Inst_Sbox_5_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T13), 
        .A2(SubBytesIns_Inst_Sbox_5_T6), .ZN(SubBytesIns_Inst_Sbox_5_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T23), 
        .A2(SubBytesIns_Inst_Sbox_5_T8), .ZN(SubBytesIns_Inst_Sbox_5_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_5_T14), 
        .B(SubBytesIns_Inst_Sbox_5_M1), .Z(SubBytesIns_Inst_Sbox_5_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T19), 
        .A2(ciphertext[40]), .ZN(SubBytesIns_Inst_Sbox_5_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_5_M4), 
        .B(SubBytesIns_Inst_Sbox_5_M1), .Z(SubBytesIns_Inst_Sbox_5_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T3), 
        .A2(SubBytesIns_Inst_Sbox_5_T16), .ZN(SubBytesIns_Inst_Sbox_5_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T22), 
        .A2(SubBytesIns_Inst_Sbox_5_T9), .ZN(SubBytesIns_Inst_Sbox_5_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_5_T26), 
        .B(SubBytesIns_Inst_Sbox_5_M6), .Z(SubBytesIns_Inst_Sbox_5_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T20), 
        .A2(SubBytesIns_Inst_Sbox_5_T17), .ZN(SubBytesIns_Inst_Sbox_5_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_5_M9), 
        .B(SubBytesIns_Inst_Sbox_5_M6), .Z(SubBytesIns_Inst_Sbox_5_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T1), 
        .A2(SubBytesIns_Inst_Sbox_5_T15), .ZN(SubBytesIns_Inst_Sbox_5_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T4), 
        .A2(SubBytesIns_Inst_Sbox_5_T27), .ZN(SubBytesIns_Inst_Sbox_5_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_5_M12), 
        .B(SubBytesIns_Inst_Sbox_5_M11), .Z(SubBytesIns_Inst_Sbox_5_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T2), 
        .A2(SubBytesIns_Inst_Sbox_5_T10), .ZN(SubBytesIns_Inst_Sbox_5_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_5_M14), 
        .B(SubBytesIns_Inst_Sbox_5_M11), .Z(SubBytesIns_Inst_Sbox_5_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_5_M3), 
        .B(SubBytesIns_Inst_Sbox_5_M2), .Z(SubBytesIns_Inst_Sbox_5_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_5_M5), 
        .B(SubBytesIns_Inst_Sbox_5_T24), .Z(SubBytesIns_Inst_Sbox_5_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_5_M8), 
        .B(SubBytesIns_Inst_Sbox_5_M7), .Z(SubBytesIns_Inst_Sbox_5_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_5_M10), 
        .B(SubBytesIns_Inst_Sbox_5_M15), .Z(SubBytesIns_Inst_Sbox_5_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_5_M16), 
        .B(SubBytesIns_Inst_Sbox_5_M13), .Z(SubBytesIns_Inst_Sbox_5_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_5_M17), 
        .B(SubBytesIns_Inst_Sbox_5_M15), .Z(SubBytesIns_Inst_Sbox_5_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_5_M18), 
        .B(SubBytesIns_Inst_Sbox_5_M13), .Z(SubBytesIns_Inst_Sbox_5_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_5_M19), 
        .B(SubBytesIns_Inst_Sbox_5_T25), .Z(SubBytesIns_Inst_Sbox_5_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_5_M22), 
        .B(SubBytesIns_Inst_Sbox_5_M23), .Z(SubBytesIns_Inst_Sbox_5_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M22), .A2(SubBytesIns_Inst_Sbox_5_M20), .ZN(SubBytesIns_Inst_Sbox_5_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_5_M21), 
        .B(SubBytesIns_Inst_Sbox_5_M25), .Z(SubBytesIns_Inst_Sbox_5_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_5_M20), 
        .B(SubBytesIns_Inst_Sbox_5_M21), .Z(SubBytesIns_Inst_Sbox_5_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_5_M23), 
        .B(SubBytesIns_Inst_Sbox_5_M25), .Z(SubBytesIns_Inst_Sbox_5_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M28), .A2(SubBytesIns_Inst_Sbox_5_M27), .ZN(SubBytesIns_Inst_Sbox_5_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M26), .A2(SubBytesIns_Inst_Sbox_5_M24), .ZN(SubBytesIns_Inst_Sbox_5_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M20), .A2(SubBytesIns_Inst_Sbox_5_M23), .ZN(SubBytesIns_Inst_Sbox_5_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M27), .A2(SubBytesIns_Inst_Sbox_5_M31), .ZN(SubBytesIns_Inst_Sbox_5_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_5_M27), 
        .B(SubBytesIns_Inst_Sbox_5_M25), .Z(SubBytesIns_Inst_Sbox_5_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M21), .A2(SubBytesIns_Inst_Sbox_5_M22), .ZN(SubBytesIns_Inst_Sbox_5_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M24), .A2(SubBytesIns_Inst_Sbox_5_M34), .ZN(SubBytesIns_Inst_Sbox_5_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_5_M24), 
        .B(SubBytesIns_Inst_Sbox_5_M25), .Z(SubBytesIns_Inst_Sbox_5_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_5_M21), 
        .B(SubBytesIns_Inst_Sbox_5_M29), .Z(SubBytesIns_Inst_Sbox_5_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_5_M32), 
        .B(SubBytesIns_Inst_Sbox_5_M33), .Z(SubBytesIns_Inst_Sbox_5_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_5_M23), 
        .B(SubBytesIns_Inst_Sbox_5_M30), .Z(SubBytesIns_Inst_Sbox_5_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_5_M35), 
        .B(SubBytesIns_Inst_Sbox_5_M36), .Z(SubBytesIns_Inst_Sbox_5_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_5_M38), 
        .B(SubBytesIns_Inst_Sbox_5_M40), .Z(SubBytesIns_Inst_Sbox_5_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_5_M37), 
        .B(SubBytesIns_Inst_Sbox_5_M39), .Z(SubBytesIns_Inst_Sbox_5_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_5_M37), 
        .B(SubBytesIns_Inst_Sbox_5_M38), .Z(SubBytesIns_Inst_Sbox_5_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_5_M39), 
        .B(SubBytesIns_Inst_Sbox_5_M40), .Z(SubBytesIns_Inst_Sbox_5_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_5_M42), 
        .B(SubBytesIns_Inst_Sbox_5_M41), .Z(SubBytesIns_Inst_Sbox_5_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M44), .A2(SubBytesIns_Inst_Sbox_5_T6), .ZN(SubBytesIns_Inst_Sbox_5_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M40), .A2(SubBytesIns_Inst_Sbox_5_T8), .ZN(SubBytesIns_Inst_Sbox_5_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M39), .A2(ciphertext[40]), .ZN(SubBytesIns_Inst_Sbox_5_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M43), .A2(SubBytesIns_Inst_Sbox_5_T16), .ZN(SubBytesIns_Inst_Sbox_5_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M38), .A2(SubBytesIns_Inst_Sbox_5_T9), .ZN(SubBytesIns_Inst_Sbox_5_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M37), .A2(SubBytesIns_Inst_Sbox_5_T17), .ZN(SubBytesIns_Inst_Sbox_5_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M42), .A2(SubBytesIns_Inst_Sbox_5_T15), .ZN(SubBytesIns_Inst_Sbox_5_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M45), .A2(SubBytesIns_Inst_Sbox_5_T27), .ZN(SubBytesIns_Inst_Sbox_5_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M41), .A2(SubBytesIns_Inst_Sbox_5_T10), .ZN(SubBytesIns_Inst_Sbox_5_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M44), .A2(SubBytesIns_Inst_Sbox_5_T13), .ZN(SubBytesIns_Inst_Sbox_5_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M40), .A2(SubBytesIns_Inst_Sbox_5_T23), .ZN(SubBytesIns_Inst_Sbox_5_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M39), .A2(SubBytesIns_Inst_Sbox_5_T19), .ZN(SubBytesIns_Inst_Sbox_5_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M43), .A2(SubBytesIns_Inst_Sbox_5_T3), .ZN(SubBytesIns_Inst_Sbox_5_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M38), .A2(SubBytesIns_Inst_Sbox_5_T22), .ZN(SubBytesIns_Inst_Sbox_5_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M37), .A2(SubBytesIns_Inst_Sbox_5_T20), .ZN(SubBytesIns_Inst_Sbox_5_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M42), .A2(SubBytesIns_Inst_Sbox_5_T1), .ZN(SubBytesIns_Inst_Sbox_5_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M45), .A2(SubBytesIns_Inst_Sbox_5_T4), .ZN(SubBytesIns_Inst_Sbox_5_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M41), .A2(SubBytesIns_Inst_Sbox_5_T2), .ZN(SubBytesIns_Inst_Sbox_5_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_5_M61), 
        .B(SubBytesIns_Inst_Sbox_5_M62), .Z(SubBytesIns_Inst_Sbox_5_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_5_M50), 
        .B(SubBytesIns_Inst_Sbox_5_M56), .Z(SubBytesIns_Inst_Sbox_5_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_5_M46), 
        .B(SubBytesIns_Inst_Sbox_5_M48), .Z(SubBytesIns_Inst_Sbox_5_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_5_M47), 
        .B(SubBytesIns_Inst_Sbox_5_M55), .Z(SubBytesIns_Inst_Sbox_5_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_5_M54), 
        .B(SubBytesIns_Inst_Sbox_5_M58), .Z(SubBytesIns_Inst_Sbox_5_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_5_M49), 
        .B(SubBytesIns_Inst_Sbox_5_M61), .Z(SubBytesIns_Inst_Sbox_5_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_5_M62), 
        .B(SubBytesIns_Inst_Sbox_5_L5), .Z(SubBytesIns_Inst_Sbox_5_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_5_M46), 
        .B(SubBytesIns_Inst_Sbox_5_L3), .Z(SubBytesIns_Inst_Sbox_5_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_5_M51), 
        .B(SubBytesIns_Inst_Sbox_5_M59), .Z(SubBytesIns_Inst_Sbox_5_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_5_M52), 
        .B(SubBytesIns_Inst_Sbox_5_M53), .Z(SubBytesIns_Inst_Sbox_5_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_5_M53), 
        .B(SubBytesIns_Inst_Sbox_5_L4), .Z(SubBytesIns_Inst_Sbox_5_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_5_M60), 
        .B(SubBytesIns_Inst_Sbox_5_L2), .Z(SubBytesIns_Inst_Sbox_5_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_5_M48), 
        .B(SubBytesIns_Inst_Sbox_5_M51), .Z(SubBytesIns_Inst_Sbox_5_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_5_M50), 
        .B(SubBytesIns_Inst_Sbox_5_L0), .Z(SubBytesIns_Inst_Sbox_5_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_5_M52), 
        .B(SubBytesIns_Inst_Sbox_5_M61), .Z(SubBytesIns_Inst_Sbox_5_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_5_M55), 
        .B(SubBytesIns_Inst_Sbox_5_L1), .Z(SubBytesIns_Inst_Sbox_5_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_5_M56), 
        .B(SubBytesIns_Inst_Sbox_5_L0), .Z(SubBytesIns_Inst_Sbox_5_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_5_M57), 
        .B(SubBytesIns_Inst_Sbox_5_L1), .Z(SubBytesIns_Inst_Sbox_5_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_5_M58), 
        .B(SubBytesIns_Inst_Sbox_5_L8), .Z(SubBytesIns_Inst_Sbox_5_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_5_M63), 
        .B(SubBytesIns_Inst_Sbox_5_L4), .Z(SubBytesIns_Inst_Sbox_5_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_5_L0), 
        .B(SubBytesIns_Inst_Sbox_5_L1), .Z(SubBytesIns_Inst_Sbox_5_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_5_L1), 
        .B(SubBytesIns_Inst_Sbox_5_L7), .Z(SubBytesIns_Inst_Sbox_5_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_5_L3), 
        .B(SubBytesIns_Inst_Sbox_5_L12), .Z(SubBytesIns_Inst_Sbox_5_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_5_L18), 
        .B(SubBytesIns_Inst_Sbox_5_L2), .Z(SubBytesIns_Inst_Sbox_5_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_5_L15), 
        .B(SubBytesIns_Inst_Sbox_5_L9), .Z(SubBytesIns_Inst_Sbox_5_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_5_L6), 
        .B(SubBytesIns_Inst_Sbox_5_L10), .Z(SubBytesIns_Inst_Sbox_5_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_5_L7), 
        .B(SubBytesIns_Inst_Sbox_5_L9), .Z(SubBytesIns_Inst_Sbox_5_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_5_L8), 
        .B(SubBytesIns_Inst_Sbox_5_L10), .Z(SubBytesIns_Inst_Sbox_5_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_5_L11), 
        .B(SubBytesIns_Inst_Sbox_5_L14), .Z(SubBytesIns_Inst_Sbox_5_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_5_L11), 
        .B(SubBytesIns_Inst_Sbox_5_L17), .Z(SubBytesIns_Inst_Sbox_5_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_5_L6), 
        .B(SubBytesIns_Inst_Sbox_5_L24), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_5_L16), 
        .B(SubBytesIns_Inst_Sbox_5_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_5_L19), 
        .B(SubBytesIns_Inst_Sbox_5_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_5_L6), 
        .B(SubBytesIns_Inst_Sbox_5_L21), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_5_L20), 
        .B(SubBytesIns_Inst_Sbox_5_L22), .Z(MixColumnsInput[107]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_5_L25), 
        .B(SubBytesIns_Inst_Sbox_5_L29), .Z(MixColumnsInput[106]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_5_L13), 
        .B(SubBytesIns_Inst_Sbox_5_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_5_L6), 
        .B(SubBytesIns_Inst_Sbox_5_L23), .ZN(MixColumnsInput[104]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T1_U1 ( .A(ciphertext[55]), .B(
        ciphertext[52]), .Z(SubBytesIns_Inst_Sbox_6_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T2_U1 ( .A(ciphertext[55]), .B(
        ciphertext[50]), .Z(SubBytesIns_Inst_Sbox_6_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T3_U1 ( .A(ciphertext[55]), .B(
        ciphertext[49]), .Z(SubBytesIns_Inst_Sbox_6_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T4_U1 ( .A(ciphertext[52]), .B(
        ciphertext[50]), .Z(SubBytesIns_Inst_Sbox_6_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T5_U1 ( .A(ciphertext[51]), .B(
        ciphertext[49]), .Z(SubBytesIns_Inst_Sbox_6_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_6_T1), 
        .B(SubBytesIns_Inst_Sbox_6_T5), .Z(SubBytesIns_Inst_Sbox_6_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T7_U1 ( .A(ciphertext[54]), .B(
        ciphertext[53]), .Z(SubBytesIns_Inst_Sbox_6_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T8_U1 ( .A(ciphertext[48]), .B(
        SubBytesIns_Inst_Sbox_6_T6), .Z(SubBytesIns_Inst_Sbox_6_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T9_U1 ( .A(ciphertext[48]), .B(
        SubBytesIns_Inst_Sbox_6_T7), .Z(SubBytesIns_Inst_Sbox_6_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_6_T6), 
        .B(SubBytesIns_Inst_Sbox_6_T7), .Z(SubBytesIns_Inst_Sbox_6_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T11_U1 ( .A(ciphertext[54]), .B(
        ciphertext[50]), .Z(SubBytesIns_Inst_Sbox_6_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T12_U1 ( .A(ciphertext[53]), .B(
        ciphertext[50]), .Z(SubBytesIns_Inst_Sbox_6_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_6_T3), 
        .B(SubBytesIns_Inst_Sbox_6_T4), .Z(SubBytesIns_Inst_Sbox_6_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_6_T6), 
        .B(SubBytesIns_Inst_Sbox_6_T11), .Z(SubBytesIns_Inst_Sbox_6_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_6_T5), 
        .B(SubBytesIns_Inst_Sbox_6_T11), .Z(SubBytesIns_Inst_Sbox_6_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_6_T5), 
        .B(SubBytesIns_Inst_Sbox_6_T12), .Z(SubBytesIns_Inst_Sbox_6_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_6_T9), 
        .B(SubBytesIns_Inst_Sbox_6_T16), .Z(SubBytesIns_Inst_Sbox_6_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T18_U1 ( .A(ciphertext[52]), .B(
        ciphertext[48]), .Z(SubBytesIns_Inst_Sbox_6_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_6_T7), 
        .B(SubBytesIns_Inst_Sbox_6_T18), .Z(SubBytesIns_Inst_Sbox_6_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_6_T1), 
        .B(SubBytesIns_Inst_Sbox_6_T19), .Z(SubBytesIns_Inst_Sbox_6_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T21_U1 ( .A(ciphertext[49]), .B(
        ciphertext[48]), .Z(SubBytesIns_Inst_Sbox_6_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_6_T7), 
        .B(SubBytesIns_Inst_Sbox_6_T21), .Z(SubBytesIns_Inst_Sbox_6_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_6_T2), 
        .B(SubBytesIns_Inst_Sbox_6_T22), .Z(SubBytesIns_Inst_Sbox_6_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_6_T2), 
        .B(SubBytesIns_Inst_Sbox_6_T10), .Z(SubBytesIns_Inst_Sbox_6_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_6_T20), 
        .B(SubBytesIns_Inst_Sbox_6_T17), .Z(SubBytesIns_Inst_Sbox_6_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_6_T3), 
        .B(SubBytesIns_Inst_Sbox_6_T16), .Z(SubBytesIns_Inst_Sbox_6_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_6_T1), 
        .B(SubBytesIns_Inst_Sbox_6_T12), .Z(SubBytesIns_Inst_Sbox_6_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T13), 
        .A2(SubBytesIns_Inst_Sbox_6_T6), .ZN(SubBytesIns_Inst_Sbox_6_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T23), 
        .A2(SubBytesIns_Inst_Sbox_6_T8), .ZN(SubBytesIns_Inst_Sbox_6_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_6_T14), 
        .B(SubBytesIns_Inst_Sbox_6_M1), .Z(SubBytesIns_Inst_Sbox_6_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T19), 
        .A2(ciphertext[48]), .ZN(SubBytesIns_Inst_Sbox_6_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_6_M4), 
        .B(SubBytesIns_Inst_Sbox_6_M1), .Z(SubBytesIns_Inst_Sbox_6_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T3), 
        .A2(SubBytesIns_Inst_Sbox_6_T16), .ZN(SubBytesIns_Inst_Sbox_6_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T22), 
        .A2(SubBytesIns_Inst_Sbox_6_T9), .ZN(SubBytesIns_Inst_Sbox_6_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_6_T26), 
        .B(SubBytesIns_Inst_Sbox_6_M6), .Z(SubBytesIns_Inst_Sbox_6_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T20), 
        .A2(SubBytesIns_Inst_Sbox_6_T17), .ZN(SubBytesIns_Inst_Sbox_6_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_6_M9), 
        .B(SubBytesIns_Inst_Sbox_6_M6), .Z(SubBytesIns_Inst_Sbox_6_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T1), 
        .A2(SubBytesIns_Inst_Sbox_6_T15), .ZN(SubBytesIns_Inst_Sbox_6_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T4), 
        .A2(SubBytesIns_Inst_Sbox_6_T27), .ZN(SubBytesIns_Inst_Sbox_6_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_6_M12), 
        .B(SubBytesIns_Inst_Sbox_6_M11), .Z(SubBytesIns_Inst_Sbox_6_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T2), 
        .A2(SubBytesIns_Inst_Sbox_6_T10), .ZN(SubBytesIns_Inst_Sbox_6_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_6_M14), 
        .B(SubBytesIns_Inst_Sbox_6_M11), .Z(SubBytesIns_Inst_Sbox_6_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_6_M3), 
        .B(SubBytesIns_Inst_Sbox_6_M2), .Z(SubBytesIns_Inst_Sbox_6_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_6_M5), 
        .B(SubBytesIns_Inst_Sbox_6_T24), .Z(SubBytesIns_Inst_Sbox_6_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_6_M8), 
        .B(SubBytesIns_Inst_Sbox_6_M7), .Z(SubBytesIns_Inst_Sbox_6_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_6_M10), 
        .B(SubBytesIns_Inst_Sbox_6_M15), .Z(SubBytesIns_Inst_Sbox_6_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_6_M16), 
        .B(SubBytesIns_Inst_Sbox_6_M13), .Z(SubBytesIns_Inst_Sbox_6_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_6_M17), 
        .B(SubBytesIns_Inst_Sbox_6_M15), .Z(SubBytesIns_Inst_Sbox_6_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_6_M18), 
        .B(SubBytesIns_Inst_Sbox_6_M13), .Z(SubBytesIns_Inst_Sbox_6_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_6_M19), 
        .B(SubBytesIns_Inst_Sbox_6_T25), .Z(SubBytesIns_Inst_Sbox_6_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_6_M22), 
        .B(SubBytesIns_Inst_Sbox_6_M23), .Z(SubBytesIns_Inst_Sbox_6_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M22), .A2(SubBytesIns_Inst_Sbox_6_M20), .ZN(SubBytesIns_Inst_Sbox_6_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_6_M21), 
        .B(SubBytesIns_Inst_Sbox_6_M25), .Z(SubBytesIns_Inst_Sbox_6_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_6_M20), 
        .B(SubBytesIns_Inst_Sbox_6_M21), .Z(SubBytesIns_Inst_Sbox_6_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_6_M23), 
        .B(SubBytesIns_Inst_Sbox_6_M25), .Z(SubBytesIns_Inst_Sbox_6_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M28), .A2(SubBytesIns_Inst_Sbox_6_M27), .ZN(SubBytesIns_Inst_Sbox_6_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M26), .A2(SubBytesIns_Inst_Sbox_6_M24), .ZN(SubBytesIns_Inst_Sbox_6_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M20), .A2(SubBytesIns_Inst_Sbox_6_M23), .ZN(SubBytesIns_Inst_Sbox_6_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M27), .A2(SubBytesIns_Inst_Sbox_6_M31), .ZN(SubBytesIns_Inst_Sbox_6_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_6_M27), 
        .B(SubBytesIns_Inst_Sbox_6_M25), .Z(SubBytesIns_Inst_Sbox_6_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M21), .A2(SubBytesIns_Inst_Sbox_6_M22), .ZN(SubBytesIns_Inst_Sbox_6_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M24), .A2(SubBytesIns_Inst_Sbox_6_M34), .ZN(SubBytesIns_Inst_Sbox_6_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_6_M24), 
        .B(SubBytesIns_Inst_Sbox_6_M25), .Z(SubBytesIns_Inst_Sbox_6_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_6_M21), 
        .B(SubBytesIns_Inst_Sbox_6_M29), .Z(SubBytesIns_Inst_Sbox_6_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_6_M32), 
        .B(SubBytesIns_Inst_Sbox_6_M33), .Z(SubBytesIns_Inst_Sbox_6_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_6_M23), 
        .B(SubBytesIns_Inst_Sbox_6_M30), .Z(SubBytesIns_Inst_Sbox_6_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_6_M35), 
        .B(SubBytesIns_Inst_Sbox_6_M36), .Z(SubBytesIns_Inst_Sbox_6_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_6_M38), 
        .B(SubBytesIns_Inst_Sbox_6_M40), .Z(SubBytesIns_Inst_Sbox_6_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_6_M37), 
        .B(SubBytesIns_Inst_Sbox_6_M39), .Z(SubBytesIns_Inst_Sbox_6_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_6_M37), 
        .B(SubBytesIns_Inst_Sbox_6_M38), .Z(SubBytesIns_Inst_Sbox_6_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_6_M39), 
        .B(SubBytesIns_Inst_Sbox_6_M40), .Z(SubBytesIns_Inst_Sbox_6_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_6_M42), 
        .B(SubBytesIns_Inst_Sbox_6_M41), .Z(SubBytesIns_Inst_Sbox_6_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M44), .A2(SubBytesIns_Inst_Sbox_6_T6), .ZN(SubBytesIns_Inst_Sbox_6_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M40), .A2(SubBytesIns_Inst_Sbox_6_T8), .ZN(SubBytesIns_Inst_Sbox_6_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M39), .A2(ciphertext[48]), .ZN(SubBytesIns_Inst_Sbox_6_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M43), .A2(SubBytesIns_Inst_Sbox_6_T16), .ZN(SubBytesIns_Inst_Sbox_6_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M38), .A2(SubBytesIns_Inst_Sbox_6_T9), .ZN(SubBytesIns_Inst_Sbox_6_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M37), .A2(SubBytesIns_Inst_Sbox_6_T17), .ZN(SubBytesIns_Inst_Sbox_6_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M42), .A2(SubBytesIns_Inst_Sbox_6_T15), .ZN(SubBytesIns_Inst_Sbox_6_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M45), .A2(SubBytesIns_Inst_Sbox_6_T27), .ZN(SubBytesIns_Inst_Sbox_6_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M41), .A2(SubBytesIns_Inst_Sbox_6_T10), .ZN(SubBytesIns_Inst_Sbox_6_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M44), .A2(SubBytesIns_Inst_Sbox_6_T13), .ZN(SubBytesIns_Inst_Sbox_6_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M40), .A2(SubBytesIns_Inst_Sbox_6_T23), .ZN(SubBytesIns_Inst_Sbox_6_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M39), .A2(SubBytesIns_Inst_Sbox_6_T19), .ZN(SubBytesIns_Inst_Sbox_6_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M43), .A2(SubBytesIns_Inst_Sbox_6_T3), .ZN(SubBytesIns_Inst_Sbox_6_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M38), .A2(SubBytesIns_Inst_Sbox_6_T22), .ZN(SubBytesIns_Inst_Sbox_6_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M37), .A2(SubBytesIns_Inst_Sbox_6_T20), .ZN(SubBytesIns_Inst_Sbox_6_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M42), .A2(SubBytesIns_Inst_Sbox_6_T1), .ZN(SubBytesIns_Inst_Sbox_6_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M45), .A2(SubBytesIns_Inst_Sbox_6_T4), .ZN(SubBytesIns_Inst_Sbox_6_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M41), .A2(SubBytesIns_Inst_Sbox_6_T2), .ZN(SubBytesIns_Inst_Sbox_6_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_6_M61), 
        .B(SubBytesIns_Inst_Sbox_6_M62), .Z(SubBytesIns_Inst_Sbox_6_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_6_M50), 
        .B(SubBytesIns_Inst_Sbox_6_M56), .Z(SubBytesIns_Inst_Sbox_6_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_6_M46), 
        .B(SubBytesIns_Inst_Sbox_6_M48), .Z(SubBytesIns_Inst_Sbox_6_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_6_M47), 
        .B(SubBytesIns_Inst_Sbox_6_M55), .Z(SubBytesIns_Inst_Sbox_6_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_6_M54), 
        .B(SubBytesIns_Inst_Sbox_6_M58), .Z(SubBytesIns_Inst_Sbox_6_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_6_M49), 
        .B(SubBytesIns_Inst_Sbox_6_M61), .Z(SubBytesIns_Inst_Sbox_6_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_6_M62), 
        .B(SubBytesIns_Inst_Sbox_6_L5), .Z(SubBytesIns_Inst_Sbox_6_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_6_M46), 
        .B(SubBytesIns_Inst_Sbox_6_L3), .Z(SubBytesIns_Inst_Sbox_6_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_6_M51), 
        .B(SubBytesIns_Inst_Sbox_6_M59), .Z(SubBytesIns_Inst_Sbox_6_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_6_M52), 
        .B(SubBytesIns_Inst_Sbox_6_M53), .Z(SubBytesIns_Inst_Sbox_6_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_6_M53), 
        .B(SubBytesIns_Inst_Sbox_6_L4), .Z(SubBytesIns_Inst_Sbox_6_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_6_M60), 
        .B(SubBytesIns_Inst_Sbox_6_L2), .Z(SubBytesIns_Inst_Sbox_6_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_6_M48), 
        .B(SubBytesIns_Inst_Sbox_6_M51), .Z(SubBytesIns_Inst_Sbox_6_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_6_M50), 
        .B(SubBytesIns_Inst_Sbox_6_L0), .Z(SubBytesIns_Inst_Sbox_6_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_6_M52), 
        .B(SubBytesIns_Inst_Sbox_6_M61), .Z(SubBytesIns_Inst_Sbox_6_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_6_M55), 
        .B(SubBytesIns_Inst_Sbox_6_L1), .Z(SubBytesIns_Inst_Sbox_6_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_6_M56), 
        .B(SubBytesIns_Inst_Sbox_6_L0), .Z(SubBytesIns_Inst_Sbox_6_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_6_M57), 
        .B(SubBytesIns_Inst_Sbox_6_L1), .Z(SubBytesIns_Inst_Sbox_6_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_6_M58), 
        .B(SubBytesIns_Inst_Sbox_6_L8), .Z(SubBytesIns_Inst_Sbox_6_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_6_M63), 
        .B(SubBytesIns_Inst_Sbox_6_L4), .Z(SubBytesIns_Inst_Sbox_6_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_6_L0), 
        .B(SubBytesIns_Inst_Sbox_6_L1), .Z(SubBytesIns_Inst_Sbox_6_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_6_L1), 
        .B(SubBytesIns_Inst_Sbox_6_L7), .Z(SubBytesIns_Inst_Sbox_6_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_6_L3), 
        .B(SubBytesIns_Inst_Sbox_6_L12), .Z(SubBytesIns_Inst_Sbox_6_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_6_L18), 
        .B(SubBytesIns_Inst_Sbox_6_L2), .Z(SubBytesIns_Inst_Sbox_6_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_6_L15), 
        .B(SubBytesIns_Inst_Sbox_6_L9), .Z(SubBytesIns_Inst_Sbox_6_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_6_L6), 
        .B(SubBytesIns_Inst_Sbox_6_L10), .Z(SubBytesIns_Inst_Sbox_6_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_6_L7), 
        .B(SubBytesIns_Inst_Sbox_6_L9), .Z(SubBytesIns_Inst_Sbox_6_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_6_L8), 
        .B(SubBytesIns_Inst_Sbox_6_L10), .Z(SubBytesIns_Inst_Sbox_6_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_6_L11), 
        .B(SubBytesIns_Inst_Sbox_6_L14), .Z(SubBytesIns_Inst_Sbox_6_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_6_L11), 
        .B(SubBytesIns_Inst_Sbox_6_L17), .Z(SubBytesIns_Inst_Sbox_6_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_6_L6), 
        .B(SubBytesIns_Inst_Sbox_6_L24), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_6_L16), 
        .B(SubBytesIns_Inst_Sbox_6_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_6_L19), 
        .B(SubBytesIns_Inst_Sbox_6_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_6_L6), 
        .B(SubBytesIns_Inst_Sbox_6_L21), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_6_L20), 
        .B(SubBytesIns_Inst_Sbox_6_L22), .Z(MixColumnsInput[83]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_6_L25), 
        .B(SubBytesIns_Inst_Sbox_6_L29), .Z(MixColumnsInput[82]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_6_L13), 
        .B(SubBytesIns_Inst_Sbox_6_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_6_L6), 
        .B(SubBytesIns_Inst_Sbox_6_L23), .ZN(MixColumnsInput[80]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T1_U1 ( .A(ciphertext[63]), .B(
        ciphertext[60]), .Z(SubBytesIns_Inst_Sbox_7_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T2_U1 ( .A(ciphertext[63]), .B(
        ciphertext[58]), .Z(SubBytesIns_Inst_Sbox_7_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T3_U1 ( .A(ciphertext[63]), .B(
        ciphertext[57]), .Z(SubBytesIns_Inst_Sbox_7_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T4_U1 ( .A(ciphertext[60]), .B(
        ciphertext[58]), .Z(SubBytesIns_Inst_Sbox_7_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T5_U1 ( .A(ciphertext[59]), .B(
        ciphertext[57]), .Z(SubBytesIns_Inst_Sbox_7_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_7_T1), 
        .B(SubBytesIns_Inst_Sbox_7_T5), .Z(SubBytesIns_Inst_Sbox_7_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T7_U1 ( .A(ciphertext[62]), .B(
        ciphertext[61]), .Z(SubBytesIns_Inst_Sbox_7_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T8_U1 ( .A(ciphertext[56]), .B(
        SubBytesIns_Inst_Sbox_7_T6), .Z(SubBytesIns_Inst_Sbox_7_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T9_U1 ( .A(ciphertext[56]), .B(
        SubBytesIns_Inst_Sbox_7_T7), .Z(SubBytesIns_Inst_Sbox_7_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_7_T6), 
        .B(SubBytesIns_Inst_Sbox_7_T7), .Z(SubBytesIns_Inst_Sbox_7_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T11_U1 ( .A(ciphertext[62]), .B(
        ciphertext[58]), .Z(SubBytesIns_Inst_Sbox_7_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T12_U1 ( .A(ciphertext[61]), .B(
        ciphertext[58]), .Z(SubBytesIns_Inst_Sbox_7_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_7_T3), 
        .B(SubBytesIns_Inst_Sbox_7_T4), .Z(SubBytesIns_Inst_Sbox_7_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_7_T6), 
        .B(SubBytesIns_Inst_Sbox_7_T11), .Z(SubBytesIns_Inst_Sbox_7_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_7_T5), 
        .B(SubBytesIns_Inst_Sbox_7_T11), .Z(SubBytesIns_Inst_Sbox_7_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_7_T5), 
        .B(SubBytesIns_Inst_Sbox_7_T12), .Z(SubBytesIns_Inst_Sbox_7_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_7_T9), 
        .B(SubBytesIns_Inst_Sbox_7_T16), .Z(SubBytesIns_Inst_Sbox_7_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T18_U1 ( .A(ciphertext[60]), .B(
        ciphertext[56]), .Z(SubBytesIns_Inst_Sbox_7_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_7_T7), 
        .B(SubBytesIns_Inst_Sbox_7_T18), .Z(SubBytesIns_Inst_Sbox_7_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_7_T1), 
        .B(SubBytesIns_Inst_Sbox_7_T19), .Z(SubBytesIns_Inst_Sbox_7_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T21_U1 ( .A(ciphertext[57]), .B(
        ciphertext[56]), .Z(SubBytesIns_Inst_Sbox_7_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_7_T7), 
        .B(SubBytesIns_Inst_Sbox_7_T21), .Z(SubBytesIns_Inst_Sbox_7_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_7_T2), 
        .B(SubBytesIns_Inst_Sbox_7_T22), .Z(SubBytesIns_Inst_Sbox_7_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_7_T2), 
        .B(SubBytesIns_Inst_Sbox_7_T10), .Z(SubBytesIns_Inst_Sbox_7_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_7_T20), 
        .B(SubBytesIns_Inst_Sbox_7_T17), .Z(SubBytesIns_Inst_Sbox_7_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_7_T3), 
        .B(SubBytesIns_Inst_Sbox_7_T16), .Z(SubBytesIns_Inst_Sbox_7_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_7_T1), 
        .B(SubBytesIns_Inst_Sbox_7_T12), .Z(SubBytesIns_Inst_Sbox_7_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T13), 
        .A2(SubBytesIns_Inst_Sbox_7_T6), .ZN(SubBytesIns_Inst_Sbox_7_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T23), 
        .A2(SubBytesIns_Inst_Sbox_7_T8), .ZN(SubBytesIns_Inst_Sbox_7_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_7_T14), 
        .B(SubBytesIns_Inst_Sbox_7_M1), .Z(SubBytesIns_Inst_Sbox_7_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T19), 
        .A2(ciphertext[56]), .ZN(SubBytesIns_Inst_Sbox_7_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_7_M4), 
        .B(SubBytesIns_Inst_Sbox_7_M1), .Z(SubBytesIns_Inst_Sbox_7_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T3), 
        .A2(SubBytesIns_Inst_Sbox_7_T16), .ZN(SubBytesIns_Inst_Sbox_7_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T22), 
        .A2(SubBytesIns_Inst_Sbox_7_T9), .ZN(SubBytesIns_Inst_Sbox_7_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_7_T26), 
        .B(SubBytesIns_Inst_Sbox_7_M6), .Z(SubBytesIns_Inst_Sbox_7_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T20), 
        .A2(SubBytesIns_Inst_Sbox_7_T17), .ZN(SubBytesIns_Inst_Sbox_7_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_7_M9), 
        .B(SubBytesIns_Inst_Sbox_7_M6), .Z(SubBytesIns_Inst_Sbox_7_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T1), 
        .A2(SubBytesIns_Inst_Sbox_7_T15), .ZN(SubBytesIns_Inst_Sbox_7_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T4), 
        .A2(SubBytesIns_Inst_Sbox_7_T27), .ZN(SubBytesIns_Inst_Sbox_7_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_7_M12), 
        .B(SubBytesIns_Inst_Sbox_7_M11), .Z(SubBytesIns_Inst_Sbox_7_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T2), 
        .A2(SubBytesIns_Inst_Sbox_7_T10), .ZN(SubBytesIns_Inst_Sbox_7_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_7_M14), 
        .B(SubBytesIns_Inst_Sbox_7_M11), .Z(SubBytesIns_Inst_Sbox_7_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_7_M3), 
        .B(SubBytesIns_Inst_Sbox_7_M2), .Z(SubBytesIns_Inst_Sbox_7_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_7_M5), 
        .B(SubBytesIns_Inst_Sbox_7_T24), .Z(SubBytesIns_Inst_Sbox_7_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_7_M8), 
        .B(SubBytesIns_Inst_Sbox_7_M7), .Z(SubBytesIns_Inst_Sbox_7_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_7_M10), 
        .B(SubBytesIns_Inst_Sbox_7_M15), .Z(SubBytesIns_Inst_Sbox_7_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_7_M16), 
        .B(SubBytesIns_Inst_Sbox_7_M13), .Z(SubBytesIns_Inst_Sbox_7_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_7_M17), 
        .B(SubBytesIns_Inst_Sbox_7_M15), .Z(SubBytesIns_Inst_Sbox_7_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_7_M18), 
        .B(SubBytesIns_Inst_Sbox_7_M13), .Z(SubBytesIns_Inst_Sbox_7_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_7_M19), 
        .B(SubBytesIns_Inst_Sbox_7_T25), .Z(SubBytesIns_Inst_Sbox_7_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_7_M22), 
        .B(SubBytesIns_Inst_Sbox_7_M23), .Z(SubBytesIns_Inst_Sbox_7_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M22), .A2(SubBytesIns_Inst_Sbox_7_M20), .ZN(SubBytesIns_Inst_Sbox_7_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_7_M21), 
        .B(SubBytesIns_Inst_Sbox_7_M25), .Z(SubBytesIns_Inst_Sbox_7_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_7_M20), 
        .B(SubBytesIns_Inst_Sbox_7_M21), .Z(SubBytesIns_Inst_Sbox_7_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_7_M23), 
        .B(SubBytesIns_Inst_Sbox_7_M25), .Z(SubBytesIns_Inst_Sbox_7_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M28), .A2(SubBytesIns_Inst_Sbox_7_M27), .ZN(SubBytesIns_Inst_Sbox_7_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M26), .A2(SubBytesIns_Inst_Sbox_7_M24), .ZN(SubBytesIns_Inst_Sbox_7_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M20), .A2(SubBytesIns_Inst_Sbox_7_M23), .ZN(SubBytesIns_Inst_Sbox_7_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M27), .A2(SubBytesIns_Inst_Sbox_7_M31), .ZN(SubBytesIns_Inst_Sbox_7_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_7_M27), 
        .B(SubBytesIns_Inst_Sbox_7_M25), .Z(SubBytesIns_Inst_Sbox_7_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M21), .A2(SubBytesIns_Inst_Sbox_7_M22), .ZN(SubBytesIns_Inst_Sbox_7_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M24), .A2(SubBytesIns_Inst_Sbox_7_M34), .ZN(SubBytesIns_Inst_Sbox_7_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_7_M24), 
        .B(SubBytesIns_Inst_Sbox_7_M25), .Z(SubBytesIns_Inst_Sbox_7_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_7_M21), 
        .B(SubBytesIns_Inst_Sbox_7_M29), .Z(SubBytesIns_Inst_Sbox_7_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_7_M32), 
        .B(SubBytesIns_Inst_Sbox_7_M33), .Z(SubBytesIns_Inst_Sbox_7_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_7_M23), 
        .B(SubBytesIns_Inst_Sbox_7_M30), .Z(SubBytesIns_Inst_Sbox_7_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_7_M35), 
        .B(SubBytesIns_Inst_Sbox_7_M36), .Z(SubBytesIns_Inst_Sbox_7_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_7_M38), 
        .B(SubBytesIns_Inst_Sbox_7_M40), .Z(SubBytesIns_Inst_Sbox_7_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_7_M37), 
        .B(SubBytesIns_Inst_Sbox_7_M39), .Z(SubBytesIns_Inst_Sbox_7_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_7_M37), 
        .B(SubBytesIns_Inst_Sbox_7_M38), .Z(SubBytesIns_Inst_Sbox_7_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_7_M39), 
        .B(SubBytesIns_Inst_Sbox_7_M40), .Z(SubBytesIns_Inst_Sbox_7_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_7_M42), 
        .B(SubBytesIns_Inst_Sbox_7_M41), .Z(SubBytesIns_Inst_Sbox_7_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M44), .A2(SubBytesIns_Inst_Sbox_7_T6), .ZN(SubBytesIns_Inst_Sbox_7_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M40), .A2(SubBytesIns_Inst_Sbox_7_T8), .ZN(SubBytesIns_Inst_Sbox_7_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M39), .A2(ciphertext[56]), .ZN(SubBytesIns_Inst_Sbox_7_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M43), .A2(SubBytesIns_Inst_Sbox_7_T16), .ZN(SubBytesIns_Inst_Sbox_7_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M38), .A2(SubBytesIns_Inst_Sbox_7_T9), .ZN(SubBytesIns_Inst_Sbox_7_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M37), .A2(SubBytesIns_Inst_Sbox_7_T17), .ZN(SubBytesIns_Inst_Sbox_7_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M42), .A2(SubBytesIns_Inst_Sbox_7_T15), .ZN(SubBytesIns_Inst_Sbox_7_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M45), .A2(SubBytesIns_Inst_Sbox_7_T27), .ZN(SubBytesIns_Inst_Sbox_7_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M41), .A2(SubBytesIns_Inst_Sbox_7_T10), .ZN(SubBytesIns_Inst_Sbox_7_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M44), .A2(SubBytesIns_Inst_Sbox_7_T13), .ZN(SubBytesIns_Inst_Sbox_7_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M40), .A2(SubBytesIns_Inst_Sbox_7_T23), .ZN(SubBytesIns_Inst_Sbox_7_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M39), .A2(SubBytesIns_Inst_Sbox_7_T19), .ZN(SubBytesIns_Inst_Sbox_7_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M43), .A2(SubBytesIns_Inst_Sbox_7_T3), .ZN(SubBytesIns_Inst_Sbox_7_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M38), .A2(SubBytesIns_Inst_Sbox_7_T22), .ZN(SubBytesIns_Inst_Sbox_7_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M37), .A2(SubBytesIns_Inst_Sbox_7_T20), .ZN(SubBytesIns_Inst_Sbox_7_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M42), .A2(SubBytesIns_Inst_Sbox_7_T1), .ZN(SubBytesIns_Inst_Sbox_7_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M45), .A2(SubBytesIns_Inst_Sbox_7_T4), .ZN(SubBytesIns_Inst_Sbox_7_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M41), .A2(SubBytesIns_Inst_Sbox_7_T2), .ZN(SubBytesIns_Inst_Sbox_7_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_7_M61), 
        .B(SubBytesIns_Inst_Sbox_7_M62), .Z(SubBytesIns_Inst_Sbox_7_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_7_M50), 
        .B(SubBytesIns_Inst_Sbox_7_M56), .Z(SubBytesIns_Inst_Sbox_7_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_7_M46), 
        .B(SubBytesIns_Inst_Sbox_7_M48), .Z(SubBytesIns_Inst_Sbox_7_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_7_M47), 
        .B(SubBytesIns_Inst_Sbox_7_M55), .Z(SubBytesIns_Inst_Sbox_7_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_7_M54), 
        .B(SubBytesIns_Inst_Sbox_7_M58), .Z(SubBytesIns_Inst_Sbox_7_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_7_M49), 
        .B(SubBytesIns_Inst_Sbox_7_M61), .Z(SubBytesIns_Inst_Sbox_7_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_7_M62), 
        .B(SubBytesIns_Inst_Sbox_7_L5), .Z(SubBytesIns_Inst_Sbox_7_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_7_M46), 
        .B(SubBytesIns_Inst_Sbox_7_L3), .Z(SubBytesIns_Inst_Sbox_7_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_7_M51), 
        .B(SubBytesIns_Inst_Sbox_7_M59), .Z(SubBytesIns_Inst_Sbox_7_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_7_M52), 
        .B(SubBytesIns_Inst_Sbox_7_M53), .Z(SubBytesIns_Inst_Sbox_7_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_7_M53), 
        .B(SubBytesIns_Inst_Sbox_7_L4), .Z(SubBytesIns_Inst_Sbox_7_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_7_M60), 
        .B(SubBytesIns_Inst_Sbox_7_L2), .Z(SubBytesIns_Inst_Sbox_7_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_7_M48), 
        .B(SubBytesIns_Inst_Sbox_7_M51), .Z(SubBytesIns_Inst_Sbox_7_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_7_M50), 
        .B(SubBytesIns_Inst_Sbox_7_L0), .Z(SubBytesIns_Inst_Sbox_7_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_7_M52), 
        .B(SubBytesIns_Inst_Sbox_7_M61), .Z(SubBytesIns_Inst_Sbox_7_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_7_M55), 
        .B(SubBytesIns_Inst_Sbox_7_L1), .Z(SubBytesIns_Inst_Sbox_7_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_7_M56), 
        .B(SubBytesIns_Inst_Sbox_7_L0), .Z(SubBytesIns_Inst_Sbox_7_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_7_M57), 
        .B(SubBytesIns_Inst_Sbox_7_L1), .Z(SubBytesIns_Inst_Sbox_7_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_7_M58), 
        .B(SubBytesIns_Inst_Sbox_7_L8), .Z(SubBytesIns_Inst_Sbox_7_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_7_M63), 
        .B(SubBytesIns_Inst_Sbox_7_L4), .Z(SubBytesIns_Inst_Sbox_7_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_7_L0), 
        .B(SubBytesIns_Inst_Sbox_7_L1), .Z(SubBytesIns_Inst_Sbox_7_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_7_L1), 
        .B(SubBytesIns_Inst_Sbox_7_L7), .Z(SubBytesIns_Inst_Sbox_7_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_7_L3), 
        .B(SubBytesIns_Inst_Sbox_7_L12), .Z(SubBytesIns_Inst_Sbox_7_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_7_L18), 
        .B(SubBytesIns_Inst_Sbox_7_L2), .Z(SubBytesIns_Inst_Sbox_7_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_7_L15), 
        .B(SubBytesIns_Inst_Sbox_7_L9), .Z(SubBytesIns_Inst_Sbox_7_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_7_L6), 
        .B(SubBytesIns_Inst_Sbox_7_L10), .Z(SubBytesIns_Inst_Sbox_7_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_7_L7), 
        .B(SubBytesIns_Inst_Sbox_7_L9), .Z(SubBytesIns_Inst_Sbox_7_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_7_L8), 
        .B(SubBytesIns_Inst_Sbox_7_L10), .Z(SubBytesIns_Inst_Sbox_7_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_7_L11), 
        .B(SubBytesIns_Inst_Sbox_7_L14), .Z(SubBytesIns_Inst_Sbox_7_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_7_L11), 
        .B(SubBytesIns_Inst_Sbox_7_L17), .Z(SubBytesIns_Inst_Sbox_7_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_7_L6), 
        .B(SubBytesIns_Inst_Sbox_7_L24), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_7_L16), 
        .B(SubBytesIns_Inst_Sbox_7_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_7_L19), 
        .B(SubBytesIns_Inst_Sbox_7_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_7_L6), 
        .B(SubBytesIns_Inst_Sbox_7_L21), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_7_L20), 
        .B(SubBytesIns_Inst_Sbox_7_L22), .Z(MixColumnsInput[59]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_7_L25), 
        .B(SubBytesIns_Inst_Sbox_7_L29), .Z(MixColumnsInput[58]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_7_L13), 
        .B(SubBytesIns_Inst_Sbox_7_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_7_L6), 
        .B(SubBytesIns_Inst_Sbox_7_L23), .ZN(MixColumnsInput[56]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T1_U1 ( .A(ciphertext[71]), .B(
        ciphertext[68]), .Z(SubBytesIns_Inst_Sbox_8_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T2_U1 ( .A(ciphertext[71]), .B(
        ciphertext[66]), .Z(SubBytesIns_Inst_Sbox_8_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T3_U1 ( .A(ciphertext[71]), .B(
        ciphertext[65]), .Z(SubBytesIns_Inst_Sbox_8_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T4_U1 ( .A(ciphertext[68]), .B(
        ciphertext[66]), .Z(SubBytesIns_Inst_Sbox_8_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T5_U1 ( .A(ciphertext[67]), .B(
        ciphertext[65]), .Z(SubBytesIns_Inst_Sbox_8_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_8_T1), 
        .B(SubBytesIns_Inst_Sbox_8_T5), .Z(SubBytesIns_Inst_Sbox_8_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T7_U1 ( .A(ciphertext[70]), .B(
        ciphertext[69]), .Z(SubBytesIns_Inst_Sbox_8_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T8_U1 ( .A(ciphertext[64]), .B(
        SubBytesIns_Inst_Sbox_8_T6), .Z(SubBytesIns_Inst_Sbox_8_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T9_U1 ( .A(ciphertext[64]), .B(
        SubBytesIns_Inst_Sbox_8_T7), .Z(SubBytesIns_Inst_Sbox_8_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_8_T6), 
        .B(SubBytesIns_Inst_Sbox_8_T7), .Z(SubBytesIns_Inst_Sbox_8_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T11_U1 ( .A(ciphertext[70]), .B(
        ciphertext[66]), .Z(SubBytesIns_Inst_Sbox_8_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T12_U1 ( .A(ciphertext[69]), .B(
        ciphertext[66]), .Z(SubBytesIns_Inst_Sbox_8_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_8_T3), 
        .B(SubBytesIns_Inst_Sbox_8_T4), .Z(SubBytesIns_Inst_Sbox_8_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_8_T6), 
        .B(SubBytesIns_Inst_Sbox_8_T11), .Z(SubBytesIns_Inst_Sbox_8_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_8_T5), 
        .B(SubBytesIns_Inst_Sbox_8_T11), .Z(SubBytesIns_Inst_Sbox_8_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_8_T5), 
        .B(SubBytesIns_Inst_Sbox_8_T12), .Z(SubBytesIns_Inst_Sbox_8_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_8_T9), 
        .B(SubBytesIns_Inst_Sbox_8_T16), .Z(SubBytesIns_Inst_Sbox_8_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T18_U1 ( .A(ciphertext[68]), .B(
        ciphertext[64]), .Z(SubBytesIns_Inst_Sbox_8_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_8_T7), 
        .B(SubBytesIns_Inst_Sbox_8_T18), .Z(SubBytesIns_Inst_Sbox_8_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_8_T1), 
        .B(SubBytesIns_Inst_Sbox_8_T19), .Z(SubBytesIns_Inst_Sbox_8_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T21_U1 ( .A(ciphertext[65]), .B(
        ciphertext[64]), .Z(SubBytesIns_Inst_Sbox_8_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_8_T7), 
        .B(SubBytesIns_Inst_Sbox_8_T21), .Z(SubBytesIns_Inst_Sbox_8_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_8_T2), 
        .B(SubBytesIns_Inst_Sbox_8_T22), .Z(SubBytesIns_Inst_Sbox_8_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_8_T2), 
        .B(SubBytesIns_Inst_Sbox_8_T10), .Z(SubBytesIns_Inst_Sbox_8_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_8_T20), 
        .B(SubBytesIns_Inst_Sbox_8_T17), .Z(SubBytesIns_Inst_Sbox_8_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_8_T3), 
        .B(SubBytesIns_Inst_Sbox_8_T16), .Z(SubBytesIns_Inst_Sbox_8_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_8_T1), 
        .B(SubBytesIns_Inst_Sbox_8_T12), .Z(SubBytesIns_Inst_Sbox_8_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T13), 
        .A2(SubBytesIns_Inst_Sbox_8_T6), .ZN(SubBytesIns_Inst_Sbox_8_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T23), 
        .A2(SubBytesIns_Inst_Sbox_8_T8), .ZN(SubBytesIns_Inst_Sbox_8_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_8_T14), 
        .B(SubBytesIns_Inst_Sbox_8_M1), .Z(SubBytesIns_Inst_Sbox_8_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T19), 
        .A2(ciphertext[64]), .ZN(SubBytesIns_Inst_Sbox_8_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_8_M4), 
        .B(SubBytesIns_Inst_Sbox_8_M1), .Z(SubBytesIns_Inst_Sbox_8_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T3), 
        .A2(SubBytesIns_Inst_Sbox_8_T16), .ZN(SubBytesIns_Inst_Sbox_8_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T22), 
        .A2(SubBytesIns_Inst_Sbox_8_T9), .ZN(SubBytesIns_Inst_Sbox_8_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_8_T26), 
        .B(SubBytesIns_Inst_Sbox_8_M6), .Z(SubBytesIns_Inst_Sbox_8_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T20), 
        .A2(SubBytesIns_Inst_Sbox_8_T17), .ZN(SubBytesIns_Inst_Sbox_8_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_8_M9), 
        .B(SubBytesIns_Inst_Sbox_8_M6), .Z(SubBytesIns_Inst_Sbox_8_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T1), 
        .A2(SubBytesIns_Inst_Sbox_8_T15), .ZN(SubBytesIns_Inst_Sbox_8_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T4), 
        .A2(SubBytesIns_Inst_Sbox_8_T27), .ZN(SubBytesIns_Inst_Sbox_8_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_8_M12), 
        .B(SubBytesIns_Inst_Sbox_8_M11), .Z(SubBytesIns_Inst_Sbox_8_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T2), 
        .A2(SubBytesIns_Inst_Sbox_8_T10), .ZN(SubBytesIns_Inst_Sbox_8_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_8_M14), 
        .B(SubBytesIns_Inst_Sbox_8_M11), .Z(SubBytesIns_Inst_Sbox_8_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_8_M3), 
        .B(SubBytesIns_Inst_Sbox_8_M2), .Z(SubBytesIns_Inst_Sbox_8_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_8_M5), 
        .B(SubBytesIns_Inst_Sbox_8_T24), .Z(SubBytesIns_Inst_Sbox_8_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_8_M8), 
        .B(SubBytesIns_Inst_Sbox_8_M7), .Z(SubBytesIns_Inst_Sbox_8_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_8_M10), 
        .B(SubBytesIns_Inst_Sbox_8_M15), .Z(SubBytesIns_Inst_Sbox_8_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_8_M16), 
        .B(SubBytesIns_Inst_Sbox_8_M13), .Z(SubBytesIns_Inst_Sbox_8_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_8_M17), 
        .B(SubBytesIns_Inst_Sbox_8_M15), .Z(SubBytesIns_Inst_Sbox_8_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_8_M18), 
        .B(SubBytesIns_Inst_Sbox_8_M13), .Z(SubBytesIns_Inst_Sbox_8_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_8_M19), 
        .B(SubBytesIns_Inst_Sbox_8_T25), .Z(SubBytesIns_Inst_Sbox_8_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_8_M22), 
        .B(SubBytesIns_Inst_Sbox_8_M23), .Z(SubBytesIns_Inst_Sbox_8_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M22), .A2(SubBytesIns_Inst_Sbox_8_M20), .ZN(SubBytesIns_Inst_Sbox_8_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_8_M21), 
        .B(SubBytesIns_Inst_Sbox_8_M25), .Z(SubBytesIns_Inst_Sbox_8_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_8_M20), 
        .B(SubBytesIns_Inst_Sbox_8_M21), .Z(SubBytesIns_Inst_Sbox_8_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_8_M23), 
        .B(SubBytesIns_Inst_Sbox_8_M25), .Z(SubBytesIns_Inst_Sbox_8_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M28), .A2(SubBytesIns_Inst_Sbox_8_M27), .ZN(SubBytesIns_Inst_Sbox_8_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M26), .A2(SubBytesIns_Inst_Sbox_8_M24), .ZN(SubBytesIns_Inst_Sbox_8_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M20), .A2(SubBytesIns_Inst_Sbox_8_M23), .ZN(SubBytesIns_Inst_Sbox_8_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M27), .A2(SubBytesIns_Inst_Sbox_8_M31), .ZN(SubBytesIns_Inst_Sbox_8_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_8_M27), 
        .B(SubBytesIns_Inst_Sbox_8_M25), .Z(SubBytesIns_Inst_Sbox_8_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M21), .A2(SubBytesIns_Inst_Sbox_8_M22), .ZN(SubBytesIns_Inst_Sbox_8_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M24), .A2(SubBytesIns_Inst_Sbox_8_M34), .ZN(SubBytesIns_Inst_Sbox_8_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_8_M24), 
        .B(SubBytesIns_Inst_Sbox_8_M25), .Z(SubBytesIns_Inst_Sbox_8_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_8_M21), 
        .B(SubBytesIns_Inst_Sbox_8_M29), .Z(SubBytesIns_Inst_Sbox_8_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_8_M32), 
        .B(SubBytesIns_Inst_Sbox_8_M33), .Z(SubBytesIns_Inst_Sbox_8_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_8_M23), 
        .B(SubBytesIns_Inst_Sbox_8_M30), .Z(SubBytesIns_Inst_Sbox_8_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_8_M35), 
        .B(SubBytesIns_Inst_Sbox_8_M36), .Z(SubBytesIns_Inst_Sbox_8_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_8_M38), 
        .B(SubBytesIns_Inst_Sbox_8_M40), .Z(SubBytesIns_Inst_Sbox_8_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_8_M37), 
        .B(SubBytesIns_Inst_Sbox_8_M39), .Z(SubBytesIns_Inst_Sbox_8_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_8_M37), 
        .B(SubBytesIns_Inst_Sbox_8_M38), .Z(SubBytesIns_Inst_Sbox_8_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_8_M39), 
        .B(SubBytesIns_Inst_Sbox_8_M40), .Z(SubBytesIns_Inst_Sbox_8_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_8_M42), 
        .B(SubBytesIns_Inst_Sbox_8_M41), .Z(SubBytesIns_Inst_Sbox_8_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M44), .A2(SubBytesIns_Inst_Sbox_8_T6), .ZN(SubBytesIns_Inst_Sbox_8_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M40), .A2(SubBytesIns_Inst_Sbox_8_T8), .ZN(SubBytesIns_Inst_Sbox_8_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M39), .A2(ciphertext[64]), .ZN(SubBytesIns_Inst_Sbox_8_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M43), .A2(SubBytesIns_Inst_Sbox_8_T16), .ZN(SubBytesIns_Inst_Sbox_8_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M38), .A2(SubBytesIns_Inst_Sbox_8_T9), .ZN(SubBytesIns_Inst_Sbox_8_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M37), .A2(SubBytesIns_Inst_Sbox_8_T17), .ZN(SubBytesIns_Inst_Sbox_8_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M42), .A2(SubBytesIns_Inst_Sbox_8_T15), .ZN(SubBytesIns_Inst_Sbox_8_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M45), .A2(SubBytesIns_Inst_Sbox_8_T27), .ZN(SubBytesIns_Inst_Sbox_8_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M41), .A2(SubBytesIns_Inst_Sbox_8_T10), .ZN(SubBytesIns_Inst_Sbox_8_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M44), .A2(SubBytesIns_Inst_Sbox_8_T13), .ZN(SubBytesIns_Inst_Sbox_8_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M40), .A2(SubBytesIns_Inst_Sbox_8_T23), .ZN(SubBytesIns_Inst_Sbox_8_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M39), .A2(SubBytesIns_Inst_Sbox_8_T19), .ZN(SubBytesIns_Inst_Sbox_8_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M43), .A2(SubBytesIns_Inst_Sbox_8_T3), .ZN(SubBytesIns_Inst_Sbox_8_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M38), .A2(SubBytesIns_Inst_Sbox_8_T22), .ZN(SubBytesIns_Inst_Sbox_8_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M37), .A2(SubBytesIns_Inst_Sbox_8_T20), .ZN(SubBytesIns_Inst_Sbox_8_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M42), .A2(SubBytesIns_Inst_Sbox_8_T1), .ZN(SubBytesIns_Inst_Sbox_8_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M45), .A2(SubBytesIns_Inst_Sbox_8_T4), .ZN(SubBytesIns_Inst_Sbox_8_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M41), .A2(SubBytesIns_Inst_Sbox_8_T2), .ZN(SubBytesIns_Inst_Sbox_8_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_8_M61), 
        .B(SubBytesIns_Inst_Sbox_8_M62), .Z(SubBytesIns_Inst_Sbox_8_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_8_M50), 
        .B(SubBytesIns_Inst_Sbox_8_M56), .Z(SubBytesIns_Inst_Sbox_8_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_8_M46), 
        .B(SubBytesIns_Inst_Sbox_8_M48), .Z(SubBytesIns_Inst_Sbox_8_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_8_M47), 
        .B(SubBytesIns_Inst_Sbox_8_M55), .Z(SubBytesIns_Inst_Sbox_8_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_8_M54), 
        .B(SubBytesIns_Inst_Sbox_8_M58), .Z(SubBytesIns_Inst_Sbox_8_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_8_M49), 
        .B(SubBytesIns_Inst_Sbox_8_M61), .Z(SubBytesIns_Inst_Sbox_8_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_8_M62), 
        .B(SubBytesIns_Inst_Sbox_8_L5), .Z(SubBytesIns_Inst_Sbox_8_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_8_M46), 
        .B(SubBytesIns_Inst_Sbox_8_L3), .Z(SubBytesIns_Inst_Sbox_8_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_8_M51), 
        .B(SubBytesIns_Inst_Sbox_8_M59), .Z(SubBytesIns_Inst_Sbox_8_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_8_M52), 
        .B(SubBytesIns_Inst_Sbox_8_M53), .Z(SubBytesIns_Inst_Sbox_8_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_8_M53), 
        .B(SubBytesIns_Inst_Sbox_8_L4), .Z(SubBytesIns_Inst_Sbox_8_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_8_M60), 
        .B(SubBytesIns_Inst_Sbox_8_L2), .Z(SubBytesIns_Inst_Sbox_8_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_8_M48), 
        .B(SubBytesIns_Inst_Sbox_8_M51), .Z(SubBytesIns_Inst_Sbox_8_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_8_M50), 
        .B(SubBytesIns_Inst_Sbox_8_L0), .Z(SubBytesIns_Inst_Sbox_8_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_8_M52), 
        .B(SubBytesIns_Inst_Sbox_8_M61), .Z(SubBytesIns_Inst_Sbox_8_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_8_M55), 
        .B(SubBytesIns_Inst_Sbox_8_L1), .Z(SubBytesIns_Inst_Sbox_8_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_8_M56), 
        .B(SubBytesIns_Inst_Sbox_8_L0), .Z(SubBytesIns_Inst_Sbox_8_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_8_M57), 
        .B(SubBytesIns_Inst_Sbox_8_L1), .Z(SubBytesIns_Inst_Sbox_8_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_8_M58), 
        .B(SubBytesIns_Inst_Sbox_8_L8), .Z(SubBytesIns_Inst_Sbox_8_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_8_M63), 
        .B(SubBytesIns_Inst_Sbox_8_L4), .Z(SubBytesIns_Inst_Sbox_8_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_8_L0), 
        .B(SubBytesIns_Inst_Sbox_8_L1), .Z(SubBytesIns_Inst_Sbox_8_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_8_L1), 
        .B(SubBytesIns_Inst_Sbox_8_L7), .Z(SubBytesIns_Inst_Sbox_8_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_8_L3), 
        .B(SubBytesIns_Inst_Sbox_8_L12), .Z(SubBytesIns_Inst_Sbox_8_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_8_L18), 
        .B(SubBytesIns_Inst_Sbox_8_L2), .Z(SubBytesIns_Inst_Sbox_8_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_8_L15), 
        .B(SubBytesIns_Inst_Sbox_8_L9), .Z(SubBytesIns_Inst_Sbox_8_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_8_L6), 
        .B(SubBytesIns_Inst_Sbox_8_L10), .Z(SubBytesIns_Inst_Sbox_8_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_8_L7), 
        .B(SubBytesIns_Inst_Sbox_8_L9), .Z(SubBytesIns_Inst_Sbox_8_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_8_L8), 
        .B(SubBytesIns_Inst_Sbox_8_L10), .Z(SubBytesIns_Inst_Sbox_8_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_8_L11), 
        .B(SubBytesIns_Inst_Sbox_8_L14), .Z(SubBytesIns_Inst_Sbox_8_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_8_L11), 
        .B(SubBytesIns_Inst_Sbox_8_L17), .Z(SubBytesIns_Inst_Sbox_8_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_8_L6), 
        .B(SubBytesIns_Inst_Sbox_8_L24), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_8_L16), 
        .B(SubBytesIns_Inst_Sbox_8_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_8_L19), 
        .B(SubBytesIns_Inst_Sbox_8_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_8_L6), 
        .B(SubBytesIns_Inst_Sbox_8_L21), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_8_L20), 
        .B(SubBytesIns_Inst_Sbox_8_L22), .Z(MixColumnsInput[35]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_8_L25), 
        .B(SubBytesIns_Inst_Sbox_8_L29), .Z(MixColumnsInput[34]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_8_L13), 
        .B(SubBytesIns_Inst_Sbox_8_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_8_L6), 
        .B(SubBytesIns_Inst_Sbox_8_L23), .ZN(MixColumnsInput[32]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T1_U1 ( .A(ciphertext[79]), .B(
        ciphertext[76]), .Z(SubBytesIns_Inst_Sbox_9_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T2_U1 ( .A(ciphertext[79]), .B(
        ciphertext[74]), .Z(SubBytesIns_Inst_Sbox_9_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T3_U1 ( .A(ciphertext[79]), .B(
        ciphertext[73]), .Z(SubBytesIns_Inst_Sbox_9_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T4_U1 ( .A(ciphertext[76]), .B(
        ciphertext[74]), .Z(SubBytesIns_Inst_Sbox_9_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T5_U1 ( .A(ciphertext[75]), .B(
        ciphertext[73]), .Z(SubBytesIns_Inst_Sbox_9_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_9_T1), 
        .B(SubBytesIns_Inst_Sbox_9_T5), .Z(SubBytesIns_Inst_Sbox_9_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T7_U1 ( .A(ciphertext[78]), .B(
        ciphertext[77]), .Z(SubBytesIns_Inst_Sbox_9_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T8_U1 ( .A(ciphertext[72]), .B(
        SubBytesIns_Inst_Sbox_9_T6), .Z(SubBytesIns_Inst_Sbox_9_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T9_U1 ( .A(ciphertext[72]), .B(
        SubBytesIns_Inst_Sbox_9_T7), .Z(SubBytesIns_Inst_Sbox_9_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_9_T6), 
        .B(SubBytesIns_Inst_Sbox_9_T7), .Z(SubBytesIns_Inst_Sbox_9_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T11_U1 ( .A(ciphertext[78]), .B(
        ciphertext[74]), .Z(SubBytesIns_Inst_Sbox_9_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T12_U1 ( .A(ciphertext[77]), .B(
        ciphertext[74]), .Z(SubBytesIns_Inst_Sbox_9_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_9_T3), 
        .B(SubBytesIns_Inst_Sbox_9_T4), .Z(SubBytesIns_Inst_Sbox_9_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_9_T6), 
        .B(SubBytesIns_Inst_Sbox_9_T11), .Z(SubBytesIns_Inst_Sbox_9_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_9_T5), 
        .B(SubBytesIns_Inst_Sbox_9_T11), .Z(SubBytesIns_Inst_Sbox_9_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_9_T5), 
        .B(SubBytesIns_Inst_Sbox_9_T12), .Z(SubBytesIns_Inst_Sbox_9_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_9_T9), 
        .B(SubBytesIns_Inst_Sbox_9_T16), .Z(SubBytesIns_Inst_Sbox_9_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T18_U1 ( .A(ciphertext[76]), .B(
        ciphertext[72]), .Z(SubBytesIns_Inst_Sbox_9_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_9_T7), 
        .B(SubBytesIns_Inst_Sbox_9_T18), .Z(SubBytesIns_Inst_Sbox_9_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_9_T1), 
        .B(SubBytesIns_Inst_Sbox_9_T19), .Z(SubBytesIns_Inst_Sbox_9_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T21_U1 ( .A(ciphertext[73]), .B(
        ciphertext[72]), .Z(SubBytesIns_Inst_Sbox_9_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_9_T7), 
        .B(SubBytesIns_Inst_Sbox_9_T21), .Z(SubBytesIns_Inst_Sbox_9_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_9_T2), 
        .B(SubBytesIns_Inst_Sbox_9_T22), .Z(SubBytesIns_Inst_Sbox_9_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_9_T2), 
        .B(SubBytesIns_Inst_Sbox_9_T10), .Z(SubBytesIns_Inst_Sbox_9_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_9_T20), 
        .B(SubBytesIns_Inst_Sbox_9_T17), .Z(SubBytesIns_Inst_Sbox_9_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_9_T3), 
        .B(SubBytesIns_Inst_Sbox_9_T16), .Z(SubBytesIns_Inst_Sbox_9_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_9_T1), 
        .B(SubBytesIns_Inst_Sbox_9_T12), .Z(SubBytesIns_Inst_Sbox_9_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T13), 
        .A2(SubBytesIns_Inst_Sbox_9_T6), .ZN(SubBytesIns_Inst_Sbox_9_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T23), 
        .A2(SubBytesIns_Inst_Sbox_9_T8), .ZN(SubBytesIns_Inst_Sbox_9_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_9_T14), 
        .B(SubBytesIns_Inst_Sbox_9_M1), .Z(SubBytesIns_Inst_Sbox_9_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T19), 
        .A2(ciphertext[72]), .ZN(SubBytesIns_Inst_Sbox_9_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_9_M4), 
        .B(SubBytesIns_Inst_Sbox_9_M1), .Z(SubBytesIns_Inst_Sbox_9_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T3), 
        .A2(SubBytesIns_Inst_Sbox_9_T16), .ZN(SubBytesIns_Inst_Sbox_9_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T22), 
        .A2(SubBytesIns_Inst_Sbox_9_T9), .ZN(SubBytesIns_Inst_Sbox_9_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_9_T26), 
        .B(SubBytesIns_Inst_Sbox_9_M6), .Z(SubBytesIns_Inst_Sbox_9_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T20), 
        .A2(SubBytesIns_Inst_Sbox_9_T17), .ZN(SubBytesIns_Inst_Sbox_9_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_9_M9), 
        .B(SubBytesIns_Inst_Sbox_9_M6), .Z(SubBytesIns_Inst_Sbox_9_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T1), 
        .A2(SubBytesIns_Inst_Sbox_9_T15), .ZN(SubBytesIns_Inst_Sbox_9_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T4), 
        .A2(SubBytesIns_Inst_Sbox_9_T27), .ZN(SubBytesIns_Inst_Sbox_9_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_9_M12), 
        .B(SubBytesIns_Inst_Sbox_9_M11), .Z(SubBytesIns_Inst_Sbox_9_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T2), 
        .A2(SubBytesIns_Inst_Sbox_9_T10), .ZN(SubBytesIns_Inst_Sbox_9_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_9_M14), 
        .B(SubBytesIns_Inst_Sbox_9_M11), .Z(SubBytesIns_Inst_Sbox_9_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_9_M3), 
        .B(SubBytesIns_Inst_Sbox_9_M2), .Z(SubBytesIns_Inst_Sbox_9_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_9_M5), 
        .B(SubBytesIns_Inst_Sbox_9_T24), .Z(SubBytesIns_Inst_Sbox_9_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_9_M8), 
        .B(SubBytesIns_Inst_Sbox_9_M7), .Z(SubBytesIns_Inst_Sbox_9_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_9_M10), 
        .B(SubBytesIns_Inst_Sbox_9_M15), .Z(SubBytesIns_Inst_Sbox_9_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_9_M16), 
        .B(SubBytesIns_Inst_Sbox_9_M13), .Z(SubBytesIns_Inst_Sbox_9_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_9_M17), 
        .B(SubBytesIns_Inst_Sbox_9_M15), .Z(SubBytesIns_Inst_Sbox_9_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_9_M18), 
        .B(SubBytesIns_Inst_Sbox_9_M13), .Z(SubBytesIns_Inst_Sbox_9_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_9_M19), 
        .B(SubBytesIns_Inst_Sbox_9_T25), .Z(SubBytesIns_Inst_Sbox_9_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_9_M22), 
        .B(SubBytesIns_Inst_Sbox_9_M23), .Z(SubBytesIns_Inst_Sbox_9_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M22), .A2(SubBytesIns_Inst_Sbox_9_M20), .ZN(SubBytesIns_Inst_Sbox_9_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_9_M21), 
        .B(SubBytesIns_Inst_Sbox_9_M25), .Z(SubBytesIns_Inst_Sbox_9_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_9_M20), 
        .B(SubBytesIns_Inst_Sbox_9_M21), .Z(SubBytesIns_Inst_Sbox_9_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_9_M23), 
        .B(SubBytesIns_Inst_Sbox_9_M25), .Z(SubBytesIns_Inst_Sbox_9_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M28), .A2(SubBytesIns_Inst_Sbox_9_M27), .ZN(SubBytesIns_Inst_Sbox_9_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M26), .A2(SubBytesIns_Inst_Sbox_9_M24), .ZN(SubBytesIns_Inst_Sbox_9_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M20), .A2(SubBytesIns_Inst_Sbox_9_M23), .ZN(SubBytesIns_Inst_Sbox_9_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M27), .A2(SubBytesIns_Inst_Sbox_9_M31), .ZN(SubBytesIns_Inst_Sbox_9_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_9_M27), 
        .B(SubBytesIns_Inst_Sbox_9_M25), .Z(SubBytesIns_Inst_Sbox_9_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M21), .A2(SubBytesIns_Inst_Sbox_9_M22), .ZN(SubBytesIns_Inst_Sbox_9_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M24), .A2(SubBytesIns_Inst_Sbox_9_M34), .ZN(SubBytesIns_Inst_Sbox_9_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_9_M24), 
        .B(SubBytesIns_Inst_Sbox_9_M25), .Z(SubBytesIns_Inst_Sbox_9_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_9_M21), 
        .B(SubBytesIns_Inst_Sbox_9_M29), .Z(SubBytesIns_Inst_Sbox_9_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_9_M32), 
        .B(SubBytesIns_Inst_Sbox_9_M33), .Z(SubBytesIns_Inst_Sbox_9_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_9_M23), 
        .B(SubBytesIns_Inst_Sbox_9_M30), .Z(SubBytesIns_Inst_Sbox_9_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_9_M35), 
        .B(SubBytesIns_Inst_Sbox_9_M36), .Z(SubBytesIns_Inst_Sbox_9_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_9_M38), 
        .B(SubBytesIns_Inst_Sbox_9_M40), .Z(SubBytesIns_Inst_Sbox_9_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_9_M37), 
        .B(SubBytesIns_Inst_Sbox_9_M39), .Z(SubBytesIns_Inst_Sbox_9_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_9_M37), 
        .B(SubBytesIns_Inst_Sbox_9_M38), .Z(SubBytesIns_Inst_Sbox_9_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_9_M39), 
        .B(SubBytesIns_Inst_Sbox_9_M40), .Z(SubBytesIns_Inst_Sbox_9_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_9_M42), 
        .B(SubBytesIns_Inst_Sbox_9_M41), .Z(SubBytesIns_Inst_Sbox_9_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M44), .A2(SubBytesIns_Inst_Sbox_9_T6), .ZN(SubBytesIns_Inst_Sbox_9_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M40), .A2(SubBytesIns_Inst_Sbox_9_T8), .ZN(SubBytesIns_Inst_Sbox_9_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M39), .A2(ciphertext[72]), .ZN(SubBytesIns_Inst_Sbox_9_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M43), .A2(SubBytesIns_Inst_Sbox_9_T16), .ZN(SubBytesIns_Inst_Sbox_9_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M38), .A2(SubBytesIns_Inst_Sbox_9_T9), .ZN(SubBytesIns_Inst_Sbox_9_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M37), .A2(SubBytesIns_Inst_Sbox_9_T17), .ZN(SubBytesIns_Inst_Sbox_9_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M42), .A2(SubBytesIns_Inst_Sbox_9_T15), .ZN(SubBytesIns_Inst_Sbox_9_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M45), .A2(SubBytesIns_Inst_Sbox_9_T27), .ZN(SubBytesIns_Inst_Sbox_9_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M41), .A2(SubBytesIns_Inst_Sbox_9_T10), .ZN(SubBytesIns_Inst_Sbox_9_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M44), .A2(SubBytesIns_Inst_Sbox_9_T13), .ZN(SubBytesIns_Inst_Sbox_9_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M40), .A2(SubBytesIns_Inst_Sbox_9_T23), .ZN(SubBytesIns_Inst_Sbox_9_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M39), .A2(SubBytesIns_Inst_Sbox_9_T19), .ZN(SubBytesIns_Inst_Sbox_9_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M43), .A2(SubBytesIns_Inst_Sbox_9_T3), .ZN(SubBytesIns_Inst_Sbox_9_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M38), .A2(SubBytesIns_Inst_Sbox_9_T22), .ZN(SubBytesIns_Inst_Sbox_9_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M37), .A2(SubBytesIns_Inst_Sbox_9_T20), .ZN(SubBytesIns_Inst_Sbox_9_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M42), .A2(SubBytesIns_Inst_Sbox_9_T1), .ZN(SubBytesIns_Inst_Sbox_9_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M45), .A2(SubBytesIns_Inst_Sbox_9_T4), .ZN(SubBytesIns_Inst_Sbox_9_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M41), .A2(SubBytesIns_Inst_Sbox_9_T2), .ZN(SubBytesIns_Inst_Sbox_9_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_9_M61), 
        .B(SubBytesIns_Inst_Sbox_9_M62), .Z(SubBytesIns_Inst_Sbox_9_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_9_M50), 
        .B(SubBytesIns_Inst_Sbox_9_M56), .Z(SubBytesIns_Inst_Sbox_9_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_9_M46), 
        .B(SubBytesIns_Inst_Sbox_9_M48), .Z(SubBytesIns_Inst_Sbox_9_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_9_M47), 
        .B(SubBytesIns_Inst_Sbox_9_M55), .Z(SubBytesIns_Inst_Sbox_9_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_9_M54), 
        .B(SubBytesIns_Inst_Sbox_9_M58), .Z(SubBytesIns_Inst_Sbox_9_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_9_M49), 
        .B(SubBytesIns_Inst_Sbox_9_M61), .Z(SubBytesIns_Inst_Sbox_9_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_9_M62), 
        .B(SubBytesIns_Inst_Sbox_9_L5), .Z(SubBytesIns_Inst_Sbox_9_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_9_M46), 
        .B(SubBytesIns_Inst_Sbox_9_L3), .Z(SubBytesIns_Inst_Sbox_9_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_9_M51), 
        .B(SubBytesIns_Inst_Sbox_9_M59), .Z(SubBytesIns_Inst_Sbox_9_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_9_M52), 
        .B(SubBytesIns_Inst_Sbox_9_M53), .Z(SubBytesIns_Inst_Sbox_9_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_9_M53), 
        .B(SubBytesIns_Inst_Sbox_9_L4), .Z(SubBytesIns_Inst_Sbox_9_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_9_M60), 
        .B(SubBytesIns_Inst_Sbox_9_L2), .Z(SubBytesIns_Inst_Sbox_9_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_9_M48), 
        .B(SubBytesIns_Inst_Sbox_9_M51), .Z(SubBytesIns_Inst_Sbox_9_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_9_M50), 
        .B(SubBytesIns_Inst_Sbox_9_L0), .Z(SubBytesIns_Inst_Sbox_9_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_9_M52), 
        .B(SubBytesIns_Inst_Sbox_9_M61), .Z(SubBytesIns_Inst_Sbox_9_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_9_M55), 
        .B(SubBytesIns_Inst_Sbox_9_L1), .Z(SubBytesIns_Inst_Sbox_9_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_9_M56), 
        .B(SubBytesIns_Inst_Sbox_9_L0), .Z(SubBytesIns_Inst_Sbox_9_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_9_M57), 
        .B(SubBytesIns_Inst_Sbox_9_L1), .Z(SubBytesIns_Inst_Sbox_9_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_9_M58), 
        .B(SubBytesIns_Inst_Sbox_9_L8), .Z(SubBytesIns_Inst_Sbox_9_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_9_M63), 
        .B(SubBytesIns_Inst_Sbox_9_L4), .Z(SubBytesIns_Inst_Sbox_9_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_9_L0), 
        .B(SubBytesIns_Inst_Sbox_9_L1), .Z(SubBytesIns_Inst_Sbox_9_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_9_L1), 
        .B(SubBytesIns_Inst_Sbox_9_L7), .Z(SubBytesIns_Inst_Sbox_9_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_9_L3), 
        .B(SubBytesIns_Inst_Sbox_9_L12), .Z(SubBytesIns_Inst_Sbox_9_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_9_L18), 
        .B(SubBytesIns_Inst_Sbox_9_L2), .Z(SubBytesIns_Inst_Sbox_9_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_9_L15), 
        .B(SubBytesIns_Inst_Sbox_9_L9), .Z(SubBytesIns_Inst_Sbox_9_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_9_L6), 
        .B(SubBytesIns_Inst_Sbox_9_L10), .Z(SubBytesIns_Inst_Sbox_9_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_9_L7), 
        .B(SubBytesIns_Inst_Sbox_9_L9), .Z(SubBytesIns_Inst_Sbox_9_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_9_L8), 
        .B(SubBytesIns_Inst_Sbox_9_L10), .Z(SubBytesIns_Inst_Sbox_9_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_9_L11), 
        .B(SubBytesIns_Inst_Sbox_9_L14), .Z(SubBytesIns_Inst_Sbox_9_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_9_L11), 
        .B(SubBytesIns_Inst_Sbox_9_L17), .Z(SubBytesIns_Inst_Sbox_9_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_9_L6), 
        .B(SubBytesIns_Inst_Sbox_9_L24), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_9_L16), 
        .B(SubBytesIns_Inst_Sbox_9_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_9_L19), 
        .B(SubBytesIns_Inst_Sbox_9_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_9_L6), 
        .B(SubBytesIns_Inst_Sbox_9_L21), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_9_L20), 
        .B(SubBytesIns_Inst_Sbox_9_L22), .Z(MixColumnsInput[11]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_9_L25), 
        .B(SubBytesIns_Inst_Sbox_9_L29), .Z(MixColumnsInput[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_9_L13), 
        .B(SubBytesIns_Inst_Sbox_9_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_9_L6), 
        .B(SubBytesIns_Inst_Sbox_9_L23), .ZN(MixColumnsInput[8]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T1_U1 ( .A(ciphertext[87]), .B(
        ciphertext[84]), .Z(SubBytesIns_Inst_Sbox_10_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T2_U1 ( .A(ciphertext[87]), .B(
        ciphertext[82]), .Z(SubBytesIns_Inst_Sbox_10_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T3_U1 ( .A(ciphertext[87]), .B(
        ciphertext[81]), .Z(SubBytesIns_Inst_Sbox_10_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T4_U1 ( .A(ciphertext[84]), .B(
        ciphertext[82]), .Z(SubBytesIns_Inst_Sbox_10_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T5_U1 ( .A(ciphertext[83]), .B(
        ciphertext[81]), .Z(SubBytesIns_Inst_Sbox_10_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_10_T1), 
        .B(SubBytesIns_Inst_Sbox_10_T5), .Z(SubBytesIns_Inst_Sbox_10_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T7_U1 ( .A(ciphertext[86]), .B(
        ciphertext[85]), .Z(SubBytesIns_Inst_Sbox_10_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T8_U1 ( .A(ciphertext[80]), .B(
        SubBytesIns_Inst_Sbox_10_T6), .Z(SubBytesIns_Inst_Sbox_10_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T9_U1 ( .A(ciphertext[80]), .B(
        SubBytesIns_Inst_Sbox_10_T7), .Z(SubBytesIns_Inst_Sbox_10_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_10_T6), .B(SubBytesIns_Inst_Sbox_10_T7), .Z(SubBytesIns_Inst_Sbox_10_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T11_U1 ( .A(ciphertext[86]), .B(
        ciphertext[82]), .Z(SubBytesIns_Inst_Sbox_10_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T12_U1 ( .A(ciphertext[85]), .B(
        ciphertext[82]), .Z(SubBytesIns_Inst_Sbox_10_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_10_T3), .B(SubBytesIns_Inst_Sbox_10_T4), .Z(SubBytesIns_Inst_Sbox_10_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_10_T6), .B(SubBytesIns_Inst_Sbox_10_T11), .Z(SubBytesIns_Inst_Sbox_10_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_10_T5), .B(SubBytesIns_Inst_Sbox_10_T11), .Z(SubBytesIns_Inst_Sbox_10_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_10_T5), .B(SubBytesIns_Inst_Sbox_10_T12), .Z(SubBytesIns_Inst_Sbox_10_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_10_T9), .B(SubBytesIns_Inst_Sbox_10_T16), .Z(SubBytesIns_Inst_Sbox_10_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T18_U1 ( .A(ciphertext[84]), .B(
        ciphertext[80]), .Z(SubBytesIns_Inst_Sbox_10_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_10_T7), .B(SubBytesIns_Inst_Sbox_10_T18), .Z(SubBytesIns_Inst_Sbox_10_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_10_T1), .B(SubBytesIns_Inst_Sbox_10_T19), .Z(SubBytesIns_Inst_Sbox_10_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T21_U1 ( .A(ciphertext[81]), .B(
        ciphertext[80]), .Z(SubBytesIns_Inst_Sbox_10_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_10_T7), .B(SubBytesIns_Inst_Sbox_10_T21), .Z(SubBytesIns_Inst_Sbox_10_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_10_T2), .B(SubBytesIns_Inst_Sbox_10_T22), .Z(SubBytesIns_Inst_Sbox_10_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_10_T2), .B(SubBytesIns_Inst_Sbox_10_T10), .Z(SubBytesIns_Inst_Sbox_10_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_T20), .B(SubBytesIns_Inst_Sbox_10_T17), .Z(
        SubBytesIns_Inst_Sbox_10_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_10_T3), .B(SubBytesIns_Inst_Sbox_10_T16), .Z(SubBytesIns_Inst_Sbox_10_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_10_T1), .B(SubBytesIns_Inst_Sbox_10_T12), .Z(SubBytesIns_Inst_Sbox_10_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T13), .A2(SubBytesIns_Inst_Sbox_10_T6), .ZN(
        SubBytesIns_Inst_Sbox_10_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T23), .A2(SubBytesIns_Inst_Sbox_10_T8), .ZN(
        SubBytesIns_Inst_Sbox_10_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_10_T14), .B(SubBytesIns_Inst_Sbox_10_M1), .Z(SubBytesIns_Inst_Sbox_10_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T19), .A2(ciphertext[80]), .ZN(
        SubBytesIns_Inst_Sbox_10_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_10_M4), 
        .B(SubBytesIns_Inst_Sbox_10_M1), .Z(SubBytesIns_Inst_Sbox_10_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_10_T3), .A2(SubBytesIns_Inst_Sbox_10_T16), .ZN(SubBytesIns_Inst_Sbox_10_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T22), .A2(SubBytesIns_Inst_Sbox_10_T9), .ZN(
        SubBytesIns_Inst_Sbox_10_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_10_T26), .B(SubBytesIns_Inst_Sbox_10_M6), .Z(SubBytesIns_Inst_Sbox_10_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T20), .A2(SubBytesIns_Inst_Sbox_10_T17), .ZN(
        SubBytesIns_Inst_Sbox_10_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_10_M9), .B(SubBytesIns_Inst_Sbox_10_M6), .Z(SubBytesIns_Inst_Sbox_10_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T1), .A2(SubBytesIns_Inst_Sbox_10_T15), .ZN(
        SubBytesIns_Inst_Sbox_10_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T4), .A2(SubBytesIns_Inst_Sbox_10_T27), .ZN(
        SubBytesIns_Inst_Sbox_10_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M12), .B(SubBytesIns_Inst_Sbox_10_M11), .Z(
        SubBytesIns_Inst_Sbox_10_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T2), .A2(SubBytesIns_Inst_Sbox_10_T10), .ZN(
        SubBytesIns_Inst_Sbox_10_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M14), .B(SubBytesIns_Inst_Sbox_10_M11), .Z(
        SubBytesIns_Inst_Sbox_10_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_10_M3), .B(SubBytesIns_Inst_Sbox_10_M2), .Z(SubBytesIns_Inst_Sbox_10_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_10_M5), .B(SubBytesIns_Inst_Sbox_10_T24), .Z(SubBytesIns_Inst_Sbox_10_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_10_M8), .B(SubBytesIns_Inst_Sbox_10_M7), .Z(SubBytesIns_Inst_Sbox_10_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M10), .B(SubBytesIns_Inst_Sbox_10_M15), .Z(
        SubBytesIns_Inst_Sbox_10_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M16), .B(SubBytesIns_Inst_Sbox_10_M13), .Z(
        SubBytesIns_Inst_Sbox_10_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M17), .B(SubBytesIns_Inst_Sbox_10_M15), .Z(
        SubBytesIns_Inst_Sbox_10_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M18), .B(SubBytesIns_Inst_Sbox_10_M13), .Z(
        SubBytesIns_Inst_Sbox_10_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M19), .B(SubBytesIns_Inst_Sbox_10_T25), .Z(
        SubBytesIns_Inst_Sbox_10_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M22), .B(SubBytesIns_Inst_Sbox_10_M23), .Z(
        SubBytesIns_Inst_Sbox_10_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M22), .A2(SubBytesIns_Inst_Sbox_10_M20), .ZN(
        SubBytesIns_Inst_Sbox_10_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M21), .B(SubBytesIns_Inst_Sbox_10_M25), .Z(
        SubBytesIns_Inst_Sbox_10_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M20), .B(SubBytesIns_Inst_Sbox_10_M21), .Z(
        SubBytesIns_Inst_Sbox_10_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M23), .B(SubBytesIns_Inst_Sbox_10_M25), .Z(
        SubBytesIns_Inst_Sbox_10_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M28), .A2(SubBytesIns_Inst_Sbox_10_M27), .ZN(
        SubBytesIns_Inst_Sbox_10_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M26), .A2(SubBytesIns_Inst_Sbox_10_M24), .ZN(
        SubBytesIns_Inst_Sbox_10_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M20), .A2(SubBytesIns_Inst_Sbox_10_M23), .ZN(
        SubBytesIns_Inst_Sbox_10_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M27), .A2(SubBytesIns_Inst_Sbox_10_M31), .ZN(
        SubBytesIns_Inst_Sbox_10_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M27), .B(SubBytesIns_Inst_Sbox_10_M25), .Z(
        SubBytesIns_Inst_Sbox_10_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M21), .A2(SubBytesIns_Inst_Sbox_10_M22), .ZN(
        SubBytesIns_Inst_Sbox_10_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M24), .A2(SubBytesIns_Inst_Sbox_10_M34), .ZN(
        SubBytesIns_Inst_Sbox_10_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M24), .B(SubBytesIns_Inst_Sbox_10_M25), .Z(
        SubBytesIns_Inst_Sbox_10_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M21), .B(SubBytesIns_Inst_Sbox_10_M29), .Z(
        SubBytesIns_Inst_Sbox_10_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M32), .B(SubBytesIns_Inst_Sbox_10_M33), .Z(
        SubBytesIns_Inst_Sbox_10_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M23), .B(SubBytesIns_Inst_Sbox_10_M30), .Z(
        SubBytesIns_Inst_Sbox_10_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M35), .B(SubBytesIns_Inst_Sbox_10_M36), .Z(
        SubBytesIns_Inst_Sbox_10_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M38), .B(SubBytesIns_Inst_Sbox_10_M40), .Z(
        SubBytesIns_Inst_Sbox_10_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M37), .B(SubBytesIns_Inst_Sbox_10_M39), .Z(
        SubBytesIns_Inst_Sbox_10_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M37), .B(SubBytesIns_Inst_Sbox_10_M38), .Z(
        SubBytesIns_Inst_Sbox_10_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M39), .B(SubBytesIns_Inst_Sbox_10_M40), .Z(
        SubBytesIns_Inst_Sbox_10_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M42), .B(SubBytesIns_Inst_Sbox_10_M41), .Z(
        SubBytesIns_Inst_Sbox_10_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M44), .A2(SubBytesIns_Inst_Sbox_10_T6), .ZN(
        SubBytesIns_Inst_Sbox_10_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M40), .A2(SubBytesIns_Inst_Sbox_10_T8), .ZN(
        SubBytesIns_Inst_Sbox_10_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M39), .A2(ciphertext[80]), .ZN(
        SubBytesIns_Inst_Sbox_10_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M43), .A2(SubBytesIns_Inst_Sbox_10_T16), .ZN(
        SubBytesIns_Inst_Sbox_10_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M38), .A2(SubBytesIns_Inst_Sbox_10_T9), .ZN(
        SubBytesIns_Inst_Sbox_10_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M37), .A2(SubBytesIns_Inst_Sbox_10_T17), .ZN(
        SubBytesIns_Inst_Sbox_10_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M42), .A2(SubBytesIns_Inst_Sbox_10_T15), .ZN(
        SubBytesIns_Inst_Sbox_10_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M45), .A2(SubBytesIns_Inst_Sbox_10_T27), .ZN(
        SubBytesIns_Inst_Sbox_10_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M41), .A2(SubBytesIns_Inst_Sbox_10_T10), .ZN(
        SubBytesIns_Inst_Sbox_10_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M44), .A2(SubBytesIns_Inst_Sbox_10_T13), .ZN(
        SubBytesIns_Inst_Sbox_10_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M40), .A2(SubBytesIns_Inst_Sbox_10_T23), .ZN(
        SubBytesIns_Inst_Sbox_10_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M39), .A2(SubBytesIns_Inst_Sbox_10_T19), .ZN(
        SubBytesIns_Inst_Sbox_10_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M43), .A2(SubBytesIns_Inst_Sbox_10_T3), .ZN(
        SubBytesIns_Inst_Sbox_10_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M38), .A2(SubBytesIns_Inst_Sbox_10_T22), .ZN(
        SubBytesIns_Inst_Sbox_10_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M37), .A2(SubBytesIns_Inst_Sbox_10_T20), .ZN(
        SubBytesIns_Inst_Sbox_10_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M42), .A2(SubBytesIns_Inst_Sbox_10_T1), .ZN(
        SubBytesIns_Inst_Sbox_10_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M45), .A2(SubBytesIns_Inst_Sbox_10_T4), .ZN(
        SubBytesIns_Inst_Sbox_10_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M41), .A2(SubBytesIns_Inst_Sbox_10_T2), .ZN(
        SubBytesIns_Inst_Sbox_10_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_10_M61), .B(SubBytesIns_Inst_Sbox_10_M62), .Z(SubBytesIns_Inst_Sbox_10_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_10_M50), .B(SubBytesIns_Inst_Sbox_10_M56), .Z(SubBytesIns_Inst_Sbox_10_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_10_M46), .B(SubBytesIns_Inst_Sbox_10_M48), .Z(SubBytesIns_Inst_Sbox_10_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_10_M47), .B(SubBytesIns_Inst_Sbox_10_M55), .Z(SubBytesIns_Inst_Sbox_10_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_10_M54), .B(SubBytesIns_Inst_Sbox_10_M58), .Z(SubBytesIns_Inst_Sbox_10_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_10_M49), .B(SubBytesIns_Inst_Sbox_10_M61), .Z(SubBytesIns_Inst_Sbox_10_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_10_M62), .B(SubBytesIns_Inst_Sbox_10_L5), .Z(SubBytesIns_Inst_Sbox_10_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_10_M46), .B(SubBytesIns_Inst_Sbox_10_L3), .Z(SubBytesIns_Inst_Sbox_10_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_10_M51), .B(SubBytesIns_Inst_Sbox_10_M59), .Z(SubBytesIns_Inst_Sbox_10_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_10_M52), .B(SubBytesIns_Inst_Sbox_10_M53), .Z(SubBytesIns_Inst_Sbox_10_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M53), .B(SubBytesIns_Inst_Sbox_10_L4), .Z(
        SubBytesIns_Inst_Sbox_10_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M60), .B(SubBytesIns_Inst_Sbox_10_L2), .Z(
        SubBytesIns_Inst_Sbox_10_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M48), .B(SubBytesIns_Inst_Sbox_10_M51), .Z(
        SubBytesIns_Inst_Sbox_10_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M50), .B(SubBytesIns_Inst_Sbox_10_L0), .Z(
        SubBytesIns_Inst_Sbox_10_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M52), .B(SubBytesIns_Inst_Sbox_10_M61), .Z(
        SubBytesIns_Inst_Sbox_10_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M55), .B(SubBytesIns_Inst_Sbox_10_L1), .Z(
        SubBytesIns_Inst_Sbox_10_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M56), .B(SubBytesIns_Inst_Sbox_10_L0), .Z(
        SubBytesIns_Inst_Sbox_10_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M57), .B(SubBytesIns_Inst_Sbox_10_L1), .Z(
        SubBytesIns_Inst_Sbox_10_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M58), .B(SubBytesIns_Inst_Sbox_10_L8), .Z(
        SubBytesIns_Inst_Sbox_10_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M63), .B(SubBytesIns_Inst_Sbox_10_L4), .Z(
        SubBytesIns_Inst_Sbox_10_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_10_L0), .B(SubBytesIns_Inst_Sbox_10_L1), .Z(SubBytesIns_Inst_Sbox_10_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_10_L1), .B(SubBytesIns_Inst_Sbox_10_L7), .Z(SubBytesIns_Inst_Sbox_10_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_10_L3), .B(SubBytesIns_Inst_Sbox_10_L12), .Z(SubBytesIns_Inst_Sbox_10_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L18), .B(SubBytesIns_Inst_Sbox_10_L2), .Z(
        SubBytesIns_Inst_Sbox_10_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L15), .B(SubBytesIns_Inst_Sbox_10_L9), .Z(
        SubBytesIns_Inst_Sbox_10_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_10_L6), .B(SubBytesIns_Inst_Sbox_10_L10), .Z(SubBytesIns_Inst_Sbox_10_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_10_L7), .B(SubBytesIns_Inst_Sbox_10_L9), .Z(SubBytesIns_Inst_Sbox_10_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_10_L8), .B(SubBytesIns_Inst_Sbox_10_L10), .Z(SubBytesIns_Inst_Sbox_10_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L11), .B(SubBytesIns_Inst_Sbox_10_L14), .Z(
        SubBytesIns_Inst_Sbox_10_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L11), .B(SubBytesIns_Inst_Sbox_10_L17), .Z(
        SubBytesIns_Inst_Sbox_10_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_10_L6), 
        .B(SubBytesIns_Inst_Sbox_10_L24), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L16), .B(SubBytesIns_Inst_Sbox_10_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L19), .B(SubBytesIns_Inst_Sbox_10_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_10_L6), 
        .B(SubBytesIns_Inst_Sbox_10_L21), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_10_L20), .B(SubBytesIns_Inst_Sbox_10_L22), .Z(MixColumnsInput[115]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_10_L25), .B(SubBytesIns_Inst_Sbox_10_L29), .Z(MixColumnsInput[114]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L13), .B(SubBytesIns_Inst_Sbox_10_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_10_L6), .B(SubBytesIns_Inst_Sbox_10_L23), .ZN(MixColumnsInput[112]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T1_U1 ( .A(ciphertext[95]), .B(
        ciphertext[92]), .Z(SubBytesIns_Inst_Sbox_11_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T2_U1 ( .A(ciphertext[95]), .B(
        ciphertext[90]), .Z(SubBytesIns_Inst_Sbox_11_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T3_U1 ( .A(ciphertext[95]), .B(
        ciphertext[89]), .Z(SubBytesIns_Inst_Sbox_11_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T4_U1 ( .A(ciphertext[92]), .B(
        ciphertext[90]), .Z(SubBytesIns_Inst_Sbox_11_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T5_U1 ( .A(ciphertext[91]), .B(
        ciphertext[89]), .Z(SubBytesIns_Inst_Sbox_11_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_11_T1), 
        .B(SubBytesIns_Inst_Sbox_11_T5), .Z(SubBytesIns_Inst_Sbox_11_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T7_U1 ( .A(ciphertext[94]), .B(
        ciphertext[93]), .Z(SubBytesIns_Inst_Sbox_11_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T8_U1 ( .A(ciphertext[88]), .B(
        SubBytesIns_Inst_Sbox_11_T6), .Z(SubBytesIns_Inst_Sbox_11_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T9_U1 ( .A(ciphertext[88]), .B(
        SubBytesIns_Inst_Sbox_11_T7), .Z(SubBytesIns_Inst_Sbox_11_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_11_T6), .B(SubBytesIns_Inst_Sbox_11_T7), .Z(SubBytesIns_Inst_Sbox_11_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T11_U1 ( .A(ciphertext[94]), .B(
        ciphertext[90]), .Z(SubBytesIns_Inst_Sbox_11_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T12_U1 ( .A(ciphertext[93]), .B(
        ciphertext[90]), .Z(SubBytesIns_Inst_Sbox_11_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_11_T3), .B(SubBytesIns_Inst_Sbox_11_T4), .Z(SubBytesIns_Inst_Sbox_11_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_11_T6), .B(SubBytesIns_Inst_Sbox_11_T11), .Z(SubBytesIns_Inst_Sbox_11_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_11_T5), .B(SubBytesIns_Inst_Sbox_11_T11), .Z(SubBytesIns_Inst_Sbox_11_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_11_T5), .B(SubBytesIns_Inst_Sbox_11_T12), .Z(SubBytesIns_Inst_Sbox_11_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_11_T9), .B(SubBytesIns_Inst_Sbox_11_T16), .Z(SubBytesIns_Inst_Sbox_11_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T18_U1 ( .A(ciphertext[92]), .B(
        ciphertext[88]), .Z(SubBytesIns_Inst_Sbox_11_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_11_T7), .B(SubBytesIns_Inst_Sbox_11_T18), .Z(SubBytesIns_Inst_Sbox_11_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_11_T1), .B(SubBytesIns_Inst_Sbox_11_T19), .Z(SubBytesIns_Inst_Sbox_11_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T21_U1 ( .A(ciphertext[89]), .B(
        ciphertext[88]), .Z(SubBytesIns_Inst_Sbox_11_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_11_T7), .B(SubBytesIns_Inst_Sbox_11_T21), .Z(SubBytesIns_Inst_Sbox_11_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_11_T2), .B(SubBytesIns_Inst_Sbox_11_T22), .Z(SubBytesIns_Inst_Sbox_11_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_11_T2), .B(SubBytesIns_Inst_Sbox_11_T10), .Z(SubBytesIns_Inst_Sbox_11_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_T20), .B(SubBytesIns_Inst_Sbox_11_T17), .Z(
        SubBytesIns_Inst_Sbox_11_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_11_T3), .B(SubBytesIns_Inst_Sbox_11_T16), .Z(SubBytesIns_Inst_Sbox_11_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_11_T1), .B(SubBytesIns_Inst_Sbox_11_T12), .Z(SubBytesIns_Inst_Sbox_11_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T13), .A2(SubBytesIns_Inst_Sbox_11_T6), .ZN(
        SubBytesIns_Inst_Sbox_11_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T23), .A2(SubBytesIns_Inst_Sbox_11_T8), .ZN(
        SubBytesIns_Inst_Sbox_11_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_11_T14), .B(SubBytesIns_Inst_Sbox_11_M1), .Z(SubBytesIns_Inst_Sbox_11_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T19), .A2(ciphertext[88]), .ZN(
        SubBytesIns_Inst_Sbox_11_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_11_M4), 
        .B(SubBytesIns_Inst_Sbox_11_M1), .Z(SubBytesIns_Inst_Sbox_11_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_11_T3), .A2(SubBytesIns_Inst_Sbox_11_T16), .ZN(SubBytesIns_Inst_Sbox_11_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T22), .A2(SubBytesIns_Inst_Sbox_11_T9), .ZN(
        SubBytesIns_Inst_Sbox_11_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_11_T26), .B(SubBytesIns_Inst_Sbox_11_M6), .Z(SubBytesIns_Inst_Sbox_11_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T20), .A2(SubBytesIns_Inst_Sbox_11_T17), .ZN(
        SubBytesIns_Inst_Sbox_11_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_11_M9), .B(SubBytesIns_Inst_Sbox_11_M6), .Z(SubBytesIns_Inst_Sbox_11_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T1), .A2(SubBytesIns_Inst_Sbox_11_T15), .ZN(
        SubBytesIns_Inst_Sbox_11_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T4), .A2(SubBytesIns_Inst_Sbox_11_T27), .ZN(
        SubBytesIns_Inst_Sbox_11_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M12), .B(SubBytesIns_Inst_Sbox_11_M11), .Z(
        SubBytesIns_Inst_Sbox_11_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T2), .A2(SubBytesIns_Inst_Sbox_11_T10), .ZN(
        SubBytesIns_Inst_Sbox_11_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M14), .B(SubBytesIns_Inst_Sbox_11_M11), .Z(
        SubBytesIns_Inst_Sbox_11_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_11_M3), .B(SubBytesIns_Inst_Sbox_11_M2), .Z(SubBytesIns_Inst_Sbox_11_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_11_M5), .B(SubBytesIns_Inst_Sbox_11_T24), .Z(SubBytesIns_Inst_Sbox_11_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_11_M8), .B(SubBytesIns_Inst_Sbox_11_M7), .Z(SubBytesIns_Inst_Sbox_11_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M10), .B(SubBytesIns_Inst_Sbox_11_M15), .Z(
        SubBytesIns_Inst_Sbox_11_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M16), .B(SubBytesIns_Inst_Sbox_11_M13), .Z(
        SubBytesIns_Inst_Sbox_11_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M17), .B(SubBytesIns_Inst_Sbox_11_M15), .Z(
        SubBytesIns_Inst_Sbox_11_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M18), .B(SubBytesIns_Inst_Sbox_11_M13), .Z(
        SubBytesIns_Inst_Sbox_11_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M19), .B(SubBytesIns_Inst_Sbox_11_T25), .Z(
        SubBytesIns_Inst_Sbox_11_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M22), .B(SubBytesIns_Inst_Sbox_11_M23), .Z(
        SubBytesIns_Inst_Sbox_11_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M22), .A2(SubBytesIns_Inst_Sbox_11_M20), .ZN(
        SubBytesIns_Inst_Sbox_11_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M21), .B(SubBytesIns_Inst_Sbox_11_M25), .Z(
        SubBytesIns_Inst_Sbox_11_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M20), .B(SubBytesIns_Inst_Sbox_11_M21), .Z(
        SubBytesIns_Inst_Sbox_11_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M23), .B(SubBytesIns_Inst_Sbox_11_M25), .Z(
        SubBytesIns_Inst_Sbox_11_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M28), .A2(SubBytesIns_Inst_Sbox_11_M27), .ZN(
        SubBytesIns_Inst_Sbox_11_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M26), .A2(SubBytesIns_Inst_Sbox_11_M24), .ZN(
        SubBytesIns_Inst_Sbox_11_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M20), .A2(SubBytesIns_Inst_Sbox_11_M23), .ZN(
        SubBytesIns_Inst_Sbox_11_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M27), .A2(SubBytesIns_Inst_Sbox_11_M31), .ZN(
        SubBytesIns_Inst_Sbox_11_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M27), .B(SubBytesIns_Inst_Sbox_11_M25), .Z(
        SubBytesIns_Inst_Sbox_11_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M21), .A2(SubBytesIns_Inst_Sbox_11_M22), .ZN(
        SubBytesIns_Inst_Sbox_11_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M24), .A2(SubBytesIns_Inst_Sbox_11_M34), .ZN(
        SubBytesIns_Inst_Sbox_11_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M24), .B(SubBytesIns_Inst_Sbox_11_M25), .Z(
        SubBytesIns_Inst_Sbox_11_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M21), .B(SubBytesIns_Inst_Sbox_11_M29), .Z(
        SubBytesIns_Inst_Sbox_11_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M32), .B(SubBytesIns_Inst_Sbox_11_M33), .Z(
        SubBytesIns_Inst_Sbox_11_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M23), .B(SubBytesIns_Inst_Sbox_11_M30), .Z(
        SubBytesIns_Inst_Sbox_11_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M35), .B(SubBytesIns_Inst_Sbox_11_M36), .Z(
        SubBytesIns_Inst_Sbox_11_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M38), .B(SubBytesIns_Inst_Sbox_11_M40), .Z(
        SubBytesIns_Inst_Sbox_11_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M37), .B(SubBytesIns_Inst_Sbox_11_M39), .Z(
        SubBytesIns_Inst_Sbox_11_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M37), .B(SubBytesIns_Inst_Sbox_11_M38), .Z(
        SubBytesIns_Inst_Sbox_11_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M39), .B(SubBytesIns_Inst_Sbox_11_M40), .Z(
        SubBytesIns_Inst_Sbox_11_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M42), .B(SubBytesIns_Inst_Sbox_11_M41), .Z(
        SubBytesIns_Inst_Sbox_11_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M44), .A2(SubBytesIns_Inst_Sbox_11_T6), .ZN(
        SubBytesIns_Inst_Sbox_11_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M40), .A2(SubBytesIns_Inst_Sbox_11_T8), .ZN(
        SubBytesIns_Inst_Sbox_11_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M39), .A2(ciphertext[88]), .ZN(
        SubBytesIns_Inst_Sbox_11_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M43), .A2(SubBytesIns_Inst_Sbox_11_T16), .ZN(
        SubBytesIns_Inst_Sbox_11_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M38), .A2(SubBytesIns_Inst_Sbox_11_T9), .ZN(
        SubBytesIns_Inst_Sbox_11_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M37), .A2(SubBytesIns_Inst_Sbox_11_T17), .ZN(
        SubBytesIns_Inst_Sbox_11_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M42), .A2(SubBytesIns_Inst_Sbox_11_T15), .ZN(
        SubBytesIns_Inst_Sbox_11_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M45), .A2(SubBytesIns_Inst_Sbox_11_T27), .ZN(
        SubBytesIns_Inst_Sbox_11_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M41), .A2(SubBytesIns_Inst_Sbox_11_T10), .ZN(
        SubBytesIns_Inst_Sbox_11_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M44), .A2(SubBytesIns_Inst_Sbox_11_T13), .ZN(
        SubBytesIns_Inst_Sbox_11_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M40), .A2(SubBytesIns_Inst_Sbox_11_T23), .ZN(
        SubBytesIns_Inst_Sbox_11_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M39), .A2(SubBytesIns_Inst_Sbox_11_T19), .ZN(
        SubBytesIns_Inst_Sbox_11_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M43), .A2(SubBytesIns_Inst_Sbox_11_T3), .ZN(
        SubBytesIns_Inst_Sbox_11_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M38), .A2(SubBytesIns_Inst_Sbox_11_T22), .ZN(
        SubBytesIns_Inst_Sbox_11_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M37), .A2(SubBytesIns_Inst_Sbox_11_T20), .ZN(
        SubBytesIns_Inst_Sbox_11_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M42), .A2(SubBytesIns_Inst_Sbox_11_T1), .ZN(
        SubBytesIns_Inst_Sbox_11_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M45), .A2(SubBytesIns_Inst_Sbox_11_T4), .ZN(
        SubBytesIns_Inst_Sbox_11_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M41), .A2(SubBytesIns_Inst_Sbox_11_T2), .ZN(
        SubBytesIns_Inst_Sbox_11_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_11_M61), .B(SubBytesIns_Inst_Sbox_11_M62), .Z(SubBytesIns_Inst_Sbox_11_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_11_M50), .B(SubBytesIns_Inst_Sbox_11_M56), .Z(SubBytesIns_Inst_Sbox_11_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_11_M46), .B(SubBytesIns_Inst_Sbox_11_M48), .Z(SubBytesIns_Inst_Sbox_11_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_11_M47), .B(SubBytesIns_Inst_Sbox_11_M55), .Z(SubBytesIns_Inst_Sbox_11_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_11_M54), .B(SubBytesIns_Inst_Sbox_11_M58), .Z(SubBytesIns_Inst_Sbox_11_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_11_M49), .B(SubBytesIns_Inst_Sbox_11_M61), .Z(SubBytesIns_Inst_Sbox_11_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_11_M62), .B(SubBytesIns_Inst_Sbox_11_L5), .Z(SubBytesIns_Inst_Sbox_11_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_11_M46), .B(SubBytesIns_Inst_Sbox_11_L3), .Z(SubBytesIns_Inst_Sbox_11_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_11_M51), .B(SubBytesIns_Inst_Sbox_11_M59), .Z(SubBytesIns_Inst_Sbox_11_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_11_M52), .B(SubBytesIns_Inst_Sbox_11_M53), .Z(SubBytesIns_Inst_Sbox_11_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M53), .B(SubBytesIns_Inst_Sbox_11_L4), .Z(
        SubBytesIns_Inst_Sbox_11_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M60), .B(SubBytesIns_Inst_Sbox_11_L2), .Z(
        SubBytesIns_Inst_Sbox_11_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M48), .B(SubBytesIns_Inst_Sbox_11_M51), .Z(
        SubBytesIns_Inst_Sbox_11_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M50), .B(SubBytesIns_Inst_Sbox_11_L0), .Z(
        SubBytesIns_Inst_Sbox_11_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M52), .B(SubBytesIns_Inst_Sbox_11_M61), .Z(
        SubBytesIns_Inst_Sbox_11_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M55), .B(SubBytesIns_Inst_Sbox_11_L1), .Z(
        SubBytesIns_Inst_Sbox_11_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M56), .B(SubBytesIns_Inst_Sbox_11_L0), .Z(
        SubBytesIns_Inst_Sbox_11_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M57), .B(SubBytesIns_Inst_Sbox_11_L1), .Z(
        SubBytesIns_Inst_Sbox_11_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M58), .B(SubBytesIns_Inst_Sbox_11_L8), .Z(
        SubBytesIns_Inst_Sbox_11_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M63), .B(SubBytesIns_Inst_Sbox_11_L4), .Z(
        SubBytesIns_Inst_Sbox_11_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_11_L0), .B(SubBytesIns_Inst_Sbox_11_L1), .Z(SubBytesIns_Inst_Sbox_11_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_11_L1), .B(SubBytesIns_Inst_Sbox_11_L7), .Z(SubBytesIns_Inst_Sbox_11_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_11_L3), .B(SubBytesIns_Inst_Sbox_11_L12), .Z(SubBytesIns_Inst_Sbox_11_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L18), .B(SubBytesIns_Inst_Sbox_11_L2), .Z(
        SubBytesIns_Inst_Sbox_11_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L15), .B(SubBytesIns_Inst_Sbox_11_L9), .Z(
        SubBytesIns_Inst_Sbox_11_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_11_L6), .B(SubBytesIns_Inst_Sbox_11_L10), .Z(SubBytesIns_Inst_Sbox_11_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_11_L7), .B(SubBytesIns_Inst_Sbox_11_L9), .Z(SubBytesIns_Inst_Sbox_11_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_11_L8), .B(SubBytesIns_Inst_Sbox_11_L10), .Z(SubBytesIns_Inst_Sbox_11_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L11), .B(SubBytesIns_Inst_Sbox_11_L14), .Z(
        SubBytesIns_Inst_Sbox_11_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L11), .B(SubBytesIns_Inst_Sbox_11_L17), .Z(
        SubBytesIns_Inst_Sbox_11_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_11_L6), 
        .B(SubBytesIns_Inst_Sbox_11_L24), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L16), .B(SubBytesIns_Inst_Sbox_11_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L19), .B(SubBytesIns_Inst_Sbox_11_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_11_L6), 
        .B(SubBytesIns_Inst_Sbox_11_L21), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_11_L20), .B(SubBytesIns_Inst_Sbox_11_L22), .Z(MixColumnsInput[91]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_11_L25), .B(SubBytesIns_Inst_Sbox_11_L29), .Z(MixColumnsInput[90]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L13), .B(SubBytesIns_Inst_Sbox_11_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_11_L6), .B(SubBytesIns_Inst_Sbox_11_L23), .ZN(MixColumnsInput[88]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T1_U1 ( .A(ciphertext[103]), .B(
        ciphertext[100]), .Z(SubBytesIns_Inst_Sbox_12_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T2_U1 ( .A(ciphertext[103]), .B(
        ciphertext[98]), .Z(SubBytesIns_Inst_Sbox_12_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T3_U1 ( .A(ciphertext[103]), .B(
        ciphertext[97]), .Z(SubBytesIns_Inst_Sbox_12_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T4_U1 ( .A(ciphertext[100]), .B(
        ciphertext[98]), .Z(SubBytesIns_Inst_Sbox_12_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T5_U1 ( .A(ciphertext[99]), .B(
        ciphertext[97]), .Z(SubBytesIns_Inst_Sbox_12_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_12_T1), 
        .B(SubBytesIns_Inst_Sbox_12_T5), .Z(SubBytesIns_Inst_Sbox_12_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T7_U1 ( .A(ciphertext[102]), .B(
        ciphertext[101]), .Z(SubBytesIns_Inst_Sbox_12_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T8_U1 ( .A(ciphertext[96]), .B(
        SubBytesIns_Inst_Sbox_12_T6), .Z(SubBytesIns_Inst_Sbox_12_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T9_U1 ( .A(ciphertext[96]), .B(
        SubBytesIns_Inst_Sbox_12_T7), .Z(SubBytesIns_Inst_Sbox_12_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_12_T6), .B(SubBytesIns_Inst_Sbox_12_T7), .Z(SubBytesIns_Inst_Sbox_12_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T11_U1 ( .A(ciphertext[102]), .B(
        ciphertext[98]), .Z(SubBytesIns_Inst_Sbox_12_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T12_U1 ( .A(ciphertext[101]), .B(
        ciphertext[98]), .Z(SubBytesIns_Inst_Sbox_12_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_12_T3), .B(SubBytesIns_Inst_Sbox_12_T4), .Z(SubBytesIns_Inst_Sbox_12_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_12_T6), .B(SubBytesIns_Inst_Sbox_12_T11), .Z(SubBytesIns_Inst_Sbox_12_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_12_T5), .B(SubBytesIns_Inst_Sbox_12_T11), .Z(SubBytesIns_Inst_Sbox_12_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_12_T5), .B(SubBytesIns_Inst_Sbox_12_T12), .Z(SubBytesIns_Inst_Sbox_12_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_12_T9), .B(SubBytesIns_Inst_Sbox_12_T16), .Z(SubBytesIns_Inst_Sbox_12_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T18_U1 ( .A(ciphertext[100]), .B(
        ciphertext[96]), .Z(SubBytesIns_Inst_Sbox_12_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_12_T7), .B(SubBytesIns_Inst_Sbox_12_T18), .Z(SubBytesIns_Inst_Sbox_12_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_12_T1), .B(SubBytesIns_Inst_Sbox_12_T19), .Z(SubBytesIns_Inst_Sbox_12_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T21_U1 ( .A(ciphertext[97]), .B(
        ciphertext[96]), .Z(SubBytesIns_Inst_Sbox_12_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_12_T7), .B(SubBytesIns_Inst_Sbox_12_T21), .Z(SubBytesIns_Inst_Sbox_12_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_12_T2), .B(SubBytesIns_Inst_Sbox_12_T22), .Z(SubBytesIns_Inst_Sbox_12_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_12_T2), .B(SubBytesIns_Inst_Sbox_12_T10), .Z(SubBytesIns_Inst_Sbox_12_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_T20), .B(SubBytesIns_Inst_Sbox_12_T17), .Z(
        SubBytesIns_Inst_Sbox_12_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_12_T3), .B(SubBytesIns_Inst_Sbox_12_T16), .Z(SubBytesIns_Inst_Sbox_12_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_12_T1), .B(SubBytesIns_Inst_Sbox_12_T12), .Z(SubBytesIns_Inst_Sbox_12_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T13), .A2(SubBytesIns_Inst_Sbox_12_T6), .ZN(
        SubBytesIns_Inst_Sbox_12_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T23), .A2(SubBytesIns_Inst_Sbox_12_T8), .ZN(
        SubBytesIns_Inst_Sbox_12_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_12_T14), .B(SubBytesIns_Inst_Sbox_12_M1), .Z(SubBytesIns_Inst_Sbox_12_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T19), .A2(ciphertext[96]), .ZN(
        SubBytesIns_Inst_Sbox_12_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_12_M4), 
        .B(SubBytesIns_Inst_Sbox_12_M1), .Z(SubBytesIns_Inst_Sbox_12_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_12_T3), .A2(SubBytesIns_Inst_Sbox_12_T16), .ZN(SubBytesIns_Inst_Sbox_12_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T22), .A2(SubBytesIns_Inst_Sbox_12_T9), .ZN(
        SubBytesIns_Inst_Sbox_12_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_12_T26), .B(SubBytesIns_Inst_Sbox_12_M6), .Z(SubBytesIns_Inst_Sbox_12_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T20), .A2(SubBytesIns_Inst_Sbox_12_T17), .ZN(
        SubBytesIns_Inst_Sbox_12_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_12_M9), .B(SubBytesIns_Inst_Sbox_12_M6), .Z(SubBytesIns_Inst_Sbox_12_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T1), .A2(SubBytesIns_Inst_Sbox_12_T15), .ZN(
        SubBytesIns_Inst_Sbox_12_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T4), .A2(SubBytesIns_Inst_Sbox_12_T27), .ZN(
        SubBytesIns_Inst_Sbox_12_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M12), .B(SubBytesIns_Inst_Sbox_12_M11), .Z(
        SubBytesIns_Inst_Sbox_12_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T2), .A2(SubBytesIns_Inst_Sbox_12_T10), .ZN(
        SubBytesIns_Inst_Sbox_12_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M14), .B(SubBytesIns_Inst_Sbox_12_M11), .Z(
        SubBytesIns_Inst_Sbox_12_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_12_M3), .B(SubBytesIns_Inst_Sbox_12_M2), .Z(SubBytesIns_Inst_Sbox_12_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_12_M5), .B(SubBytesIns_Inst_Sbox_12_T24), .Z(SubBytesIns_Inst_Sbox_12_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_12_M8), .B(SubBytesIns_Inst_Sbox_12_M7), .Z(SubBytesIns_Inst_Sbox_12_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M10), .B(SubBytesIns_Inst_Sbox_12_M15), .Z(
        SubBytesIns_Inst_Sbox_12_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M16), .B(SubBytesIns_Inst_Sbox_12_M13), .Z(
        SubBytesIns_Inst_Sbox_12_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M17), .B(SubBytesIns_Inst_Sbox_12_M15), .Z(
        SubBytesIns_Inst_Sbox_12_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M18), .B(SubBytesIns_Inst_Sbox_12_M13), .Z(
        SubBytesIns_Inst_Sbox_12_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M19), .B(SubBytesIns_Inst_Sbox_12_T25), .Z(
        SubBytesIns_Inst_Sbox_12_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M22), .B(SubBytesIns_Inst_Sbox_12_M23), .Z(
        SubBytesIns_Inst_Sbox_12_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M22), .A2(SubBytesIns_Inst_Sbox_12_M20), .ZN(
        SubBytesIns_Inst_Sbox_12_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M21), .B(SubBytesIns_Inst_Sbox_12_M25), .Z(
        SubBytesIns_Inst_Sbox_12_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M20), .B(SubBytesIns_Inst_Sbox_12_M21), .Z(
        SubBytesIns_Inst_Sbox_12_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M23), .B(SubBytesIns_Inst_Sbox_12_M25), .Z(
        SubBytesIns_Inst_Sbox_12_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M28), .A2(SubBytesIns_Inst_Sbox_12_M27), .ZN(
        SubBytesIns_Inst_Sbox_12_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M26), .A2(SubBytesIns_Inst_Sbox_12_M24), .ZN(
        SubBytesIns_Inst_Sbox_12_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M20), .A2(SubBytesIns_Inst_Sbox_12_M23), .ZN(
        SubBytesIns_Inst_Sbox_12_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M27), .A2(SubBytesIns_Inst_Sbox_12_M31), .ZN(
        SubBytesIns_Inst_Sbox_12_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M27), .B(SubBytesIns_Inst_Sbox_12_M25), .Z(
        SubBytesIns_Inst_Sbox_12_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M21), .A2(SubBytesIns_Inst_Sbox_12_M22), .ZN(
        SubBytesIns_Inst_Sbox_12_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M24), .A2(SubBytesIns_Inst_Sbox_12_M34), .ZN(
        SubBytesIns_Inst_Sbox_12_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M24), .B(SubBytesIns_Inst_Sbox_12_M25), .Z(
        SubBytesIns_Inst_Sbox_12_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M21), .B(SubBytesIns_Inst_Sbox_12_M29), .Z(
        SubBytesIns_Inst_Sbox_12_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M32), .B(SubBytesIns_Inst_Sbox_12_M33), .Z(
        SubBytesIns_Inst_Sbox_12_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M23), .B(SubBytesIns_Inst_Sbox_12_M30), .Z(
        SubBytesIns_Inst_Sbox_12_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M35), .B(SubBytesIns_Inst_Sbox_12_M36), .Z(
        SubBytesIns_Inst_Sbox_12_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M38), .B(SubBytesIns_Inst_Sbox_12_M40), .Z(
        SubBytesIns_Inst_Sbox_12_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M37), .B(SubBytesIns_Inst_Sbox_12_M39), .Z(
        SubBytesIns_Inst_Sbox_12_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M37), .B(SubBytesIns_Inst_Sbox_12_M38), .Z(
        SubBytesIns_Inst_Sbox_12_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M39), .B(SubBytesIns_Inst_Sbox_12_M40), .Z(
        SubBytesIns_Inst_Sbox_12_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M42), .B(SubBytesIns_Inst_Sbox_12_M41), .Z(
        SubBytesIns_Inst_Sbox_12_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M44), .A2(SubBytesIns_Inst_Sbox_12_T6), .ZN(
        SubBytesIns_Inst_Sbox_12_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M40), .A2(SubBytesIns_Inst_Sbox_12_T8), .ZN(
        SubBytesIns_Inst_Sbox_12_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M39), .A2(ciphertext[96]), .ZN(
        SubBytesIns_Inst_Sbox_12_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M43), .A2(SubBytesIns_Inst_Sbox_12_T16), .ZN(
        SubBytesIns_Inst_Sbox_12_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M38), .A2(SubBytesIns_Inst_Sbox_12_T9), .ZN(
        SubBytesIns_Inst_Sbox_12_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M37), .A2(SubBytesIns_Inst_Sbox_12_T17), .ZN(
        SubBytesIns_Inst_Sbox_12_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M42), .A2(SubBytesIns_Inst_Sbox_12_T15), .ZN(
        SubBytesIns_Inst_Sbox_12_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M45), .A2(SubBytesIns_Inst_Sbox_12_T27), .ZN(
        SubBytesIns_Inst_Sbox_12_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M41), .A2(SubBytesIns_Inst_Sbox_12_T10), .ZN(
        SubBytesIns_Inst_Sbox_12_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M44), .A2(SubBytesIns_Inst_Sbox_12_T13), .ZN(
        SubBytesIns_Inst_Sbox_12_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M40), .A2(SubBytesIns_Inst_Sbox_12_T23), .ZN(
        SubBytesIns_Inst_Sbox_12_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M39), .A2(SubBytesIns_Inst_Sbox_12_T19), .ZN(
        SubBytesIns_Inst_Sbox_12_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M43), .A2(SubBytesIns_Inst_Sbox_12_T3), .ZN(
        SubBytesIns_Inst_Sbox_12_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M38), .A2(SubBytesIns_Inst_Sbox_12_T22), .ZN(
        SubBytesIns_Inst_Sbox_12_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M37), .A2(SubBytesIns_Inst_Sbox_12_T20), .ZN(
        SubBytesIns_Inst_Sbox_12_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M42), .A2(SubBytesIns_Inst_Sbox_12_T1), .ZN(
        SubBytesIns_Inst_Sbox_12_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M45), .A2(SubBytesIns_Inst_Sbox_12_T4), .ZN(
        SubBytesIns_Inst_Sbox_12_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M41), .A2(SubBytesIns_Inst_Sbox_12_T2), .ZN(
        SubBytesIns_Inst_Sbox_12_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_12_M61), .B(SubBytesIns_Inst_Sbox_12_M62), .Z(SubBytesIns_Inst_Sbox_12_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_12_M50), .B(SubBytesIns_Inst_Sbox_12_M56), .Z(SubBytesIns_Inst_Sbox_12_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_12_M46), .B(SubBytesIns_Inst_Sbox_12_M48), .Z(SubBytesIns_Inst_Sbox_12_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_12_M47), .B(SubBytesIns_Inst_Sbox_12_M55), .Z(SubBytesIns_Inst_Sbox_12_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_12_M54), .B(SubBytesIns_Inst_Sbox_12_M58), .Z(SubBytesIns_Inst_Sbox_12_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_12_M49), .B(SubBytesIns_Inst_Sbox_12_M61), .Z(SubBytesIns_Inst_Sbox_12_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_12_M62), .B(SubBytesIns_Inst_Sbox_12_L5), .Z(SubBytesIns_Inst_Sbox_12_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_12_M46), .B(SubBytesIns_Inst_Sbox_12_L3), .Z(SubBytesIns_Inst_Sbox_12_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_12_M51), .B(SubBytesIns_Inst_Sbox_12_M59), .Z(SubBytesIns_Inst_Sbox_12_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_12_M52), .B(SubBytesIns_Inst_Sbox_12_M53), .Z(SubBytesIns_Inst_Sbox_12_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M53), .B(SubBytesIns_Inst_Sbox_12_L4), .Z(
        SubBytesIns_Inst_Sbox_12_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M60), .B(SubBytesIns_Inst_Sbox_12_L2), .Z(
        SubBytesIns_Inst_Sbox_12_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M48), .B(SubBytesIns_Inst_Sbox_12_M51), .Z(
        SubBytesIns_Inst_Sbox_12_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M50), .B(SubBytesIns_Inst_Sbox_12_L0), .Z(
        SubBytesIns_Inst_Sbox_12_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M52), .B(SubBytesIns_Inst_Sbox_12_M61), .Z(
        SubBytesIns_Inst_Sbox_12_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M55), .B(SubBytesIns_Inst_Sbox_12_L1), .Z(
        SubBytesIns_Inst_Sbox_12_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M56), .B(SubBytesIns_Inst_Sbox_12_L0), .Z(
        SubBytesIns_Inst_Sbox_12_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M57), .B(SubBytesIns_Inst_Sbox_12_L1), .Z(
        SubBytesIns_Inst_Sbox_12_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M58), .B(SubBytesIns_Inst_Sbox_12_L8), .Z(
        SubBytesIns_Inst_Sbox_12_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M63), .B(SubBytesIns_Inst_Sbox_12_L4), .Z(
        SubBytesIns_Inst_Sbox_12_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_12_L0), .B(SubBytesIns_Inst_Sbox_12_L1), .Z(SubBytesIns_Inst_Sbox_12_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_12_L1), .B(SubBytesIns_Inst_Sbox_12_L7), .Z(SubBytesIns_Inst_Sbox_12_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_12_L3), .B(SubBytesIns_Inst_Sbox_12_L12), .Z(SubBytesIns_Inst_Sbox_12_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L18), .B(SubBytesIns_Inst_Sbox_12_L2), .Z(
        SubBytesIns_Inst_Sbox_12_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L15), .B(SubBytesIns_Inst_Sbox_12_L9), .Z(
        SubBytesIns_Inst_Sbox_12_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_12_L6), .B(SubBytesIns_Inst_Sbox_12_L10), .Z(SubBytesIns_Inst_Sbox_12_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_12_L7), .B(SubBytesIns_Inst_Sbox_12_L9), .Z(SubBytesIns_Inst_Sbox_12_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_12_L8), .B(SubBytesIns_Inst_Sbox_12_L10), .Z(SubBytesIns_Inst_Sbox_12_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L11), .B(SubBytesIns_Inst_Sbox_12_L14), .Z(
        SubBytesIns_Inst_Sbox_12_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L11), .B(SubBytesIns_Inst_Sbox_12_L17), .Z(
        SubBytesIns_Inst_Sbox_12_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_12_L6), 
        .B(SubBytesIns_Inst_Sbox_12_L24), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L16), .B(SubBytesIns_Inst_Sbox_12_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L19), .B(SubBytesIns_Inst_Sbox_12_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_12_L6), 
        .B(SubBytesIns_Inst_Sbox_12_L21), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_12_L20), .B(SubBytesIns_Inst_Sbox_12_L22), .Z(MixColumnsInput[67]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_12_L25), .B(SubBytesIns_Inst_Sbox_12_L29), .Z(MixColumnsInput[66]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L13), .B(SubBytesIns_Inst_Sbox_12_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_12_L6), .B(SubBytesIns_Inst_Sbox_12_L23), .ZN(MixColumnsInput[64]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T1_U1 ( .A(ciphertext[111]), .B(
        ciphertext[108]), .Z(SubBytesIns_Inst_Sbox_13_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T2_U1 ( .A(ciphertext[111]), .B(
        ciphertext[106]), .Z(SubBytesIns_Inst_Sbox_13_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T3_U1 ( .A(ciphertext[111]), .B(
        ciphertext[105]), .Z(SubBytesIns_Inst_Sbox_13_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T4_U1 ( .A(ciphertext[108]), .B(
        ciphertext[106]), .Z(SubBytesIns_Inst_Sbox_13_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T5_U1 ( .A(ciphertext[107]), .B(
        ciphertext[105]), .Z(SubBytesIns_Inst_Sbox_13_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_13_T1), 
        .B(SubBytesIns_Inst_Sbox_13_T5), .Z(SubBytesIns_Inst_Sbox_13_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T7_U1 ( .A(ciphertext[110]), .B(
        ciphertext[109]), .Z(SubBytesIns_Inst_Sbox_13_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T8_U1 ( .A(ciphertext[104]), .B(
        SubBytesIns_Inst_Sbox_13_T6), .Z(SubBytesIns_Inst_Sbox_13_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T9_U1 ( .A(ciphertext[104]), .B(
        SubBytesIns_Inst_Sbox_13_T7), .Z(SubBytesIns_Inst_Sbox_13_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_13_T6), .B(SubBytesIns_Inst_Sbox_13_T7), .Z(SubBytesIns_Inst_Sbox_13_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T11_U1 ( .A(ciphertext[110]), .B(
        ciphertext[106]), .Z(SubBytesIns_Inst_Sbox_13_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T12_U1 ( .A(ciphertext[109]), .B(
        ciphertext[106]), .Z(SubBytesIns_Inst_Sbox_13_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_13_T3), .B(SubBytesIns_Inst_Sbox_13_T4), .Z(SubBytesIns_Inst_Sbox_13_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_13_T6), .B(SubBytesIns_Inst_Sbox_13_T11), .Z(SubBytesIns_Inst_Sbox_13_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_13_T5), .B(SubBytesIns_Inst_Sbox_13_T11), .Z(SubBytesIns_Inst_Sbox_13_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_13_T5), .B(SubBytesIns_Inst_Sbox_13_T12), .Z(SubBytesIns_Inst_Sbox_13_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_13_T9), .B(SubBytesIns_Inst_Sbox_13_T16), .Z(SubBytesIns_Inst_Sbox_13_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T18_U1 ( .A(ciphertext[108]), .B(
        ciphertext[104]), .Z(SubBytesIns_Inst_Sbox_13_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_13_T7), .B(SubBytesIns_Inst_Sbox_13_T18), .Z(SubBytesIns_Inst_Sbox_13_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_13_T1), .B(SubBytesIns_Inst_Sbox_13_T19), .Z(SubBytesIns_Inst_Sbox_13_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T21_U1 ( .A(ciphertext[105]), .B(
        ciphertext[104]), .Z(SubBytesIns_Inst_Sbox_13_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_13_T7), .B(SubBytesIns_Inst_Sbox_13_T21), .Z(SubBytesIns_Inst_Sbox_13_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_13_T2), .B(SubBytesIns_Inst_Sbox_13_T22), .Z(SubBytesIns_Inst_Sbox_13_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_13_T2), .B(SubBytesIns_Inst_Sbox_13_T10), .Z(SubBytesIns_Inst_Sbox_13_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_T20), .B(SubBytesIns_Inst_Sbox_13_T17), .Z(
        SubBytesIns_Inst_Sbox_13_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_13_T3), .B(SubBytesIns_Inst_Sbox_13_T16), .Z(SubBytesIns_Inst_Sbox_13_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_13_T1), .B(SubBytesIns_Inst_Sbox_13_T12), .Z(SubBytesIns_Inst_Sbox_13_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T13), .A2(SubBytesIns_Inst_Sbox_13_T6), .ZN(
        SubBytesIns_Inst_Sbox_13_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T23), .A2(SubBytesIns_Inst_Sbox_13_T8), .ZN(
        SubBytesIns_Inst_Sbox_13_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_13_T14), .B(SubBytesIns_Inst_Sbox_13_M1), .Z(SubBytesIns_Inst_Sbox_13_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T19), .A2(ciphertext[104]), .ZN(
        SubBytesIns_Inst_Sbox_13_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_13_M4), 
        .B(SubBytesIns_Inst_Sbox_13_M1), .Z(SubBytesIns_Inst_Sbox_13_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_13_T3), .A2(SubBytesIns_Inst_Sbox_13_T16), .ZN(SubBytesIns_Inst_Sbox_13_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T22), .A2(SubBytesIns_Inst_Sbox_13_T9), .ZN(
        SubBytesIns_Inst_Sbox_13_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_13_T26), .B(SubBytesIns_Inst_Sbox_13_M6), .Z(SubBytesIns_Inst_Sbox_13_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T20), .A2(SubBytesIns_Inst_Sbox_13_T17), .ZN(
        SubBytesIns_Inst_Sbox_13_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_13_M9), .B(SubBytesIns_Inst_Sbox_13_M6), .Z(SubBytesIns_Inst_Sbox_13_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T1), .A2(SubBytesIns_Inst_Sbox_13_T15), .ZN(
        SubBytesIns_Inst_Sbox_13_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T4), .A2(SubBytesIns_Inst_Sbox_13_T27), .ZN(
        SubBytesIns_Inst_Sbox_13_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M12), .B(SubBytesIns_Inst_Sbox_13_M11), .Z(
        SubBytesIns_Inst_Sbox_13_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T2), .A2(SubBytesIns_Inst_Sbox_13_T10), .ZN(
        SubBytesIns_Inst_Sbox_13_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M14), .B(SubBytesIns_Inst_Sbox_13_M11), .Z(
        SubBytesIns_Inst_Sbox_13_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_13_M3), .B(SubBytesIns_Inst_Sbox_13_M2), .Z(SubBytesIns_Inst_Sbox_13_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_13_M5), .B(SubBytesIns_Inst_Sbox_13_T24), .Z(SubBytesIns_Inst_Sbox_13_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_13_M8), .B(SubBytesIns_Inst_Sbox_13_M7), .Z(SubBytesIns_Inst_Sbox_13_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M10), .B(SubBytesIns_Inst_Sbox_13_M15), .Z(
        SubBytesIns_Inst_Sbox_13_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M16), .B(SubBytesIns_Inst_Sbox_13_M13), .Z(
        SubBytesIns_Inst_Sbox_13_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M17), .B(SubBytesIns_Inst_Sbox_13_M15), .Z(
        SubBytesIns_Inst_Sbox_13_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M18), .B(SubBytesIns_Inst_Sbox_13_M13), .Z(
        SubBytesIns_Inst_Sbox_13_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M19), .B(SubBytesIns_Inst_Sbox_13_T25), .Z(
        SubBytesIns_Inst_Sbox_13_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M22), .B(SubBytesIns_Inst_Sbox_13_M23), .Z(
        SubBytesIns_Inst_Sbox_13_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M22), .A2(SubBytesIns_Inst_Sbox_13_M20), .ZN(
        SubBytesIns_Inst_Sbox_13_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M21), .B(SubBytesIns_Inst_Sbox_13_M25), .Z(
        SubBytesIns_Inst_Sbox_13_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M20), .B(SubBytesIns_Inst_Sbox_13_M21), .Z(
        SubBytesIns_Inst_Sbox_13_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M23), .B(SubBytesIns_Inst_Sbox_13_M25), .Z(
        SubBytesIns_Inst_Sbox_13_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M28), .A2(SubBytesIns_Inst_Sbox_13_M27), .ZN(
        SubBytesIns_Inst_Sbox_13_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M26), .A2(SubBytesIns_Inst_Sbox_13_M24), .ZN(
        SubBytesIns_Inst_Sbox_13_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M20), .A2(SubBytesIns_Inst_Sbox_13_M23), .ZN(
        SubBytesIns_Inst_Sbox_13_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M27), .A2(SubBytesIns_Inst_Sbox_13_M31), .ZN(
        SubBytesIns_Inst_Sbox_13_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M27), .B(SubBytesIns_Inst_Sbox_13_M25), .Z(
        SubBytesIns_Inst_Sbox_13_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M21), .A2(SubBytesIns_Inst_Sbox_13_M22), .ZN(
        SubBytesIns_Inst_Sbox_13_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M24), .A2(SubBytesIns_Inst_Sbox_13_M34), .ZN(
        SubBytesIns_Inst_Sbox_13_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M24), .B(SubBytesIns_Inst_Sbox_13_M25), .Z(
        SubBytesIns_Inst_Sbox_13_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M21), .B(SubBytesIns_Inst_Sbox_13_M29), .Z(
        SubBytesIns_Inst_Sbox_13_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M32), .B(SubBytesIns_Inst_Sbox_13_M33), .Z(
        SubBytesIns_Inst_Sbox_13_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M23), .B(SubBytesIns_Inst_Sbox_13_M30), .Z(
        SubBytesIns_Inst_Sbox_13_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M35), .B(SubBytesIns_Inst_Sbox_13_M36), .Z(
        SubBytesIns_Inst_Sbox_13_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M38), .B(SubBytesIns_Inst_Sbox_13_M40), .Z(
        SubBytesIns_Inst_Sbox_13_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M37), .B(SubBytesIns_Inst_Sbox_13_M39), .Z(
        SubBytesIns_Inst_Sbox_13_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M37), .B(SubBytesIns_Inst_Sbox_13_M38), .Z(
        SubBytesIns_Inst_Sbox_13_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M39), .B(SubBytesIns_Inst_Sbox_13_M40), .Z(
        SubBytesIns_Inst_Sbox_13_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M42), .B(SubBytesIns_Inst_Sbox_13_M41), .Z(
        SubBytesIns_Inst_Sbox_13_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M44), .A2(SubBytesIns_Inst_Sbox_13_T6), .ZN(
        SubBytesIns_Inst_Sbox_13_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M40), .A2(SubBytesIns_Inst_Sbox_13_T8), .ZN(
        SubBytesIns_Inst_Sbox_13_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M39), .A2(ciphertext[104]), .ZN(
        SubBytesIns_Inst_Sbox_13_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M43), .A2(SubBytesIns_Inst_Sbox_13_T16), .ZN(
        SubBytesIns_Inst_Sbox_13_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M38), .A2(SubBytesIns_Inst_Sbox_13_T9), .ZN(
        SubBytesIns_Inst_Sbox_13_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M37), .A2(SubBytesIns_Inst_Sbox_13_T17), .ZN(
        SubBytesIns_Inst_Sbox_13_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M42), .A2(SubBytesIns_Inst_Sbox_13_T15), .ZN(
        SubBytesIns_Inst_Sbox_13_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M45), .A2(SubBytesIns_Inst_Sbox_13_T27), .ZN(
        SubBytesIns_Inst_Sbox_13_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M41), .A2(SubBytesIns_Inst_Sbox_13_T10), .ZN(
        SubBytesIns_Inst_Sbox_13_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M44), .A2(SubBytesIns_Inst_Sbox_13_T13), .ZN(
        SubBytesIns_Inst_Sbox_13_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M40), .A2(SubBytesIns_Inst_Sbox_13_T23), .ZN(
        SubBytesIns_Inst_Sbox_13_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M39), .A2(SubBytesIns_Inst_Sbox_13_T19), .ZN(
        SubBytesIns_Inst_Sbox_13_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M43), .A2(SubBytesIns_Inst_Sbox_13_T3), .ZN(
        SubBytesIns_Inst_Sbox_13_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M38), .A2(SubBytesIns_Inst_Sbox_13_T22), .ZN(
        SubBytesIns_Inst_Sbox_13_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M37), .A2(SubBytesIns_Inst_Sbox_13_T20), .ZN(
        SubBytesIns_Inst_Sbox_13_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M42), .A2(SubBytesIns_Inst_Sbox_13_T1), .ZN(
        SubBytesIns_Inst_Sbox_13_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M45), .A2(SubBytesIns_Inst_Sbox_13_T4), .ZN(
        SubBytesIns_Inst_Sbox_13_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M41), .A2(SubBytesIns_Inst_Sbox_13_T2), .ZN(
        SubBytesIns_Inst_Sbox_13_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_13_M61), .B(SubBytesIns_Inst_Sbox_13_M62), .Z(SubBytesIns_Inst_Sbox_13_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_13_M50), .B(SubBytesIns_Inst_Sbox_13_M56), .Z(SubBytesIns_Inst_Sbox_13_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_13_M46), .B(SubBytesIns_Inst_Sbox_13_M48), .Z(SubBytesIns_Inst_Sbox_13_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_13_M47), .B(SubBytesIns_Inst_Sbox_13_M55), .Z(SubBytesIns_Inst_Sbox_13_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_13_M54), .B(SubBytesIns_Inst_Sbox_13_M58), .Z(SubBytesIns_Inst_Sbox_13_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_13_M49), .B(SubBytesIns_Inst_Sbox_13_M61), .Z(SubBytesIns_Inst_Sbox_13_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_13_M62), .B(SubBytesIns_Inst_Sbox_13_L5), .Z(SubBytesIns_Inst_Sbox_13_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_13_M46), .B(SubBytesIns_Inst_Sbox_13_L3), .Z(SubBytesIns_Inst_Sbox_13_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_13_M51), .B(SubBytesIns_Inst_Sbox_13_M59), .Z(SubBytesIns_Inst_Sbox_13_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_13_M52), .B(SubBytesIns_Inst_Sbox_13_M53), .Z(SubBytesIns_Inst_Sbox_13_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M53), .B(SubBytesIns_Inst_Sbox_13_L4), .Z(
        SubBytesIns_Inst_Sbox_13_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M60), .B(SubBytesIns_Inst_Sbox_13_L2), .Z(
        SubBytesIns_Inst_Sbox_13_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M48), .B(SubBytesIns_Inst_Sbox_13_M51), .Z(
        SubBytesIns_Inst_Sbox_13_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M50), .B(SubBytesIns_Inst_Sbox_13_L0), .Z(
        SubBytesIns_Inst_Sbox_13_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M52), .B(SubBytesIns_Inst_Sbox_13_M61), .Z(
        SubBytesIns_Inst_Sbox_13_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M55), .B(SubBytesIns_Inst_Sbox_13_L1), .Z(
        SubBytesIns_Inst_Sbox_13_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M56), .B(SubBytesIns_Inst_Sbox_13_L0), .Z(
        SubBytesIns_Inst_Sbox_13_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M57), .B(SubBytesIns_Inst_Sbox_13_L1), .Z(
        SubBytesIns_Inst_Sbox_13_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M58), .B(SubBytesIns_Inst_Sbox_13_L8), .Z(
        SubBytesIns_Inst_Sbox_13_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M63), .B(SubBytesIns_Inst_Sbox_13_L4), .Z(
        SubBytesIns_Inst_Sbox_13_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_13_L0), .B(SubBytesIns_Inst_Sbox_13_L1), .Z(SubBytesIns_Inst_Sbox_13_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_13_L1), .B(SubBytesIns_Inst_Sbox_13_L7), .Z(SubBytesIns_Inst_Sbox_13_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_13_L3), .B(SubBytesIns_Inst_Sbox_13_L12), .Z(SubBytesIns_Inst_Sbox_13_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L18), .B(SubBytesIns_Inst_Sbox_13_L2), .Z(
        SubBytesIns_Inst_Sbox_13_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L15), .B(SubBytesIns_Inst_Sbox_13_L9), .Z(
        SubBytesIns_Inst_Sbox_13_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_13_L6), .B(SubBytesIns_Inst_Sbox_13_L10), .Z(SubBytesIns_Inst_Sbox_13_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_13_L7), .B(SubBytesIns_Inst_Sbox_13_L9), .Z(SubBytesIns_Inst_Sbox_13_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_13_L8), .B(SubBytesIns_Inst_Sbox_13_L10), .Z(SubBytesIns_Inst_Sbox_13_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L11), .B(SubBytesIns_Inst_Sbox_13_L14), .Z(
        SubBytesIns_Inst_Sbox_13_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L11), .B(SubBytesIns_Inst_Sbox_13_L17), .Z(
        SubBytesIns_Inst_Sbox_13_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_13_L6), 
        .B(SubBytesIns_Inst_Sbox_13_L24), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L16), .B(SubBytesIns_Inst_Sbox_13_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L19), .B(SubBytesIns_Inst_Sbox_13_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_13_L6), 
        .B(SubBytesIns_Inst_Sbox_13_L21), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_13_L20), .B(SubBytesIns_Inst_Sbox_13_L22), .Z(MixColumnsInput[43]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_13_L25), .B(SubBytesIns_Inst_Sbox_13_L29), .Z(MixColumnsInput[42]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L13), .B(SubBytesIns_Inst_Sbox_13_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_13_L6), .B(SubBytesIns_Inst_Sbox_13_L23), .ZN(MixColumnsInput[40]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T1_U1 ( .A(ciphertext[119]), .B(
        ciphertext[116]), .Z(SubBytesIns_Inst_Sbox_14_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T2_U1 ( .A(ciphertext[119]), .B(
        ciphertext[114]), .Z(SubBytesIns_Inst_Sbox_14_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T3_U1 ( .A(ciphertext[119]), .B(
        ciphertext[113]), .Z(SubBytesIns_Inst_Sbox_14_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T4_U1 ( .A(ciphertext[116]), .B(
        ciphertext[114]), .Z(SubBytesIns_Inst_Sbox_14_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T5_U1 ( .A(ciphertext[115]), .B(
        ciphertext[113]), .Z(SubBytesIns_Inst_Sbox_14_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_14_T1), 
        .B(SubBytesIns_Inst_Sbox_14_T5), .Z(SubBytesIns_Inst_Sbox_14_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T7_U1 ( .A(ciphertext[118]), .B(
        ciphertext[117]), .Z(SubBytesIns_Inst_Sbox_14_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T8_U1 ( .A(ciphertext[112]), .B(
        SubBytesIns_Inst_Sbox_14_T6), .Z(SubBytesIns_Inst_Sbox_14_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T9_U1 ( .A(ciphertext[112]), .B(
        SubBytesIns_Inst_Sbox_14_T7), .Z(SubBytesIns_Inst_Sbox_14_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_14_T6), .B(SubBytesIns_Inst_Sbox_14_T7), .Z(SubBytesIns_Inst_Sbox_14_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T11_U1 ( .A(ciphertext[118]), .B(
        ciphertext[114]), .Z(SubBytesIns_Inst_Sbox_14_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T12_U1 ( .A(ciphertext[117]), .B(
        ciphertext[114]), .Z(SubBytesIns_Inst_Sbox_14_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_14_T3), .B(SubBytesIns_Inst_Sbox_14_T4), .Z(SubBytesIns_Inst_Sbox_14_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_14_T6), .B(SubBytesIns_Inst_Sbox_14_T11), .Z(SubBytesIns_Inst_Sbox_14_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_14_T5), .B(SubBytesIns_Inst_Sbox_14_T11), .Z(SubBytesIns_Inst_Sbox_14_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_14_T5), .B(SubBytesIns_Inst_Sbox_14_T12), .Z(SubBytesIns_Inst_Sbox_14_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_14_T9), .B(SubBytesIns_Inst_Sbox_14_T16), .Z(SubBytesIns_Inst_Sbox_14_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T18_U1 ( .A(ciphertext[116]), .B(
        ciphertext[112]), .Z(SubBytesIns_Inst_Sbox_14_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_14_T7), .B(SubBytesIns_Inst_Sbox_14_T18), .Z(SubBytesIns_Inst_Sbox_14_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_14_T1), .B(SubBytesIns_Inst_Sbox_14_T19), .Z(SubBytesIns_Inst_Sbox_14_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T21_U1 ( .A(ciphertext[113]), .B(
        ciphertext[112]), .Z(SubBytesIns_Inst_Sbox_14_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_14_T7), .B(SubBytesIns_Inst_Sbox_14_T21), .Z(SubBytesIns_Inst_Sbox_14_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_14_T2), .B(SubBytesIns_Inst_Sbox_14_T22), .Z(SubBytesIns_Inst_Sbox_14_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_14_T2), .B(SubBytesIns_Inst_Sbox_14_T10), .Z(SubBytesIns_Inst_Sbox_14_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_T20), .B(SubBytesIns_Inst_Sbox_14_T17), .Z(
        SubBytesIns_Inst_Sbox_14_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_14_T3), .B(SubBytesIns_Inst_Sbox_14_T16), .Z(SubBytesIns_Inst_Sbox_14_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_14_T1), .B(SubBytesIns_Inst_Sbox_14_T12), .Z(SubBytesIns_Inst_Sbox_14_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T13), .A2(SubBytesIns_Inst_Sbox_14_T6), .ZN(
        SubBytesIns_Inst_Sbox_14_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T23), .A2(SubBytesIns_Inst_Sbox_14_T8), .ZN(
        SubBytesIns_Inst_Sbox_14_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_14_T14), .B(SubBytesIns_Inst_Sbox_14_M1), .Z(SubBytesIns_Inst_Sbox_14_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T19), .A2(ciphertext[112]), .ZN(
        SubBytesIns_Inst_Sbox_14_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_14_M4), 
        .B(SubBytesIns_Inst_Sbox_14_M1), .Z(SubBytesIns_Inst_Sbox_14_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_14_T3), .A2(SubBytesIns_Inst_Sbox_14_T16), .ZN(SubBytesIns_Inst_Sbox_14_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T22), .A2(SubBytesIns_Inst_Sbox_14_T9), .ZN(
        SubBytesIns_Inst_Sbox_14_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_14_T26), .B(SubBytesIns_Inst_Sbox_14_M6), .Z(SubBytesIns_Inst_Sbox_14_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T20), .A2(SubBytesIns_Inst_Sbox_14_T17), .ZN(
        SubBytesIns_Inst_Sbox_14_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_14_M9), .B(SubBytesIns_Inst_Sbox_14_M6), .Z(SubBytesIns_Inst_Sbox_14_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T1), .A2(SubBytesIns_Inst_Sbox_14_T15), .ZN(
        SubBytesIns_Inst_Sbox_14_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T4), .A2(SubBytesIns_Inst_Sbox_14_T27), .ZN(
        SubBytesIns_Inst_Sbox_14_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M12), .B(SubBytesIns_Inst_Sbox_14_M11), .Z(
        SubBytesIns_Inst_Sbox_14_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T2), .A2(SubBytesIns_Inst_Sbox_14_T10), .ZN(
        SubBytesIns_Inst_Sbox_14_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M14), .B(SubBytesIns_Inst_Sbox_14_M11), .Z(
        SubBytesIns_Inst_Sbox_14_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_14_M3), .B(SubBytesIns_Inst_Sbox_14_M2), .Z(SubBytesIns_Inst_Sbox_14_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_14_M5), .B(SubBytesIns_Inst_Sbox_14_T24), .Z(SubBytesIns_Inst_Sbox_14_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_14_M8), .B(SubBytesIns_Inst_Sbox_14_M7), .Z(SubBytesIns_Inst_Sbox_14_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M10), .B(SubBytesIns_Inst_Sbox_14_M15), .Z(
        SubBytesIns_Inst_Sbox_14_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M16), .B(SubBytesIns_Inst_Sbox_14_M13), .Z(
        SubBytesIns_Inst_Sbox_14_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M17), .B(SubBytesIns_Inst_Sbox_14_M15), .Z(
        SubBytesIns_Inst_Sbox_14_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M18), .B(SubBytesIns_Inst_Sbox_14_M13), .Z(
        SubBytesIns_Inst_Sbox_14_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M19), .B(SubBytesIns_Inst_Sbox_14_T25), .Z(
        SubBytesIns_Inst_Sbox_14_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M22), .B(SubBytesIns_Inst_Sbox_14_M23), .Z(
        SubBytesIns_Inst_Sbox_14_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M22), .A2(SubBytesIns_Inst_Sbox_14_M20), .ZN(
        SubBytesIns_Inst_Sbox_14_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M21), .B(SubBytesIns_Inst_Sbox_14_M25), .Z(
        SubBytesIns_Inst_Sbox_14_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M20), .B(SubBytesIns_Inst_Sbox_14_M21), .Z(
        SubBytesIns_Inst_Sbox_14_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M23), .B(SubBytesIns_Inst_Sbox_14_M25), .Z(
        SubBytesIns_Inst_Sbox_14_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M28), .A2(SubBytesIns_Inst_Sbox_14_M27), .ZN(
        SubBytesIns_Inst_Sbox_14_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M26), .A2(SubBytesIns_Inst_Sbox_14_M24), .ZN(
        SubBytesIns_Inst_Sbox_14_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M20), .A2(SubBytesIns_Inst_Sbox_14_M23), .ZN(
        SubBytesIns_Inst_Sbox_14_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M27), .A2(SubBytesIns_Inst_Sbox_14_M31), .ZN(
        SubBytesIns_Inst_Sbox_14_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M27), .B(SubBytesIns_Inst_Sbox_14_M25), .Z(
        SubBytesIns_Inst_Sbox_14_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M21), .A2(SubBytesIns_Inst_Sbox_14_M22), .ZN(
        SubBytesIns_Inst_Sbox_14_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M24), .A2(SubBytesIns_Inst_Sbox_14_M34), .ZN(
        SubBytesIns_Inst_Sbox_14_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M24), .B(SubBytesIns_Inst_Sbox_14_M25), .Z(
        SubBytesIns_Inst_Sbox_14_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M21), .B(SubBytesIns_Inst_Sbox_14_M29), .Z(
        SubBytesIns_Inst_Sbox_14_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M32), .B(SubBytesIns_Inst_Sbox_14_M33), .Z(
        SubBytesIns_Inst_Sbox_14_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M23), .B(SubBytesIns_Inst_Sbox_14_M30), .Z(
        SubBytesIns_Inst_Sbox_14_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M35), .B(SubBytesIns_Inst_Sbox_14_M36), .Z(
        SubBytesIns_Inst_Sbox_14_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M38), .B(SubBytesIns_Inst_Sbox_14_M40), .Z(
        SubBytesIns_Inst_Sbox_14_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M37), .B(SubBytesIns_Inst_Sbox_14_M39), .Z(
        SubBytesIns_Inst_Sbox_14_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M37), .B(SubBytesIns_Inst_Sbox_14_M38), .Z(
        SubBytesIns_Inst_Sbox_14_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M39), .B(SubBytesIns_Inst_Sbox_14_M40), .Z(
        SubBytesIns_Inst_Sbox_14_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M42), .B(SubBytesIns_Inst_Sbox_14_M41), .Z(
        SubBytesIns_Inst_Sbox_14_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M44), .A2(SubBytesIns_Inst_Sbox_14_T6), .ZN(
        SubBytesIns_Inst_Sbox_14_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M40), .A2(SubBytesIns_Inst_Sbox_14_T8), .ZN(
        SubBytesIns_Inst_Sbox_14_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M39), .A2(ciphertext[112]), .ZN(
        SubBytesIns_Inst_Sbox_14_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M43), .A2(SubBytesIns_Inst_Sbox_14_T16), .ZN(
        SubBytesIns_Inst_Sbox_14_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M38), .A2(SubBytesIns_Inst_Sbox_14_T9), .ZN(
        SubBytesIns_Inst_Sbox_14_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M37), .A2(SubBytesIns_Inst_Sbox_14_T17), .ZN(
        SubBytesIns_Inst_Sbox_14_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M42), .A2(SubBytesIns_Inst_Sbox_14_T15), .ZN(
        SubBytesIns_Inst_Sbox_14_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M45), .A2(SubBytesIns_Inst_Sbox_14_T27), .ZN(
        SubBytesIns_Inst_Sbox_14_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M41), .A2(SubBytesIns_Inst_Sbox_14_T10), .ZN(
        SubBytesIns_Inst_Sbox_14_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M44), .A2(SubBytesIns_Inst_Sbox_14_T13), .ZN(
        SubBytesIns_Inst_Sbox_14_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M40), .A2(SubBytesIns_Inst_Sbox_14_T23), .ZN(
        SubBytesIns_Inst_Sbox_14_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M39), .A2(SubBytesIns_Inst_Sbox_14_T19), .ZN(
        SubBytesIns_Inst_Sbox_14_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M43), .A2(SubBytesIns_Inst_Sbox_14_T3), .ZN(
        SubBytesIns_Inst_Sbox_14_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M38), .A2(SubBytesIns_Inst_Sbox_14_T22), .ZN(
        SubBytesIns_Inst_Sbox_14_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M37), .A2(SubBytesIns_Inst_Sbox_14_T20), .ZN(
        SubBytesIns_Inst_Sbox_14_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M42), .A2(SubBytesIns_Inst_Sbox_14_T1), .ZN(
        SubBytesIns_Inst_Sbox_14_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M45), .A2(SubBytesIns_Inst_Sbox_14_T4), .ZN(
        SubBytesIns_Inst_Sbox_14_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M41), .A2(SubBytesIns_Inst_Sbox_14_T2), .ZN(
        SubBytesIns_Inst_Sbox_14_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_14_M61), .B(SubBytesIns_Inst_Sbox_14_M62), .Z(SubBytesIns_Inst_Sbox_14_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_14_M50), .B(SubBytesIns_Inst_Sbox_14_M56), .Z(SubBytesIns_Inst_Sbox_14_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_14_M46), .B(SubBytesIns_Inst_Sbox_14_M48), .Z(SubBytesIns_Inst_Sbox_14_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_14_M47), .B(SubBytesIns_Inst_Sbox_14_M55), .Z(SubBytesIns_Inst_Sbox_14_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_14_M54), .B(SubBytesIns_Inst_Sbox_14_M58), .Z(SubBytesIns_Inst_Sbox_14_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_14_M49), .B(SubBytesIns_Inst_Sbox_14_M61), .Z(SubBytesIns_Inst_Sbox_14_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_14_M62), .B(SubBytesIns_Inst_Sbox_14_L5), .Z(SubBytesIns_Inst_Sbox_14_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_14_M46), .B(SubBytesIns_Inst_Sbox_14_L3), .Z(SubBytesIns_Inst_Sbox_14_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_14_M51), .B(SubBytesIns_Inst_Sbox_14_M59), .Z(SubBytesIns_Inst_Sbox_14_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_14_M52), .B(SubBytesIns_Inst_Sbox_14_M53), .Z(SubBytesIns_Inst_Sbox_14_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M53), .B(SubBytesIns_Inst_Sbox_14_L4), .Z(
        SubBytesIns_Inst_Sbox_14_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M60), .B(SubBytesIns_Inst_Sbox_14_L2), .Z(
        SubBytesIns_Inst_Sbox_14_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M48), .B(SubBytesIns_Inst_Sbox_14_M51), .Z(
        SubBytesIns_Inst_Sbox_14_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M50), .B(SubBytesIns_Inst_Sbox_14_L0), .Z(
        SubBytesIns_Inst_Sbox_14_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M52), .B(SubBytesIns_Inst_Sbox_14_M61), .Z(
        SubBytesIns_Inst_Sbox_14_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M55), .B(SubBytesIns_Inst_Sbox_14_L1), .Z(
        SubBytesIns_Inst_Sbox_14_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M56), .B(SubBytesIns_Inst_Sbox_14_L0), .Z(
        SubBytesIns_Inst_Sbox_14_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M57), .B(SubBytesIns_Inst_Sbox_14_L1), .Z(
        SubBytesIns_Inst_Sbox_14_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M58), .B(SubBytesIns_Inst_Sbox_14_L8), .Z(
        SubBytesIns_Inst_Sbox_14_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M63), .B(SubBytesIns_Inst_Sbox_14_L4), .Z(
        SubBytesIns_Inst_Sbox_14_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_14_L0), .B(SubBytesIns_Inst_Sbox_14_L1), .Z(SubBytesIns_Inst_Sbox_14_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_14_L1), .B(SubBytesIns_Inst_Sbox_14_L7), .Z(SubBytesIns_Inst_Sbox_14_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_14_L3), .B(SubBytesIns_Inst_Sbox_14_L12), .Z(SubBytesIns_Inst_Sbox_14_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L18), .B(SubBytesIns_Inst_Sbox_14_L2), .Z(
        SubBytesIns_Inst_Sbox_14_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L15), .B(SubBytesIns_Inst_Sbox_14_L9), .Z(
        SubBytesIns_Inst_Sbox_14_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_14_L6), .B(SubBytesIns_Inst_Sbox_14_L10), .Z(SubBytesIns_Inst_Sbox_14_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_14_L7), .B(SubBytesIns_Inst_Sbox_14_L9), .Z(SubBytesIns_Inst_Sbox_14_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_14_L8), .B(SubBytesIns_Inst_Sbox_14_L10), .Z(SubBytesIns_Inst_Sbox_14_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L11), .B(SubBytesIns_Inst_Sbox_14_L14), .Z(
        SubBytesIns_Inst_Sbox_14_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L11), .B(SubBytesIns_Inst_Sbox_14_L17), .Z(
        SubBytesIns_Inst_Sbox_14_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_14_L6), 
        .B(SubBytesIns_Inst_Sbox_14_L24), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L16), .B(SubBytesIns_Inst_Sbox_14_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L19), .B(SubBytesIns_Inst_Sbox_14_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_14_L6), 
        .B(SubBytesIns_Inst_Sbox_14_L21), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_14_L20), .B(SubBytesIns_Inst_Sbox_14_L22), .Z(MixColumnsInput[19]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_14_L25), .B(SubBytesIns_Inst_Sbox_14_L29), .Z(MixColumnsInput[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L13), .B(SubBytesIns_Inst_Sbox_14_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_14_L6), .B(SubBytesIns_Inst_Sbox_14_L23), .ZN(MixColumnsInput[16]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T1_U1 ( .A(ciphertext[127]), .B(
        ciphertext[124]), .Z(SubBytesIns_Inst_Sbox_15_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T2_U1 ( .A(ciphertext[127]), .B(
        ciphertext[122]), .Z(SubBytesIns_Inst_Sbox_15_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T3_U1 ( .A(ciphertext[127]), .B(
        ciphertext[121]), .Z(SubBytesIns_Inst_Sbox_15_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T4_U1 ( .A(ciphertext[124]), .B(
        ciphertext[122]), .Z(SubBytesIns_Inst_Sbox_15_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T5_U1 ( .A(ciphertext[123]), .B(
        ciphertext[121]), .Z(SubBytesIns_Inst_Sbox_15_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_15_T1), 
        .B(SubBytesIns_Inst_Sbox_15_T5), .Z(SubBytesIns_Inst_Sbox_15_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T7_U1 ( .A(ciphertext[126]), .B(
        ciphertext[125]), .Z(SubBytesIns_Inst_Sbox_15_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T8_U1 ( .A(ciphertext[120]), .B(
        SubBytesIns_Inst_Sbox_15_T6), .Z(SubBytesIns_Inst_Sbox_15_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T9_U1 ( .A(ciphertext[120]), .B(
        SubBytesIns_Inst_Sbox_15_T7), .Z(SubBytesIns_Inst_Sbox_15_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_15_T6), .B(SubBytesIns_Inst_Sbox_15_T7), .Z(SubBytesIns_Inst_Sbox_15_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T11_U1 ( .A(ciphertext[126]), .B(
        ciphertext[122]), .Z(SubBytesIns_Inst_Sbox_15_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T12_U1 ( .A(ciphertext[125]), .B(
        ciphertext[122]), .Z(SubBytesIns_Inst_Sbox_15_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_15_T3), .B(SubBytesIns_Inst_Sbox_15_T4), .Z(SubBytesIns_Inst_Sbox_15_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_15_T6), .B(SubBytesIns_Inst_Sbox_15_T11), .Z(SubBytesIns_Inst_Sbox_15_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_15_T5), .B(SubBytesIns_Inst_Sbox_15_T11), .Z(SubBytesIns_Inst_Sbox_15_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_15_T5), .B(SubBytesIns_Inst_Sbox_15_T12), .Z(SubBytesIns_Inst_Sbox_15_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_15_T9), .B(SubBytesIns_Inst_Sbox_15_T16), .Z(SubBytesIns_Inst_Sbox_15_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T18_U1 ( .A(ciphertext[124]), .B(
        ciphertext[120]), .Z(SubBytesIns_Inst_Sbox_15_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_15_T7), .B(SubBytesIns_Inst_Sbox_15_T18), .Z(SubBytesIns_Inst_Sbox_15_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_15_T1), .B(SubBytesIns_Inst_Sbox_15_T19), .Z(SubBytesIns_Inst_Sbox_15_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T21_U1 ( .A(ciphertext[121]), .B(
        ciphertext[120]), .Z(SubBytesIns_Inst_Sbox_15_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_15_T7), .B(SubBytesIns_Inst_Sbox_15_T21), .Z(SubBytesIns_Inst_Sbox_15_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_15_T2), .B(SubBytesIns_Inst_Sbox_15_T22), .Z(SubBytesIns_Inst_Sbox_15_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_15_T2), .B(SubBytesIns_Inst_Sbox_15_T10), .Z(SubBytesIns_Inst_Sbox_15_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_T20), .B(SubBytesIns_Inst_Sbox_15_T17), .Z(
        SubBytesIns_Inst_Sbox_15_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_15_T3), .B(SubBytesIns_Inst_Sbox_15_T16), .Z(SubBytesIns_Inst_Sbox_15_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_15_T1), .B(SubBytesIns_Inst_Sbox_15_T12), .Z(SubBytesIns_Inst_Sbox_15_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T13), .A2(SubBytesIns_Inst_Sbox_15_T6), .ZN(
        SubBytesIns_Inst_Sbox_15_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T23), .A2(SubBytesIns_Inst_Sbox_15_T8), .ZN(
        SubBytesIns_Inst_Sbox_15_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_15_T14), .B(SubBytesIns_Inst_Sbox_15_M1), .Z(SubBytesIns_Inst_Sbox_15_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T19), .A2(ciphertext[120]), .ZN(
        SubBytesIns_Inst_Sbox_15_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_15_M4), 
        .B(SubBytesIns_Inst_Sbox_15_M1), .Z(SubBytesIns_Inst_Sbox_15_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_15_T3), .A2(SubBytesIns_Inst_Sbox_15_T16), .ZN(SubBytesIns_Inst_Sbox_15_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T22), .A2(SubBytesIns_Inst_Sbox_15_T9), .ZN(
        SubBytesIns_Inst_Sbox_15_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_15_T26), .B(SubBytesIns_Inst_Sbox_15_M6), .Z(SubBytesIns_Inst_Sbox_15_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T20), .A2(SubBytesIns_Inst_Sbox_15_T17), .ZN(
        SubBytesIns_Inst_Sbox_15_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_15_M9), .B(SubBytesIns_Inst_Sbox_15_M6), .Z(SubBytesIns_Inst_Sbox_15_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T1), .A2(SubBytesIns_Inst_Sbox_15_T15), .ZN(
        SubBytesIns_Inst_Sbox_15_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T4), .A2(SubBytesIns_Inst_Sbox_15_T27), .ZN(
        SubBytesIns_Inst_Sbox_15_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M12), .B(SubBytesIns_Inst_Sbox_15_M11), .Z(
        SubBytesIns_Inst_Sbox_15_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T2), .A2(SubBytesIns_Inst_Sbox_15_T10), .ZN(
        SubBytesIns_Inst_Sbox_15_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M14), .B(SubBytesIns_Inst_Sbox_15_M11), .Z(
        SubBytesIns_Inst_Sbox_15_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_15_M3), .B(SubBytesIns_Inst_Sbox_15_M2), .Z(SubBytesIns_Inst_Sbox_15_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_15_M5), .B(SubBytesIns_Inst_Sbox_15_T24), .Z(SubBytesIns_Inst_Sbox_15_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_15_M8), .B(SubBytesIns_Inst_Sbox_15_M7), .Z(SubBytesIns_Inst_Sbox_15_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M10), .B(SubBytesIns_Inst_Sbox_15_M15), .Z(
        SubBytesIns_Inst_Sbox_15_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M16), .B(SubBytesIns_Inst_Sbox_15_M13), .Z(
        SubBytesIns_Inst_Sbox_15_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M17), .B(SubBytesIns_Inst_Sbox_15_M15), .Z(
        SubBytesIns_Inst_Sbox_15_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M18), .B(SubBytesIns_Inst_Sbox_15_M13), .Z(
        SubBytesIns_Inst_Sbox_15_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M19), .B(SubBytesIns_Inst_Sbox_15_T25), .Z(
        SubBytesIns_Inst_Sbox_15_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M22), .B(SubBytesIns_Inst_Sbox_15_M23), .Z(
        SubBytesIns_Inst_Sbox_15_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M22), .A2(SubBytesIns_Inst_Sbox_15_M20), .ZN(
        SubBytesIns_Inst_Sbox_15_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M21), .B(SubBytesIns_Inst_Sbox_15_M25), .Z(
        SubBytesIns_Inst_Sbox_15_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M20), .B(SubBytesIns_Inst_Sbox_15_M21), .Z(
        SubBytesIns_Inst_Sbox_15_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M23), .B(SubBytesIns_Inst_Sbox_15_M25), .Z(
        SubBytesIns_Inst_Sbox_15_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M28), .A2(SubBytesIns_Inst_Sbox_15_M27), .ZN(
        SubBytesIns_Inst_Sbox_15_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M26), .A2(SubBytesIns_Inst_Sbox_15_M24), .ZN(
        SubBytesIns_Inst_Sbox_15_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M20), .A2(SubBytesIns_Inst_Sbox_15_M23), .ZN(
        SubBytesIns_Inst_Sbox_15_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M27), .A2(SubBytesIns_Inst_Sbox_15_M31), .ZN(
        SubBytesIns_Inst_Sbox_15_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M27), .B(SubBytesIns_Inst_Sbox_15_M25), .Z(
        SubBytesIns_Inst_Sbox_15_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M21), .A2(SubBytesIns_Inst_Sbox_15_M22), .ZN(
        SubBytesIns_Inst_Sbox_15_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M24), .A2(SubBytesIns_Inst_Sbox_15_M34), .ZN(
        SubBytesIns_Inst_Sbox_15_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M24), .B(SubBytesIns_Inst_Sbox_15_M25), .Z(
        SubBytesIns_Inst_Sbox_15_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M21), .B(SubBytesIns_Inst_Sbox_15_M29), .Z(
        SubBytesIns_Inst_Sbox_15_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M32), .B(SubBytesIns_Inst_Sbox_15_M33), .Z(
        SubBytesIns_Inst_Sbox_15_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M23), .B(SubBytesIns_Inst_Sbox_15_M30), .Z(
        SubBytesIns_Inst_Sbox_15_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M35), .B(SubBytesIns_Inst_Sbox_15_M36), .Z(
        SubBytesIns_Inst_Sbox_15_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M38), .B(SubBytesIns_Inst_Sbox_15_M40), .Z(
        SubBytesIns_Inst_Sbox_15_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M37), .B(SubBytesIns_Inst_Sbox_15_M39), .Z(
        SubBytesIns_Inst_Sbox_15_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M37), .B(SubBytesIns_Inst_Sbox_15_M38), .Z(
        SubBytesIns_Inst_Sbox_15_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M39), .B(SubBytesIns_Inst_Sbox_15_M40), .Z(
        SubBytesIns_Inst_Sbox_15_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M42), .B(SubBytesIns_Inst_Sbox_15_M41), .Z(
        SubBytesIns_Inst_Sbox_15_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M44), .A2(SubBytesIns_Inst_Sbox_15_T6), .ZN(
        SubBytesIns_Inst_Sbox_15_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M40), .A2(SubBytesIns_Inst_Sbox_15_T8), .ZN(
        SubBytesIns_Inst_Sbox_15_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M39), .A2(ciphertext[120]), .ZN(
        SubBytesIns_Inst_Sbox_15_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M43), .A2(SubBytesIns_Inst_Sbox_15_T16), .ZN(
        SubBytesIns_Inst_Sbox_15_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M38), .A2(SubBytesIns_Inst_Sbox_15_T9), .ZN(
        SubBytesIns_Inst_Sbox_15_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M37), .A2(SubBytesIns_Inst_Sbox_15_T17), .ZN(
        SubBytesIns_Inst_Sbox_15_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M42), .A2(SubBytesIns_Inst_Sbox_15_T15), .ZN(
        SubBytesIns_Inst_Sbox_15_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M45), .A2(SubBytesIns_Inst_Sbox_15_T27), .ZN(
        SubBytesIns_Inst_Sbox_15_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M41), .A2(SubBytesIns_Inst_Sbox_15_T10), .ZN(
        SubBytesIns_Inst_Sbox_15_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M44), .A2(SubBytesIns_Inst_Sbox_15_T13), .ZN(
        SubBytesIns_Inst_Sbox_15_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M40), .A2(SubBytesIns_Inst_Sbox_15_T23), .ZN(
        SubBytesIns_Inst_Sbox_15_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M39), .A2(SubBytesIns_Inst_Sbox_15_T19), .ZN(
        SubBytesIns_Inst_Sbox_15_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M43), .A2(SubBytesIns_Inst_Sbox_15_T3), .ZN(
        SubBytesIns_Inst_Sbox_15_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M38), .A2(SubBytesIns_Inst_Sbox_15_T22), .ZN(
        SubBytesIns_Inst_Sbox_15_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M37), .A2(SubBytesIns_Inst_Sbox_15_T20), .ZN(
        SubBytesIns_Inst_Sbox_15_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M42), .A2(SubBytesIns_Inst_Sbox_15_T1), .ZN(
        SubBytesIns_Inst_Sbox_15_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M45), .A2(SubBytesIns_Inst_Sbox_15_T4), .ZN(
        SubBytesIns_Inst_Sbox_15_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M41), .A2(SubBytesIns_Inst_Sbox_15_T2), .ZN(
        SubBytesIns_Inst_Sbox_15_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_15_M61), .B(SubBytesIns_Inst_Sbox_15_M62), .Z(SubBytesIns_Inst_Sbox_15_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_15_M50), .B(SubBytesIns_Inst_Sbox_15_M56), .Z(SubBytesIns_Inst_Sbox_15_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_15_M46), .B(SubBytesIns_Inst_Sbox_15_M48), .Z(SubBytesIns_Inst_Sbox_15_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_15_M47), .B(SubBytesIns_Inst_Sbox_15_M55), .Z(SubBytesIns_Inst_Sbox_15_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_15_M54), .B(SubBytesIns_Inst_Sbox_15_M58), .Z(SubBytesIns_Inst_Sbox_15_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_15_M49), .B(SubBytesIns_Inst_Sbox_15_M61), .Z(SubBytesIns_Inst_Sbox_15_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_15_M62), .B(SubBytesIns_Inst_Sbox_15_L5), .Z(SubBytesIns_Inst_Sbox_15_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_15_M46), .B(SubBytesIns_Inst_Sbox_15_L3), .Z(SubBytesIns_Inst_Sbox_15_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_15_M51), .B(SubBytesIns_Inst_Sbox_15_M59), .Z(SubBytesIns_Inst_Sbox_15_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_15_M52), .B(SubBytesIns_Inst_Sbox_15_M53), .Z(SubBytesIns_Inst_Sbox_15_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M53), .B(SubBytesIns_Inst_Sbox_15_L4), .Z(
        SubBytesIns_Inst_Sbox_15_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M60), .B(SubBytesIns_Inst_Sbox_15_L2), .Z(
        SubBytesIns_Inst_Sbox_15_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M48), .B(SubBytesIns_Inst_Sbox_15_M51), .Z(
        SubBytesIns_Inst_Sbox_15_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M50), .B(SubBytesIns_Inst_Sbox_15_L0), .Z(
        SubBytesIns_Inst_Sbox_15_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M52), .B(SubBytesIns_Inst_Sbox_15_M61), .Z(
        SubBytesIns_Inst_Sbox_15_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M55), .B(SubBytesIns_Inst_Sbox_15_L1), .Z(
        SubBytesIns_Inst_Sbox_15_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M56), .B(SubBytesIns_Inst_Sbox_15_L0), .Z(
        SubBytesIns_Inst_Sbox_15_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M57), .B(SubBytesIns_Inst_Sbox_15_L1), .Z(
        SubBytesIns_Inst_Sbox_15_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M58), .B(SubBytesIns_Inst_Sbox_15_L8), .Z(
        SubBytesIns_Inst_Sbox_15_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M63), .B(SubBytesIns_Inst_Sbox_15_L4), .Z(
        SubBytesIns_Inst_Sbox_15_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_15_L0), .B(SubBytesIns_Inst_Sbox_15_L1), .Z(SubBytesIns_Inst_Sbox_15_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_15_L1), .B(SubBytesIns_Inst_Sbox_15_L7), .Z(SubBytesIns_Inst_Sbox_15_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_15_L3), .B(SubBytesIns_Inst_Sbox_15_L12), .Z(SubBytesIns_Inst_Sbox_15_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L18), .B(SubBytesIns_Inst_Sbox_15_L2), .Z(
        SubBytesIns_Inst_Sbox_15_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L15), .B(SubBytesIns_Inst_Sbox_15_L9), .Z(
        SubBytesIns_Inst_Sbox_15_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_15_L6), .B(SubBytesIns_Inst_Sbox_15_L10), .Z(SubBytesIns_Inst_Sbox_15_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_15_L7), .B(SubBytesIns_Inst_Sbox_15_L9), .Z(SubBytesIns_Inst_Sbox_15_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_15_L8), .B(SubBytesIns_Inst_Sbox_15_L10), .Z(SubBytesIns_Inst_Sbox_15_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L11), .B(SubBytesIns_Inst_Sbox_15_L14), .Z(
        SubBytesIns_Inst_Sbox_15_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L11), .B(SubBytesIns_Inst_Sbox_15_L17), .Z(
        SubBytesIns_Inst_Sbox_15_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_15_L6), 
        .B(SubBytesIns_Inst_Sbox_15_L24), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L16), .B(SubBytesIns_Inst_Sbox_15_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L19), .B(SubBytesIns_Inst_Sbox_15_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_15_L6), 
        .B(SubBytesIns_Inst_Sbox_15_L21), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_15_L20), .B(SubBytesIns_Inst_Sbox_15_L22), .Z(MixColumnsInput[123]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_15_L25), .B(SubBytesIns_Inst_Sbox_15_L29), .Z(MixColumnsInput[122]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L13), .B(SubBytesIns_Inst_Sbox_15_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_15_L6), .B(SubBytesIns_Inst_Sbox_15_L23), .ZN(MixColumnsInput[120]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U96 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n64), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .ZN(
        MixColumnsOutput[105]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U95 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n63), .B(
        MixColumnsIns_MixOneColumnInst_0_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n64) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U94 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n61), .B(
        MixColumnsIns_MixOneColumnInst_0_n60), .ZN(MixColumnsOutput[104]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U93 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n59), .B(MixColumnsInput[112]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n61) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U92 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n58), .B(
        MixColumnsIns_MixOneColumnInst_0_n57), .ZN(MixColumnsOutput[103]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U91 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n56), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n58) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U90 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n55), .B(
        MixColumnsIns_MixOneColumnInst_0_n54), .ZN(MixColumnsOutput[102]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U89 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n53), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n55) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U88 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n52), .B(
        MixColumnsIns_MixOneColumnInst_0_n51), .ZN(MixColumnsOutput[101]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U87 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n50), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n52) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U86 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n49), .B(
        MixColumnsIns_MixOneColumnInst_0_n48), .ZN(MixColumnsOutput[100]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U85 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n47), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n49) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U84 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n46), .B(
        MixColumnsIns_MixOneColumnInst_0_n45), .ZN(MixColumnsOutput[99]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U83 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n44), .B(MixColumnsInput[107]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n46) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U82 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n43), .B(
        MixColumnsIns_MixOneColumnInst_0_n57), .ZN(MixColumnsOutput[127]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U81 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n57) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U80 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_0_n42), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n43) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U79 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n41), .B(
        MixColumnsIns_MixOneColumnInst_0_n54), .ZN(MixColumnsOutput[126]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U78 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n54) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U77 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_0_n40), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n41) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U76 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n39), .B(
        MixColumnsIns_MixOneColumnInst_0_n38), .ZN(MixColumnsOutput[98]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U75 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n37), .B(MixColumnsInput[106]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n39) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U74 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n36), .B(
        MixColumnsIns_MixOneColumnInst_0_n51), .ZN(MixColumnsOutput[125]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U73 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n51) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U72 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_0_n35), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n36) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U71 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n34), .B(
        MixColumnsIns_MixOneColumnInst_0_n48), .ZN(MixColumnsOutput[124]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U70 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n48) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U69 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_0_n33), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n34) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U68 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n32), .B(
        MixColumnsIns_MixOneColumnInst_0_n45), .ZN(MixColumnsOutput[123]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U67 ( .A(MixColumnsInput[115]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n45) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U66 ( .A(MixColumnsInput[99]), .B(
        MixColumnsIns_MixOneColumnInst_0_n31), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n32) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U65 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n30), .B(
        MixColumnsIns_MixOneColumnInst_0_n38), .ZN(MixColumnsOutput[122]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U64 ( .A(MixColumnsInput[114]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n38) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U63 ( .A(MixColumnsInput[98]), .B(
        MixColumnsIns_MixOneColumnInst_0_n29), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n30) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U62 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n28), .B(
        MixColumnsIns_MixOneColumnInst_0_n27), .ZN(MixColumnsOutput[121]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U61 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .B(
        MixColumnsIns_MixOneColumnInst_0_n26), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n28) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U60 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n25), .B(
        MixColumnsIns_MixOneColumnInst_0_n24), .ZN(MixColumnsOutput[120]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U59 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n23), .B(MixColumnsInput[96]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n25) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U58 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n22), .B(
        MixColumnsIns_MixOneColumnInst_0_n42), .ZN(MixColumnsOutput[119]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U57 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n42) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U56 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B(
        MixColumnsIns_MixOneColumnInst_0_n21), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n22) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U55 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n20), .B(
        MixColumnsIns_MixOneColumnInst_0_n40), .ZN(MixColumnsOutput[118]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U54 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n40) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U53 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .B(
        MixColumnsIns_MixOneColumnInst_0_n19), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n20) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U52 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n18), .B(
        MixColumnsIns_MixOneColumnInst_0_n35), .ZN(MixColumnsOutput[117]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U51 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n35) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U50 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .B(
        MixColumnsIns_MixOneColumnInst_0_n17), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n18) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U49 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n16), .B(
        MixColumnsIns_MixOneColumnInst_0_n33), .ZN(MixColumnsOutput[116]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U48 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n33) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U47 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .B(
        MixColumnsIns_MixOneColumnInst_0_n15), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n16) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U46 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n14), .B(
        MixColumnsIns_MixOneColumnInst_0_n27), .ZN(MixColumnsOutput[97]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U45 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n27) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U44 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .B(
        MixColumnsIns_MixOneColumnInst_0_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n14) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U43 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n62) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U42 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n13), .B(
        MixColumnsIns_MixOneColumnInst_0_n31), .ZN(MixColumnsOutput[115]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U41 ( .A(MixColumnsInput[107]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n31) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U40 ( .A(MixColumnsInput[123]), 
        .B(MixColumnsIns_MixOneColumnInst_0_n12), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n13) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U39 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n11), .B(
        MixColumnsIns_MixOneColumnInst_0_n29), .ZN(MixColumnsOutput[114]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U38 ( .A(MixColumnsInput[106]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n29) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U37 ( .A(MixColumnsInput[122]), 
        .B(MixColumnsIns_MixOneColumnInst_0_n10), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n11) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U36 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n9), .B(
        MixColumnsIns_MixOneColumnInst_0_n26), .ZN(MixColumnsOutput[113]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U35 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n26) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U34 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n63), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n9) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U33 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n63) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U32 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n8), .B(
        MixColumnsIns_MixOneColumnInst_0_n24), .ZN(MixColumnsOutput[112]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U31 ( .A(MixColumnsInput[104]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n24) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U30 ( .A(MixColumnsInput[120]), 
        .B(MixColumnsIns_MixOneColumnInst_0_n60), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n8) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U29 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsInput[96]), .Z(MixColumnsIns_MixOneColumnInst_0_n60) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U28 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n7), .B(
        MixColumnsIns_MixOneColumnInst_0_n21), .ZN(MixColumnsOutput[111]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U27 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n21) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U26 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n56), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n7) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U25 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n56) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U24 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n6), .B(
        MixColumnsIns_MixOneColumnInst_0_n19), .ZN(MixColumnsOutput[110]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U23 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n19) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U22 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n53), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n6) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U21 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n53) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U20 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n5), .B(
        MixColumnsIns_MixOneColumnInst_0_n17), .ZN(MixColumnsOutput[109]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U19 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n17) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U18 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n50), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n5) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U17 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n50) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U16 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n4), .B(
        MixColumnsIns_MixOneColumnInst_0_n15), .ZN(MixColumnsOutput[108]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U15 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n15) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U14 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n47), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n4) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U13 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n47) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U12 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n3), .B(
        MixColumnsIns_MixOneColumnInst_0_n12), .ZN(MixColumnsOutput[107]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U11 ( .A(MixColumnsInput[99]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n12) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U10 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n44), .B(MixColumnsInput[115]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n3) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U9 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]), .B(
        MixColumnsInput[123]), .Z(MixColumnsIns_MixOneColumnInst_0_n44) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U8 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n2), .B(
        MixColumnsIns_MixOneColumnInst_0_n10), .ZN(MixColumnsOutput[106]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U7 ( .A(MixColumnsInput[98]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n10) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U6 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n37), .B(MixColumnsInput[114]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n2) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U5 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .B(
        MixColumnsInput[122]), .Z(MixColumnsIns_MixOneColumnInst_0_n37) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U4 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n1), .B(MixColumnsInput[104]), .ZN(
        MixColumnsOutput[96]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n59), .B(
        MixColumnsIns_MixOneColumnInst_0_n23), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n1) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U2 ( .A(MixColumnsInput[112]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n23) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsInput[120]), .Z(MixColumnsIns_MixOneColumnInst_0_n59) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B(
        MixColumnsInput[123]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B(
        MixColumnsInput[122]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B(
        MixColumnsInput[120]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B(
        MixColumnsInput[115]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B(
        MixColumnsInput[114]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B(
        MixColumnsInput[112]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsInput[107]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsInput[106]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsInput[104]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsInput[99]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsInput[98]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsInput[96]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U96 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n64), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .ZN(
        MixColumnsOutput[73]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U95 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n63), .B(
        MixColumnsIns_MixOneColumnInst_1_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n64) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U94 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n61), .B(
        MixColumnsIns_MixOneColumnInst_1_n60), .ZN(MixColumnsOutput[72]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U93 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n59), .B(MixColumnsInput[80]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n61) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U92 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n58), .B(
        MixColumnsIns_MixOneColumnInst_1_n57), .ZN(MixColumnsOutput[71]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U91 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n56), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n58) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U90 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n55), .B(
        MixColumnsIns_MixOneColumnInst_1_n54), .ZN(MixColumnsOutput[70]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U89 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n53), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n55) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U88 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n52), .B(
        MixColumnsIns_MixOneColumnInst_1_n51), .ZN(MixColumnsOutput[69]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U87 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n50), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n52) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U86 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n49), .B(
        MixColumnsIns_MixOneColumnInst_1_n48), .ZN(MixColumnsOutput[68]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U85 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n47), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n49) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U84 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n46), .B(
        MixColumnsIns_MixOneColumnInst_1_n45), .ZN(MixColumnsOutput[67]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U83 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n44), .B(MixColumnsInput[75]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n46) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U82 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n43), .B(
        MixColumnsIns_MixOneColumnInst_1_n57), .ZN(MixColumnsOutput[95]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U81 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n57) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U80 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_1_n42), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n43) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U79 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n41), .B(
        MixColumnsIns_MixOneColumnInst_1_n54), .ZN(MixColumnsOutput[94]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U78 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n54) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U77 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_1_n40), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n41) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U76 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n39), .B(
        MixColumnsIns_MixOneColumnInst_1_n38), .ZN(MixColumnsOutput[66]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U75 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n37), .B(MixColumnsInput[74]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n39) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U74 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n36), .B(
        MixColumnsIns_MixOneColumnInst_1_n51), .ZN(MixColumnsOutput[93]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U73 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n51) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U72 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_1_n35), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n36) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U71 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n34), .B(
        MixColumnsIns_MixOneColumnInst_1_n48), .ZN(MixColumnsOutput[92]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U70 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n48) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U69 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_1_n33), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n34) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U68 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n32), .B(
        MixColumnsIns_MixOneColumnInst_1_n45), .ZN(MixColumnsOutput[91]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U67 ( .A(MixColumnsInput[83]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n45) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U66 ( .A(MixColumnsInput[67]), .B(
        MixColumnsIns_MixOneColumnInst_1_n31), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n32) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U65 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n30), .B(
        MixColumnsIns_MixOneColumnInst_1_n38), .ZN(MixColumnsOutput[90]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U64 ( .A(MixColumnsInput[82]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n38) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U63 ( .A(MixColumnsInput[66]), .B(
        MixColumnsIns_MixOneColumnInst_1_n29), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n30) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U62 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n28), .B(
        MixColumnsIns_MixOneColumnInst_1_n27), .ZN(MixColumnsOutput[89]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U61 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .B(
        MixColumnsIns_MixOneColumnInst_1_n26), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n28) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U60 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n25), .B(
        MixColumnsIns_MixOneColumnInst_1_n24), .ZN(MixColumnsOutput[88]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U59 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n23), .B(MixColumnsInput[64]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n25) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U58 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n22), .B(
        MixColumnsIns_MixOneColumnInst_1_n42), .ZN(MixColumnsOutput[87]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U57 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n42) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U56 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B(
        MixColumnsIns_MixOneColumnInst_1_n21), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n22) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U55 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n20), .B(
        MixColumnsIns_MixOneColumnInst_1_n40), .ZN(MixColumnsOutput[86]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U54 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n40) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U53 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .B(
        MixColumnsIns_MixOneColumnInst_1_n19), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n20) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U52 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n18), .B(
        MixColumnsIns_MixOneColumnInst_1_n35), .ZN(MixColumnsOutput[85]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U51 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n35) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U50 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .B(
        MixColumnsIns_MixOneColumnInst_1_n17), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n18) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U49 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n16), .B(
        MixColumnsIns_MixOneColumnInst_1_n33), .ZN(MixColumnsOutput[84]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U48 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n33) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U47 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .B(
        MixColumnsIns_MixOneColumnInst_1_n15), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n16) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U46 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n14), .B(
        MixColumnsIns_MixOneColumnInst_1_n27), .ZN(MixColumnsOutput[65]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U45 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n27) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U44 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .B(
        MixColumnsIns_MixOneColumnInst_1_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n14) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U43 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n62) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U42 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n13), .B(
        MixColumnsIns_MixOneColumnInst_1_n31), .ZN(MixColumnsOutput[83]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U41 ( .A(MixColumnsInput[75]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n31) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U40 ( .A(MixColumnsInput[91]), .B(
        MixColumnsIns_MixOneColumnInst_1_n12), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n13) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U39 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n11), .B(
        MixColumnsIns_MixOneColumnInst_1_n29), .ZN(MixColumnsOutput[82]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U38 ( .A(MixColumnsInput[74]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n29) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U37 ( .A(MixColumnsInput[90]), .B(
        MixColumnsIns_MixOneColumnInst_1_n10), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n11) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U36 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n9), .B(
        MixColumnsIns_MixOneColumnInst_1_n26), .ZN(MixColumnsOutput[81]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U35 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n26) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U34 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n63), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n9) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U33 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n63) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U32 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n8), .B(
        MixColumnsIns_MixOneColumnInst_1_n24), .ZN(MixColumnsOutput[80]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U31 ( .A(MixColumnsInput[72]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n24) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U30 ( .A(MixColumnsInput[88]), .B(
        MixColumnsIns_MixOneColumnInst_1_n60), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n8) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U29 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsInput[64]), .Z(MixColumnsIns_MixOneColumnInst_1_n60) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U28 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n7), .B(
        MixColumnsIns_MixOneColumnInst_1_n21), .ZN(MixColumnsOutput[79]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U27 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n21) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U26 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n56), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n7) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U25 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n56) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U24 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n6), .B(
        MixColumnsIns_MixOneColumnInst_1_n19), .ZN(MixColumnsOutput[78]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U23 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n19) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U22 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n53), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n6) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U21 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n53) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U20 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n5), .B(
        MixColumnsIns_MixOneColumnInst_1_n17), .ZN(MixColumnsOutput[77]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U19 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n17) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U18 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n50), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n5) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U17 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n50) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U16 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n4), .B(
        MixColumnsIns_MixOneColumnInst_1_n15), .ZN(MixColumnsOutput[76]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U15 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n15) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U14 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n47), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n4) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U13 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n47) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U12 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n3), .B(
        MixColumnsIns_MixOneColumnInst_1_n12), .ZN(MixColumnsOutput[75]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U11 ( .A(MixColumnsInput[67]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n12) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U10 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n44), .B(MixColumnsInput[83]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n3) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U9 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]), .B(
        MixColumnsInput[91]), .Z(MixColumnsIns_MixOneColumnInst_1_n44) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U8 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n2), .B(
        MixColumnsIns_MixOneColumnInst_1_n10), .ZN(MixColumnsOutput[74]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U7 ( .A(MixColumnsInput[66]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n10) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U6 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n37), .B(MixColumnsInput[82]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n2) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U5 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .B(
        MixColumnsInput[90]), .Z(MixColumnsIns_MixOneColumnInst_1_n37) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U4 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n1), .B(MixColumnsInput[72]), .ZN(
        MixColumnsOutput[64]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n59), .B(
        MixColumnsIns_MixOneColumnInst_1_n23), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n1) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U2 ( .A(MixColumnsInput[80]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n23) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsInput[88]), .Z(MixColumnsIns_MixOneColumnInst_1_n59) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B(
        MixColumnsInput[91]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B(
        MixColumnsInput[90]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B(
        MixColumnsInput[88]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B(
        MixColumnsInput[83]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B(
        MixColumnsInput[82]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B(
        MixColumnsInput[80]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsInput[75]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsInput[74]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsInput[72]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsInput[67]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsInput[66]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsInput[64]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U96 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n64), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .ZN(
        MixColumnsOutput[41]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U95 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n63), .B(
        MixColumnsIns_MixOneColumnInst_2_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n64) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U94 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n61), .B(
        MixColumnsIns_MixOneColumnInst_2_n60), .ZN(MixColumnsOutput[40]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U93 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n59), .B(MixColumnsInput[48]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n61) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U92 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n58), .B(
        MixColumnsIns_MixOneColumnInst_2_n57), .ZN(MixColumnsOutput[39]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U91 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n56), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n58) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U90 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n55), .B(
        MixColumnsIns_MixOneColumnInst_2_n54), .ZN(MixColumnsOutput[38]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U89 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n53), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n55) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U88 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n52), .B(
        MixColumnsIns_MixOneColumnInst_2_n51), .ZN(MixColumnsOutput[37]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U87 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n50), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n52) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U86 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n49), .B(
        MixColumnsIns_MixOneColumnInst_2_n48), .ZN(MixColumnsOutput[36]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U85 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n47), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n49) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U84 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n46), .B(
        MixColumnsIns_MixOneColumnInst_2_n45), .ZN(MixColumnsOutput[35]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U83 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n44), .B(MixColumnsInput[43]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n46) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U82 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n43), .B(
        MixColumnsIns_MixOneColumnInst_2_n57), .ZN(MixColumnsOutput[63]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U81 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n57) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U80 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_2_n42), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n43) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U79 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n41), .B(
        MixColumnsIns_MixOneColumnInst_2_n54), .ZN(MixColumnsOutput[62]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U78 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n54) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U77 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_2_n40), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n41) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U76 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n39), .B(
        MixColumnsIns_MixOneColumnInst_2_n38), .ZN(MixColumnsOutput[34]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U75 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n37), .B(MixColumnsInput[42]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n39) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U74 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n36), .B(
        MixColumnsIns_MixOneColumnInst_2_n51), .ZN(MixColumnsOutput[61]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U73 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n51) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U72 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_2_n35), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n36) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U71 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n34), .B(
        MixColumnsIns_MixOneColumnInst_2_n48), .ZN(MixColumnsOutput[60]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U70 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n48) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U69 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_2_n33), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n34) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U68 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n32), .B(
        MixColumnsIns_MixOneColumnInst_2_n45), .ZN(MixColumnsOutput[59]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U67 ( .A(MixColumnsInput[51]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n45) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U66 ( .A(MixColumnsInput[35]), .B(
        MixColumnsIns_MixOneColumnInst_2_n31), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n32) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U65 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n30), .B(
        MixColumnsIns_MixOneColumnInst_2_n38), .ZN(MixColumnsOutput[58]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U64 ( .A(MixColumnsInput[50]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n38) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U63 ( .A(MixColumnsInput[34]), .B(
        MixColumnsIns_MixOneColumnInst_2_n29), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n30) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U62 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n28), .B(
        MixColumnsIns_MixOneColumnInst_2_n27), .ZN(MixColumnsOutput[57]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U61 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .B(
        MixColumnsIns_MixOneColumnInst_2_n26), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n28) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U60 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n25), .B(
        MixColumnsIns_MixOneColumnInst_2_n24), .ZN(MixColumnsOutput[56]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U59 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n23), .B(MixColumnsInput[32]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n25) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U58 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n22), .B(
        MixColumnsIns_MixOneColumnInst_2_n42), .ZN(MixColumnsOutput[55]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U57 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n42) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U56 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B(
        MixColumnsIns_MixOneColumnInst_2_n21), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n22) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U55 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n20), .B(
        MixColumnsIns_MixOneColumnInst_2_n40), .ZN(MixColumnsOutput[54]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U54 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n40) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U53 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .B(
        MixColumnsIns_MixOneColumnInst_2_n19), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n20) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U52 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n18), .B(
        MixColumnsIns_MixOneColumnInst_2_n35), .ZN(MixColumnsOutput[53]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U51 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n35) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U50 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .B(
        MixColumnsIns_MixOneColumnInst_2_n17), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n18) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U49 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n16), .B(
        MixColumnsIns_MixOneColumnInst_2_n33), .ZN(MixColumnsOutput[52]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U48 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n33) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U47 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .B(
        MixColumnsIns_MixOneColumnInst_2_n15), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n16) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U46 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n14), .B(
        MixColumnsIns_MixOneColumnInst_2_n27), .ZN(MixColumnsOutput[33]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U45 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n27) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U44 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .B(
        MixColumnsIns_MixOneColumnInst_2_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n14) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U43 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n62) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U42 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n13), .B(
        MixColumnsIns_MixOneColumnInst_2_n31), .ZN(MixColumnsOutput[51]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U41 ( .A(MixColumnsInput[43]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n31) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U40 ( .A(MixColumnsInput[59]), .B(
        MixColumnsIns_MixOneColumnInst_2_n12), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n13) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U39 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n11), .B(
        MixColumnsIns_MixOneColumnInst_2_n29), .ZN(MixColumnsOutput[50]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U38 ( .A(MixColumnsInput[42]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n29) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U37 ( .A(MixColumnsInput[58]), .B(
        MixColumnsIns_MixOneColumnInst_2_n10), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n11) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U36 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n9), .B(
        MixColumnsIns_MixOneColumnInst_2_n26), .ZN(MixColumnsOutput[49]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U35 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n26) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U34 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n63), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n9) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U33 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n63) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U32 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n8), .B(
        MixColumnsIns_MixOneColumnInst_2_n24), .ZN(MixColumnsOutput[48]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U31 ( .A(MixColumnsInput[40]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n24) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U30 ( .A(MixColumnsInput[56]), .B(
        MixColumnsIns_MixOneColumnInst_2_n60), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n8) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U29 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsInput[32]), .Z(MixColumnsIns_MixOneColumnInst_2_n60) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U28 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n7), .B(
        MixColumnsIns_MixOneColumnInst_2_n21), .ZN(MixColumnsOutput[47]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U27 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n21) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U26 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n56), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n7) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U25 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n56) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U24 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n6), .B(
        MixColumnsIns_MixOneColumnInst_2_n19), .ZN(MixColumnsOutput[46]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U23 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n19) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U22 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n53), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n6) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U21 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n53) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U20 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n5), .B(
        MixColumnsIns_MixOneColumnInst_2_n17), .ZN(MixColumnsOutput[45]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U19 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n17) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U18 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n50), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n5) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U17 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n50) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U16 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n4), .B(
        MixColumnsIns_MixOneColumnInst_2_n15), .ZN(MixColumnsOutput[44]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U15 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n15) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U14 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n47), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n4) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U13 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n47) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U12 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n3), .B(
        MixColumnsIns_MixOneColumnInst_2_n12), .ZN(MixColumnsOutput[43]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U11 ( .A(MixColumnsInput[35]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n12) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U10 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n44), .B(MixColumnsInput[51]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n3) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U9 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]), .B(
        MixColumnsInput[59]), .Z(MixColumnsIns_MixOneColumnInst_2_n44) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U8 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n2), .B(
        MixColumnsIns_MixOneColumnInst_2_n10), .ZN(MixColumnsOutput[42]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U7 ( .A(MixColumnsInput[34]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n10) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U6 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n37), .B(MixColumnsInput[50]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n2) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U5 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .B(
        MixColumnsInput[58]), .Z(MixColumnsIns_MixOneColumnInst_2_n37) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U4 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n1), .B(MixColumnsInput[40]), .ZN(
        MixColumnsOutput[32]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n59), .B(
        MixColumnsIns_MixOneColumnInst_2_n23), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n1) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U2 ( .A(MixColumnsInput[48]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n23) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsInput[56]), .Z(MixColumnsIns_MixOneColumnInst_2_n59) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B(
        MixColumnsInput[59]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B(
        MixColumnsInput[58]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B(
        MixColumnsInput[56]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B(
        MixColumnsInput[51]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B(
        MixColumnsInput[50]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B(
        MixColumnsInput[48]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsInput[43]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsInput[42]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsInput[40]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsInput[35]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsInput[34]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsInput[32]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U96 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n64), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .ZN(
        MixColumnsOutput[9]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U95 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n63), .B(
        MixColumnsIns_MixOneColumnInst_3_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n64) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U94 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n61), .B(
        MixColumnsIns_MixOneColumnInst_3_n60), .ZN(MixColumnsOutput[8]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U93 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n59), .B(MixColumnsInput[16]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n61) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U92 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n58), .B(
        MixColumnsIns_MixOneColumnInst_3_n57), .ZN(MixColumnsOutput[7]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U91 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n56), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n58) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U90 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n55), .B(
        MixColumnsIns_MixOneColumnInst_3_n54), .ZN(MixColumnsOutput[6]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U89 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n53), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n55) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U88 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n52), .B(
        MixColumnsIns_MixOneColumnInst_3_n51), .ZN(MixColumnsOutput[5]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U87 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n50), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n52) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U86 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n49), .B(
        MixColumnsIns_MixOneColumnInst_3_n48), .ZN(MixColumnsOutput[4]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U85 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n47), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n49) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U84 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n46), .B(
        MixColumnsIns_MixOneColumnInst_3_n45), .ZN(MixColumnsOutput[3]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U83 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n44), .B(MixColumnsInput[11]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n46) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U82 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n43), .B(
        MixColumnsIns_MixOneColumnInst_3_n57), .ZN(MixColumnsOutput[31]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U81 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n57) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U80 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_3_n42), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n43) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U79 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n41), .B(
        MixColumnsIns_MixOneColumnInst_3_n54), .ZN(MixColumnsOutput[30]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U78 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n54) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U77 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_3_n40), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n41) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U76 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n39), .B(
        MixColumnsIns_MixOneColumnInst_3_n38), .ZN(MixColumnsOutput[2]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U75 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n37), .B(MixColumnsInput[10]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n39) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U74 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n36), .B(
        MixColumnsIns_MixOneColumnInst_3_n51), .ZN(MixColumnsOutput[29]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U73 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n51) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U72 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_3_n35), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n36) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U71 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n34), .B(
        MixColumnsIns_MixOneColumnInst_3_n48), .ZN(MixColumnsOutput[28]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U70 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n48) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U69 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_3_n33), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n34) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U68 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n32), .B(
        MixColumnsIns_MixOneColumnInst_3_n45), .ZN(MixColumnsOutput[27]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U67 ( .A(MixColumnsInput[19]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n45) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U66 ( .A(MixColumnsInput[3]), .B(
        MixColumnsIns_MixOneColumnInst_3_n31), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n32) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U65 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n30), .B(
        MixColumnsIns_MixOneColumnInst_3_n38), .ZN(MixColumnsOutput[26]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U64 ( .A(MixColumnsInput[18]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n38) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U63 ( .A(MixColumnsInput[2]), .B(
        MixColumnsIns_MixOneColumnInst_3_n29), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n30) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U62 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n28), .B(
        MixColumnsIns_MixOneColumnInst_3_n27), .ZN(MixColumnsOutput[25]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U61 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .B(
        MixColumnsIns_MixOneColumnInst_3_n26), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n28) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U60 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n25), .B(
        MixColumnsIns_MixOneColumnInst_3_n24), .ZN(MixColumnsOutput[24]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U59 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n23), .B(MixColumnsInput[0]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n25) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U58 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n22), .B(
        MixColumnsIns_MixOneColumnInst_3_n42), .ZN(MixColumnsOutput[23]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U57 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n42) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U56 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B(
        MixColumnsIns_MixOneColumnInst_3_n21), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n22) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U55 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n20), .B(
        MixColumnsIns_MixOneColumnInst_3_n40), .ZN(MixColumnsOutput[22]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U54 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n40) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U53 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .B(
        MixColumnsIns_MixOneColumnInst_3_n19), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n20) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U52 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n18), .B(
        MixColumnsIns_MixOneColumnInst_3_n35), .ZN(MixColumnsOutput[21]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U51 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n35) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U50 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .B(
        MixColumnsIns_MixOneColumnInst_3_n17), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n18) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U49 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n16), .B(
        MixColumnsIns_MixOneColumnInst_3_n33), .ZN(MixColumnsOutput[20]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U48 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n33) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U47 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .B(
        MixColumnsIns_MixOneColumnInst_3_n15), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n16) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U46 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n14), .B(
        MixColumnsIns_MixOneColumnInst_3_n27), .ZN(MixColumnsOutput[1]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U45 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n27) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U44 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .B(
        MixColumnsIns_MixOneColumnInst_3_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n14) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U43 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n62) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U42 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n13), .B(
        MixColumnsIns_MixOneColumnInst_3_n31), .ZN(MixColumnsOutput[19]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U41 ( .A(MixColumnsInput[11]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n31) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U40 ( .A(MixColumnsInput[27]), .B(
        MixColumnsIns_MixOneColumnInst_3_n12), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n13) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U39 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n11), .B(
        MixColumnsIns_MixOneColumnInst_3_n29), .ZN(MixColumnsOutput[18]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U38 ( .A(MixColumnsInput[10]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n29) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U37 ( .A(MixColumnsInput[26]), .B(
        MixColumnsIns_MixOneColumnInst_3_n10), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n11) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U36 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n9), .B(
        MixColumnsIns_MixOneColumnInst_3_n26), .ZN(MixColumnsOutput[17]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U35 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n26) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U34 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n63), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n9) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U33 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n63) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U32 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n8), .B(
        MixColumnsIns_MixOneColumnInst_3_n24), .ZN(MixColumnsOutput[16]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U31 ( .A(MixColumnsInput[8]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n24) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U30 ( .A(MixColumnsInput[24]), .B(
        MixColumnsIns_MixOneColumnInst_3_n60), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n8) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U29 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsInput[0]), .Z(MixColumnsIns_MixOneColumnInst_3_n60) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U28 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n7), .B(
        MixColumnsIns_MixOneColumnInst_3_n21), .ZN(MixColumnsOutput[15]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U27 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n21) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U26 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n56), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n7) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U25 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n56) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U24 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n6), .B(
        MixColumnsIns_MixOneColumnInst_3_n19), .ZN(MixColumnsOutput[14]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U23 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n19) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U22 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n53), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n6) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U21 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n53) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U20 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n5), .B(
        MixColumnsIns_MixOneColumnInst_3_n17), .ZN(MixColumnsOutput[13]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U19 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n17) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U18 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n50), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n5) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U17 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n50) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U16 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n4), .B(
        MixColumnsIns_MixOneColumnInst_3_n15), .ZN(MixColumnsOutput[12]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U15 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n15) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U14 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n47), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n4) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U13 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n47) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U12 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n3), .B(
        MixColumnsIns_MixOneColumnInst_3_n12), .ZN(MixColumnsOutput[11]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U11 ( .A(MixColumnsInput[3]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n12) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U10 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n44), .B(MixColumnsInput[19]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n3) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U9 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]), .B(
        MixColumnsInput[27]), .Z(MixColumnsIns_MixOneColumnInst_3_n44) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U8 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n2), .B(
        MixColumnsIns_MixOneColumnInst_3_n10), .ZN(MixColumnsOutput[10]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U7 ( .A(MixColumnsInput[2]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n10) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U6 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n37), .B(MixColumnsInput[18]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n2) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U5 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .B(
        MixColumnsInput[26]), .Z(MixColumnsIns_MixOneColumnInst_3_n37) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U4 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n1), .B(MixColumnsInput[8]), .ZN(
        MixColumnsOutput[0]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n59), .B(
        MixColumnsIns_MixOneColumnInst_3_n23), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n1) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U2 ( .A(MixColumnsInput[16]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n23) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsInput[24]), .Z(MixColumnsIns_MixOneColumnInst_3_n59) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B(
        MixColumnsInput[27]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B(
        MixColumnsInput[26]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B(
        MixColumnsInput[24]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B(
        MixColumnsInput[19]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B(
        MixColumnsInput[18]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B(
        MixColumnsInput[16]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsInput[11]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsInput[10]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsInput[8]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsInput[3]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsInput[2]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsInput[0]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]) );
  MUX2_X1 KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .A(KeyExpansionOutput[0]), .B(
        key[0]), .S(reset), .Z(KeyReg_Inst_ff_SDE_0_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_0_current_state_reg_U1 ( .A(RoundKey[0]), .ZN(
        KeyReg_Inst_ff_SDE_0_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_0_next_state), .CK(clk), .Q(RoundKey[0]), .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .A(KeyExpansionOutput[1]), .B(
        key[1]), .S(reset), .Z(KeyReg_Inst_ff_SDE_1_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_1_current_state_reg_U1 ( .A(RoundKey[1]), .ZN(
        KeyReg_Inst_ff_SDE_1_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_1_next_state), .CK(clk), .Q(RoundKey[1]), .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .A(KeyExpansionOutput[2]), .B(
        key[2]), .S(reset), .Z(KeyReg_Inst_ff_SDE_2_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_2_current_state_reg_U1 ( .A(RoundKey[2]), .ZN(
        KeyReg_Inst_ff_SDE_2_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_2_next_state), .CK(clk), .Q(RoundKey[2]), .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .A(KeyExpansionOutput[3]), .B(
        key[3]), .S(reset), .Z(KeyReg_Inst_ff_SDE_3_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_3_current_state_reg_U1 ( .A(RoundKey[3]), .ZN(
        KeyReg_Inst_ff_SDE_3_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_3_next_state), .CK(clk), .Q(RoundKey[3]), .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .A(KeyExpansionOutput[4]), .B(
        key[4]), .S(reset), .Z(KeyReg_Inst_ff_SDE_4_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_4_current_state_reg_U1 ( .A(RoundKey[4]), .ZN(
        KeyReg_Inst_ff_SDE_4_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_4_next_state), .CK(clk), .Q(RoundKey[4]), .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .A(KeyExpansionOutput[5]), .B(
        key[5]), .S(reset), .Z(KeyReg_Inst_ff_SDE_5_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_5_current_state_reg_U1 ( .A(RoundKey[5]), .ZN(
        KeyReg_Inst_ff_SDE_5_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_5_next_state), .CK(clk), .Q(RoundKey[5]), .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .A(KeyExpansionOutput[6]), .B(
        key[6]), .S(reset), .Z(KeyReg_Inst_ff_SDE_6_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_6_current_state_reg_U1 ( .A(RoundKey[6]), .ZN(
        KeyReg_Inst_ff_SDE_6_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_6_next_state), .CK(clk), .Q(RoundKey[6]), .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .A(KeyExpansionOutput[7]), .B(
        key[7]), .S(reset), .Z(KeyReg_Inst_ff_SDE_7_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_7_current_state_reg_U1 ( .A(RoundKey[7]), .ZN(
        KeyReg_Inst_ff_SDE_7_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_7_next_state), .CK(clk), .Q(RoundKey[7]), .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .A(KeyExpansionOutput[8]), .B(
        key[8]), .S(reset), .Z(KeyReg_Inst_ff_SDE_8_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_8_current_state_reg_U1 ( .A(RoundKey[8]), .ZN(
        KeyReg_Inst_ff_SDE_8_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_8_next_state), .CK(clk), .Q(RoundKey[8]), .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .A(KeyExpansionOutput[9]), .B(
        key[9]), .S(reset), .Z(KeyReg_Inst_ff_SDE_9_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_9_current_state_reg_U1 ( .A(RoundKey[9]), .ZN(
        KeyReg_Inst_ff_SDE_9_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_9_next_state), .CK(clk), .Q(RoundKey[9]), .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .A(KeyExpansionOutput[10]), .B(
        key[10]), .S(reset), .Z(KeyReg_Inst_ff_SDE_10_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_10_current_state_reg_U1 ( .A(RoundKey[10]), .ZN(
        KeyReg_Inst_ff_SDE_10_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_10_next_state), .CK(clk), .Q(RoundKey[10]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .A(KeyExpansionOutput[11]), .B(
        key[11]), .S(reset), .Z(KeyReg_Inst_ff_SDE_11_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_11_current_state_reg_U1 ( .A(RoundKey[11]), .ZN(
        KeyReg_Inst_ff_SDE_11_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_11_next_state), .CK(clk), .Q(RoundKey[11]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .A(KeyExpansionOutput[12]), .B(
        key[12]), .S(reset), .Z(KeyReg_Inst_ff_SDE_12_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_12_current_state_reg_U1 ( .A(RoundKey[12]), .ZN(
        KeyReg_Inst_ff_SDE_12_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_12_next_state), .CK(clk), .Q(RoundKey[12]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .A(KeyExpansionOutput[13]), .B(
        key[13]), .S(reset), .Z(KeyReg_Inst_ff_SDE_13_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_13_current_state_reg_U1 ( .A(RoundKey[13]), .ZN(
        KeyReg_Inst_ff_SDE_13_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_13_next_state), .CK(clk), .Q(RoundKey[13]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .A(KeyExpansionOutput[14]), .B(
        key[14]), .S(reset), .Z(KeyReg_Inst_ff_SDE_14_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_14_current_state_reg_U1 ( .A(RoundKey[14]), .ZN(
        KeyReg_Inst_ff_SDE_14_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_14_next_state), .CK(clk), .Q(RoundKey[14]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .A(KeyExpansionOutput[15]), .B(
        key[15]), .S(reset), .Z(KeyReg_Inst_ff_SDE_15_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_15_current_state_reg_U1 ( .A(RoundKey[15]), .ZN(
        KeyReg_Inst_ff_SDE_15_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_15_next_state), .CK(clk), .Q(RoundKey[15]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .A(KeyExpansionOutput[16]), .B(
        key[16]), .S(reset), .Z(KeyReg_Inst_ff_SDE_16_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_16_current_state_reg_U1 ( .A(RoundKey[16]), .ZN(
        KeyReg_Inst_ff_SDE_16_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_16_next_state), .CK(clk), .Q(RoundKey[16]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .A(KeyExpansionOutput[17]), .B(
        key[17]), .S(reset), .Z(KeyReg_Inst_ff_SDE_17_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_17_current_state_reg_U1 ( .A(RoundKey[17]), .ZN(
        KeyReg_Inst_ff_SDE_17_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_17_next_state), .CK(clk), .Q(RoundKey[17]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .A(KeyExpansionOutput[18]), .B(
        key[18]), .S(reset), .Z(KeyReg_Inst_ff_SDE_18_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_18_current_state_reg_U1 ( .A(RoundKey[18]), .ZN(
        KeyReg_Inst_ff_SDE_18_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_18_next_state), .CK(clk), .Q(RoundKey[18]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .A(KeyExpansionOutput[19]), .B(
        key[19]), .S(reset), .Z(KeyReg_Inst_ff_SDE_19_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_19_current_state_reg_U1 ( .A(RoundKey[19]), .ZN(
        KeyReg_Inst_ff_SDE_19_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_19_next_state), .CK(clk), .Q(RoundKey[19]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .A(KeyExpansionOutput[20]), .B(
        key[20]), .S(reset), .Z(KeyReg_Inst_ff_SDE_20_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_20_current_state_reg_U1 ( .A(RoundKey[20]), .ZN(
        KeyReg_Inst_ff_SDE_20_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_20_next_state), .CK(clk), .Q(RoundKey[20]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .A(KeyExpansionOutput[21]), .B(
        key[21]), .S(reset), .Z(KeyReg_Inst_ff_SDE_21_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_21_current_state_reg_U1 ( .A(RoundKey[21]), .ZN(
        KeyReg_Inst_ff_SDE_21_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_21_next_state), .CK(clk), .Q(RoundKey[21]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .A(KeyExpansionOutput[22]), .B(
        key[22]), .S(reset), .Z(KeyReg_Inst_ff_SDE_22_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_22_current_state_reg_U1 ( .A(RoundKey[22]), .ZN(
        KeyReg_Inst_ff_SDE_22_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_22_next_state), .CK(clk), .Q(RoundKey[22]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .A(KeyExpansionOutput[23]), .B(
        key[23]), .S(reset), .Z(KeyReg_Inst_ff_SDE_23_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_23_current_state_reg_U1 ( .A(RoundKey[23]), .ZN(
        KeyReg_Inst_ff_SDE_23_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_23_next_state), .CK(clk), .Q(RoundKey[23]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .A(KeyExpansionOutput[24]), .B(
        key[24]), .S(reset), .Z(KeyReg_Inst_ff_SDE_24_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_24_current_state_reg_U1 ( .A(RoundKey[24]), .ZN(
        KeyReg_Inst_ff_SDE_24_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_24_next_state), .CK(clk), .Q(RoundKey[24]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .A(KeyExpansionOutput[25]), .B(
        key[25]), .S(reset), .Z(KeyReg_Inst_ff_SDE_25_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_25_current_state_reg_U1 ( .A(RoundKey[25]), .ZN(
        KeyReg_Inst_ff_SDE_25_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_25_next_state), .CK(clk), .Q(RoundKey[25]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .A(KeyExpansionOutput[26]), .B(
        key[26]), .S(reset), .Z(KeyReg_Inst_ff_SDE_26_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_26_current_state_reg_U1 ( .A(RoundKey[26]), .ZN(
        KeyReg_Inst_ff_SDE_26_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_26_next_state), .CK(clk), .Q(RoundKey[26]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .A(KeyExpansionOutput[27]), .B(
        key[27]), .S(reset), .Z(KeyReg_Inst_ff_SDE_27_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_27_current_state_reg_U1 ( .A(RoundKey[27]), .ZN(
        KeyReg_Inst_ff_SDE_27_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_27_next_state), .CK(clk), .Q(RoundKey[27]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .A(KeyExpansionOutput[28]), .B(
        key[28]), .S(reset), .Z(KeyReg_Inst_ff_SDE_28_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_28_current_state_reg_U1 ( .A(RoundKey[28]), .ZN(
        KeyReg_Inst_ff_SDE_28_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_28_next_state), .CK(clk), .Q(RoundKey[28]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .A(KeyExpansionOutput[29]), .B(
        key[29]), .S(reset), .Z(KeyReg_Inst_ff_SDE_29_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_29_current_state_reg_U1 ( .A(RoundKey[29]), .ZN(
        KeyReg_Inst_ff_SDE_29_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_29_next_state), .CK(clk), .Q(RoundKey[29]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .A(KeyExpansionOutput[30]), .B(
        key[30]), .S(reset), .Z(KeyReg_Inst_ff_SDE_30_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_30_current_state_reg_U1 ( .A(RoundKey[30]), .ZN(
        KeyReg_Inst_ff_SDE_30_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_30_next_state), .CK(clk), .Q(RoundKey[30]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .A(KeyExpansionOutput[31]), .B(
        key[31]), .S(reset), .Z(KeyReg_Inst_ff_SDE_31_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_31_current_state_reg_U1 ( .A(RoundKey[31]), .ZN(
        KeyReg_Inst_ff_SDE_31_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_31_next_state), .CK(clk), .Q(RoundKey[31]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .A(KeyExpansionOutput[32]), .B(
        key[32]), .S(reset), .Z(KeyReg_Inst_ff_SDE_32_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_32_current_state_reg_U1 ( .A(RoundKey[32]), .ZN(
        KeyReg_Inst_ff_SDE_32_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_32_next_state), .CK(clk), .Q(RoundKey[32]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .A(KeyExpansionOutput[33]), .B(
        key[33]), .S(reset), .Z(KeyReg_Inst_ff_SDE_33_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_33_current_state_reg_U1 ( .A(RoundKey[33]), .ZN(
        KeyReg_Inst_ff_SDE_33_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_33_next_state), .CK(clk), .Q(RoundKey[33]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .A(KeyExpansionOutput[34]), .B(
        key[34]), .S(reset), .Z(KeyReg_Inst_ff_SDE_34_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_34_current_state_reg_U1 ( .A(RoundKey[34]), .ZN(
        KeyReg_Inst_ff_SDE_34_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_34_next_state), .CK(clk), .Q(RoundKey[34]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .A(KeyExpansionOutput[35]), .B(
        key[35]), .S(reset), .Z(KeyReg_Inst_ff_SDE_35_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_35_current_state_reg_U1 ( .A(RoundKey[35]), .ZN(
        KeyReg_Inst_ff_SDE_35_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_35_next_state), .CK(clk), .Q(RoundKey[35]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .A(KeyExpansionOutput[36]), .B(
        key[36]), .S(reset), .Z(KeyReg_Inst_ff_SDE_36_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_36_current_state_reg_U1 ( .A(RoundKey[36]), .ZN(
        KeyReg_Inst_ff_SDE_36_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_36_next_state), .CK(clk), .Q(RoundKey[36]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .A(KeyExpansionOutput[37]), .B(
        key[37]), .S(reset), .Z(KeyReg_Inst_ff_SDE_37_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_37_current_state_reg_U1 ( .A(RoundKey[37]), .ZN(
        KeyReg_Inst_ff_SDE_37_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_37_next_state), .CK(clk), .Q(RoundKey[37]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .A(KeyExpansionOutput[38]), .B(
        key[38]), .S(reset), .Z(KeyReg_Inst_ff_SDE_38_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_38_current_state_reg_U1 ( .A(RoundKey[38]), .ZN(
        KeyReg_Inst_ff_SDE_38_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_38_next_state), .CK(clk), .Q(RoundKey[38]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .A(KeyExpansionOutput[39]), .B(
        key[39]), .S(reset), .Z(KeyReg_Inst_ff_SDE_39_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_39_current_state_reg_U1 ( .A(RoundKey[39]), .ZN(
        KeyReg_Inst_ff_SDE_39_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_39_next_state), .CK(clk), .Q(RoundKey[39]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .A(KeyExpansionOutput[40]), .B(
        key[40]), .S(reset), .Z(KeyReg_Inst_ff_SDE_40_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_40_current_state_reg_U1 ( .A(RoundKey[40]), .ZN(
        KeyReg_Inst_ff_SDE_40_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_40_next_state), .CK(clk), .Q(RoundKey[40]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .A(KeyExpansionOutput[41]), .B(
        key[41]), .S(reset), .Z(KeyReg_Inst_ff_SDE_41_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_41_current_state_reg_U1 ( .A(RoundKey[41]), .ZN(
        KeyReg_Inst_ff_SDE_41_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_41_next_state), .CK(clk), .Q(RoundKey[41]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .A(KeyExpansionOutput[42]), .B(
        key[42]), .S(reset), .Z(KeyReg_Inst_ff_SDE_42_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_42_current_state_reg_U1 ( .A(RoundKey[42]), .ZN(
        KeyReg_Inst_ff_SDE_42_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_42_next_state), .CK(clk), .Q(RoundKey[42]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .A(KeyExpansionOutput[43]), .B(
        key[43]), .S(reset), .Z(KeyReg_Inst_ff_SDE_43_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_43_current_state_reg_U1 ( .A(RoundKey[43]), .ZN(
        KeyReg_Inst_ff_SDE_43_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_43_next_state), .CK(clk), .Q(RoundKey[43]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .A(KeyExpansionOutput[44]), .B(
        key[44]), .S(reset), .Z(KeyReg_Inst_ff_SDE_44_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_44_current_state_reg_U1 ( .A(RoundKey[44]), .ZN(
        KeyReg_Inst_ff_SDE_44_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_44_next_state), .CK(clk), .Q(RoundKey[44]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .A(KeyExpansionOutput[45]), .B(
        key[45]), .S(reset), .Z(KeyReg_Inst_ff_SDE_45_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_45_current_state_reg_U1 ( .A(RoundKey[45]), .ZN(
        KeyReg_Inst_ff_SDE_45_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_45_next_state), .CK(clk), .Q(RoundKey[45]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .A(KeyExpansionOutput[46]), .B(
        key[46]), .S(reset), .Z(KeyReg_Inst_ff_SDE_46_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_46_current_state_reg_U1 ( .A(RoundKey[46]), .ZN(
        KeyReg_Inst_ff_SDE_46_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_46_next_state), .CK(clk), .Q(RoundKey[46]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .A(KeyExpansionOutput[47]), .B(
        key[47]), .S(reset), .Z(KeyReg_Inst_ff_SDE_47_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_47_current_state_reg_U1 ( .A(RoundKey[47]), .ZN(
        KeyReg_Inst_ff_SDE_47_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_47_next_state), .CK(clk), .Q(RoundKey[47]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .A(KeyExpansionOutput[48]), .B(
        key[48]), .S(reset), .Z(KeyReg_Inst_ff_SDE_48_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_48_current_state_reg_U1 ( .A(RoundKey[48]), .ZN(
        KeyReg_Inst_ff_SDE_48_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_48_next_state), .CK(clk), .Q(RoundKey[48]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .A(KeyExpansionOutput[49]), .B(
        key[49]), .S(reset), .Z(KeyReg_Inst_ff_SDE_49_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_49_current_state_reg_U1 ( .A(RoundKey[49]), .ZN(
        KeyReg_Inst_ff_SDE_49_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_49_next_state), .CK(clk), .Q(RoundKey[49]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .A(KeyExpansionOutput[50]), .B(
        key[50]), .S(reset), .Z(KeyReg_Inst_ff_SDE_50_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_50_current_state_reg_U1 ( .A(RoundKey[50]), .ZN(
        KeyReg_Inst_ff_SDE_50_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_50_next_state), .CK(clk), .Q(RoundKey[50]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .A(KeyExpansionOutput[51]), .B(
        key[51]), .S(reset), .Z(KeyReg_Inst_ff_SDE_51_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_51_current_state_reg_U1 ( .A(RoundKey[51]), .ZN(
        KeyReg_Inst_ff_SDE_51_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_51_next_state), .CK(clk), .Q(RoundKey[51]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .A(KeyExpansionOutput[52]), .B(
        key[52]), .S(reset), .Z(KeyReg_Inst_ff_SDE_52_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_52_current_state_reg_U1 ( .A(RoundKey[52]), .ZN(
        KeyReg_Inst_ff_SDE_52_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_52_next_state), .CK(clk), .Q(RoundKey[52]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .A(KeyExpansionOutput[53]), .B(
        key[53]), .S(reset), .Z(KeyReg_Inst_ff_SDE_53_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_53_current_state_reg_U1 ( .A(RoundKey[53]), .ZN(
        KeyReg_Inst_ff_SDE_53_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_53_next_state), .CK(clk), .Q(RoundKey[53]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .A(KeyExpansionOutput[54]), .B(
        key[54]), .S(reset), .Z(KeyReg_Inst_ff_SDE_54_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_54_current_state_reg_U1 ( .A(RoundKey[54]), .ZN(
        KeyReg_Inst_ff_SDE_54_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_54_next_state), .CK(clk), .Q(RoundKey[54]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .A(KeyExpansionOutput[55]), .B(
        key[55]), .S(reset), .Z(KeyReg_Inst_ff_SDE_55_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_55_current_state_reg_U1 ( .A(RoundKey[55]), .ZN(
        KeyReg_Inst_ff_SDE_55_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_55_next_state), .CK(clk), .Q(RoundKey[55]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .A(KeyExpansionOutput[56]), .B(
        key[56]), .S(reset), .Z(KeyReg_Inst_ff_SDE_56_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_56_current_state_reg_U1 ( .A(RoundKey[56]), .ZN(
        KeyReg_Inst_ff_SDE_56_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_56_next_state), .CK(clk), .Q(RoundKey[56]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .A(KeyExpansionOutput[57]), .B(
        key[57]), .S(reset), .Z(KeyReg_Inst_ff_SDE_57_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_57_current_state_reg_U1 ( .A(RoundKey[57]), .ZN(
        KeyReg_Inst_ff_SDE_57_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_57_next_state), .CK(clk), .Q(RoundKey[57]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .A(KeyExpansionOutput[58]), .B(
        key[58]), .S(reset), .Z(KeyReg_Inst_ff_SDE_58_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_58_current_state_reg_U1 ( .A(RoundKey[58]), .ZN(
        KeyReg_Inst_ff_SDE_58_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_58_next_state), .CK(clk), .Q(RoundKey[58]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .A(KeyExpansionOutput[59]), .B(
        key[59]), .S(reset), .Z(KeyReg_Inst_ff_SDE_59_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_59_current_state_reg_U1 ( .A(RoundKey[59]), .ZN(
        KeyReg_Inst_ff_SDE_59_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_59_next_state), .CK(clk), .Q(RoundKey[59]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .A(KeyExpansionOutput[60]), .B(
        key[60]), .S(reset), .Z(KeyReg_Inst_ff_SDE_60_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_60_current_state_reg_U1 ( .A(RoundKey[60]), .ZN(
        KeyReg_Inst_ff_SDE_60_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_60_next_state), .CK(clk), .Q(RoundKey[60]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .A(KeyExpansionOutput[61]), .B(
        key[61]), .S(reset), .Z(KeyReg_Inst_ff_SDE_61_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_61_current_state_reg_U1 ( .A(RoundKey[61]), .ZN(
        KeyReg_Inst_ff_SDE_61_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_61_next_state), .CK(clk), .Q(RoundKey[61]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .A(KeyExpansionOutput[62]), .B(
        key[62]), .S(reset), .Z(KeyReg_Inst_ff_SDE_62_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_62_current_state_reg_U1 ( .A(RoundKey[62]), .ZN(
        KeyReg_Inst_ff_SDE_62_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_62_next_state), .CK(clk), .Q(RoundKey[62]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .A(KeyExpansionOutput[63]), .B(
        key[63]), .S(reset), .Z(KeyReg_Inst_ff_SDE_63_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_63_current_state_reg_U1 ( .A(RoundKey[63]), .ZN(
        KeyReg_Inst_ff_SDE_63_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_63_next_state), .CK(clk), .Q(RoundKey[63]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .A(KeyExpansionOutput[64]), .B(
        key[64]), .S(reset), .Z(KeyReg_Inst_ff_SDE_64_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_64_current_state_reg_U1 ( .A(RoundKey[64]), .ZN(
        KeyReg_Inst_ff_SDE_64_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_64_next_state), .CK(clk), .Q(RoundKey[64]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .A(KeyExpansionOutput[65]), .B(
        key[65]), .S(reset), .Z(KeyReg_Inst_ff_SDE_65_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_65_current_state_reg_U1 ( .A(RoundKey[65]), .ZN(
        KeyReg_Inst_ff_SDE_65_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_65_next_state), .CK(clk), .Q(RoundKey[65]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .A(KeyExpansionOutput[66]), .B(
        key[66]), .S(reset), .Z(KeyReg_Inst_ff_SDE_66_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_66_current_state_reg_U1 ( .A(RoundKey[66]), .ZN(
        KeyReg_Inst_ff_SDE_66_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_66_next_state), .CK(clk), .Q(RoundKey[66]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .A(KeyExpansionOutput[67]), .B(
        key[67]), .S(reset), .Z(KeyReg_Inst_ff_SDE_67_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_67_current_state_reg_U1 ( .A(RoundKey[67]), .ZN(
        KeyReg_Inst_ff_SDE_67_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_67_next_state), .CK(clk), .Q(RoundKey[67]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .A(KeyExpansionOutput[68]), .B(
        key[68]), .S(reset), .Z(KeyReg_Inst_ff_SDE_68_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_68_current_state_reg_U1 ( .A(RoundKey[68]), .ZN(
        KeyReg_Inst_ff_SDE_68_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_68_next_state), .CK(clk), .Q(RoundKey[68]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .A(KeyExpansionOutput[69]), .B(
        key[69]), .S(reset), .Z(KeyReg_Inst_ff_SDE_69_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_69_current_state_reg_U1 ( .A(RoundKey[69]), .ZN(
        KeyReg_Inst_ff_SDE_69_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_69_next_state), .CK(clk), .Q(RoundKey[69]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .A(KeyExpansionOutput[70]), .B(
        key[70]), .S(reset), .Z(KeyReg_Inst_ff_SDE_70_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_70_current_state_reg_U1 ( .A(RoundKey[70]), .ZN(
        KeyReg_Inst_ff_SDE_70_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_70_next_state), .CK(clk), .Q(RoundKey[70]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .A(KeyExpansionOutput[71]), .B(
        key[71]), .S(reset), .Z(KeyReg_Inst_ff_SDE_71_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_71_current_state_reg_U1 ( .A(RoundKey[71]), .ZN(
        KeyReg_Inst_ff_SDE_71_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_71_next_state), .CK(clk), .Q(RoundKey[71]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .A(KeyExpansionOutput[72]), .B(
        key[72]), .S(reset), .Z(KeyReg_Inst_ff_SDE_72_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_72_current_state_reg_U1 ( .A(RoundKey[72]), .ZN(
        KeyReg_Inst_ff_SDE_72_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_72_next_state), .CK(clk), .Q(RoundKey[72]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .A(KeyExpansionOutput[73]), .B(
        key[73]), .S(reset), .Z(KeyReg_Inst_ff_SDE_73_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_73_current_state_reg_U1 ( .A(RoundKey[73]), .ZN(
        KeyReg_Inst_ff_SDE_73_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_73_next_state), .CK(clk), .Q(RoundKey[73]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .A(KeyExpansionOutput[74]), .B(
        key[74]), .S(reset), .Z(KeyReg_Inst_ff_SDE_74_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_74_current_state_reg_U1 ( .A(RoundKey[74]), .ZN(
        KeyReg_Inst_ff_SDE_74_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_74_next_state), .CK(clk), .Q(RoundKey[74]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .A(KeyExpansionOutput[75]), .B(
        key[75]), .S(reset), .Z(KeyReg_Inst_ff_SDE_75_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_75_current_state_reg_U1 ( .A(RoundKey[75]), .ZN(
        KeyReg_Inst_ff_SDE_75_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_75_next_state), .CK(clk), .Q(RoundKey[75]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .A(KeyExpansionOutput[76]), .B(
        key[76]), .S(reset), .Z(KeyReg_Inst_ff_SDE_76_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_76_current_state_reg_U1 ( .A(RoundKey[76]), .ZN(
        KeyReg_Inst_ff_SDE_76_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_76_next_state), .CK(clk), .Q(RoundKey[76]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .A(KeyExpansionOutput[77]), .B(
        key[77]), .S(reset), .Z(KeyReg_Inst_ff_SDE_77_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_77_current_state_reg_U1 ( .A(RoundKey[77]), .ZN(
        KeyReg_Inst_ff_SDE_77_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_77_next_state), .CK(clk), .Q(RoundKey[77]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .A(KeyExpansionOutput[78]), .B(
        key[78]), .S(reset), .Z(KeyReg_Inst_ff_SDE_78_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_78_current_state_reg_U1 ( .A(RoundKey[78]), .ZN(
        KeyReg_Inst_ff_SDE_78_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_78_next_state), .CK(clk), .Q(RoundKey[78]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .A(KeyExpansionOutput[79]), .B(
        key[79]), .S(reset), .Z(KeyReg_Inst_ff_SDE_79_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_79_current_state_reg_U1 ( .A(RoundKey[79]), .ZN(
        KeyReg_Inst_ff_SDE_79_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_79_next_state), .CK(clk), .Q(RoundKey[79]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .A(KeyExpansionOutput[80]), .B(
        key[80]), .S(reset), .Z(KeyReg_Inst_ff_SDE_80_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_80_current_state_reg_U1 ( .A(RoundKey[80]), .ZN(
        KeyReg_Inst_ff_SDE_80_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_80_next_state), .CK(clk), .Q(RoundKey[80]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .A(KeyExpansionOutput[81]), .B(
        key[81]), .S(reset), .Z(KeyReg_Inst_ff_SDE_81_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_81_current_state_reg_U1 ( .A(RoundKey[81]), .ZN(
        KeyReg_Inst_ff_SDE_81_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_81_next_state), .CK(clk), .Q(RoundKey[81]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .A(KeyExpansionOutput[82]), .B(
        key[82]), .S(reset), .Z(KeyReg_Inst_ff_SDE_82_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_82_current_state_reg_U1 ( .A(RoundKey[82]), .ZN(
        KeyReg_Inst_ff_SDE_82_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_82_next_state), .CK(clk), .Q(RoundKey[82]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .A(KeyExpansionOutput[83]), .B(
        key[83]), .S(reset), .Z(KeyReg_Inst_ff_SDE_83_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_83_current_state_reg_U1 ( .A(RoundKey[83]), .ZN(
        KeyReg_Inst_ff_SDE_83_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_83_next_state), .CK(clk), .Q(RoundKey[83]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .A(KeyExpansionOutput[84]), .B(
        key[84]), .S(reset), .Z(KeyReg_Inst_ff_SDE_84_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_84_current_state_reg_U1 ( .A(RoundKey[84]), .ZN(
        KeyReg_Inst_ff_SDE_84_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_84_next_state), .CK(clk), .Q(RoundKey[84]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .A(KeyExpansionOutput[85]), .B(
        key[85]), .S(reset), .Z(KeyReg_Inst_ff_SDE_85_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_85_current_state_reg_U1 ( .A(RoundKey[85]), .ZN(
        KeyReg_Inst_ff_SDE_85_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_85_next_state), .CK(clk), .Q(RoundKey[85]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .A(KeyExpansionOutput[86]), .B(
        key[86]), .S(reset), .Z(KeyReg_Inst_ff_SDE_86_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_86_current_state_reg_U1 ( .A(RoundKey[86]), .ZN(
        KeyReg_Inst_ff_SDE_86_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_86_next_state), .CK(clk), .Q(RoundKey[86]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .A(KeyExpansionOutput[87]), .B(
        key[87]), .S(reset), .Z(KeyReg_Inst_ff_SDE_87_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_87_current_state_reg_U1 ( .A(RoundKey[87]), .ZN(
        KeyReg_Inst_ff_SDE_87_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_87_next_state), .CK(clk), .Q(RoundKey[87]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .A(KeyExpansionOutput[88]), .B(
        key[88]), .S(reset), .Z(KeyReg_Inst_ff_SDE_88_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_88_current_state_reg_U1 ( .A(RoundKey[88]), .ZN(
        KeyReg_Inst_ff_SDE_88_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_88_next_state), .CK(clk), .Q(RoundKey[88]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .A(KeyExpansionOutput[89]), .B(
        key[89]), .S(reset), .Z(KeyReg_Inst_ff_SDE_89_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_89_current_state_reg_U1 ( .A(RoundKey[89]), .ZN(
        KeyReg_Inst_ff_SDE_89_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_89_next_state), .CK(clk), .Q(RoundKey[89]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .A(KeyExpansionOutput[90]), .B(
        key[90]), .S(reset), .Z(KeyReg_Inst_ff_SDE_90_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_90_current_state_reg_U1 ( .A(RoundKey[90]), .ZN(
        KeyReg_Inst_ff_SDE_90_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_90_next_state), .CK(clk), .Q(RoundKey[90]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .A(KeyExpansionOutput[91]), .B(
        key[91]), .S(reset), .Z(KeyReg_Inst_ff_SDE_91_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_91_current_state_reg_U1 ( .A(RoundKey[91]), .ZN(
        KeyReg_Inst_ff_SDE_91_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_91_next_state), .CK(clk), .Q(RoundKey[91]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .A(KeyExpansionOutput[92]), .B(
        key[92]), .S(reset), .Z(KeyReg_Inst_ff_SDE_92_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_92_current_state_reg_U1 ( .A(RoundKey[92]), .ZN(
        KeyReg_Inst_ff_SDE_92_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_92_next_state), .CK(clk), .Q(RoundKey[92]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .A(KeyExpansionOutput[93]), .B(
        key[93]), .S(reset), .Z(KeyReg_Inst_ff_SDE_93_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_93_current_state_reg_U1 ( .A(RoundKey[93]), .ZN(
        KeyReg_Inst_ff_SDE_93_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_93_next_state), .CK(clk), .Q(RoundKey[93]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .A(KeyExpansionOutput[94]), .B(
        key[94]), .S(reset), .Z(KeyReg_Inst_ff_SDE_94_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_94_current_state_reg_U1 ( .A(RoundKey[94]), .ZN(
        KeyReg_Inst_ff_SDE_94_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_94_next_state), .CK(clk), .Q(RoundKey[94]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .A(KeyExpansionOutput[95]), .B(
        key[95]), .S(reset), .Z(KeyReg_Inst_ff_SDE_95_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_95_current_state_reg_U1 ( .A(RoundKey[95]), .ZN(
        KeyReg_Inst_ff_SDE_95_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_95_next_state), .CK(clk), .Q(RoundKey[95]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .A(KeyExpansionOutput[96]), .B(
        key[96]), .S(reset), .Z(KeyReg_Inst_ff_SDE_96_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_96_current_state_reg_U1 ( .A(RoundKey[96]), .ZN(
        KeyReg_Inst_ff_SDE_96_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_96_next_state), .CK(clk), .Q(RoundKey[96]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .A(KeyExpansionOutput[97]), .B(
        key[97]), .S(reset), .Z(KeyReg_Inst_ff_SDE_97_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_97_current_state_reg_U1 ( .A(RoundKey[97]), .ZN(
        KeyReg_Inst_ff_SDE_97_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_97_next_state), .CK(clk), .Q(RoundKey[97]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .A(KeyExpansionOutput[98]), .B(
        key[98]), .S(reset), .Z(KeyReg_Inst_ff_SDE_98_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_98_current_state_reg_U1 ( .A(RoundKey[98]), .ZN(
        KeyReg_Inst_ff_SDE_98_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_98_next_state), .CK(clk), .Q(RoundKey[98]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .A(KeyExpansionOutput[99]), .B(
        key[99]), .S(reset), .Z(KeyReg_Inst_ff_SDE_99_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_99_current_state_reg_U1 ( .A(RoundKey[99]), .ZN(
        KeyReg_Inst_ff_SDE_99_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_99_next_state), .CK(clk), .Q(RoundKey[99]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .A(KeyExpansionOutput[100]), 
        .B(key[100]), .S(reset), .Z(KeyReg_Inst_ff_SDE_100_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_100_current_state_reg_U1 ( .A(RoundKey[100]), .ZN(
        KeyReg_Inst_ff_SDE_100_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_100_next_state), .CK(clk), .Q(RoundKey[100]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .A(KeyExpansionOutput[101]), 
        .B(key[101]), .S(reset), .Z(KeyReg_Inst_ff_SDE_101_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_101_current_state_reg_U1 ( .A(RoundKey[101]), .ZN(
        KeyReg_Inst_ff_SDE_101_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_101_next_state), .CK(clk), .Q(RoundKey[101]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .A(KeyExpansionOutput[102]), 
        .B(key[102]), .S(reset), .Z(KeyReg_Inst_ff_SDE_102_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_102_current_state_reg_U1 ( .A(RoundKey[102]), .ZN(
        KeyReg_Inst_ff_SDE_102_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_102_next_state), .CK(clk), .Q(RoundKey[102]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .A(KeyExpansionOutput[103]), 
        .B(key[103]), .S(reset), .Z(KeyReg_Inst_ff_SDE_103_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_103_current_state_reg_U1 ( .A(RoundKey[103]), .ZN(
        KeyReg_Inst_ff_SDE_103_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_103_next_state), .CK(clk), .Q(RoundKey[103]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .A(KeyExpansionOutput[104]), 
        .B(key[104]), .S(reset), .Z(KeyReg_Inst_ff_SDE_104_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_104_current_state_reg_U1 ( .A(RoundKey[104]), .ZN(
        KeyReg_Inst_ff_SDE_104_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_104_next_state), .CK(clk), .Q(RoundKey[104]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .A(KeyExpansionOutput[105]), 
        .B(key[105]), .S(reset), .Z(KeyReg_Inst_ff_SDE_105_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_105_current_state_reg_U1 ( .A(RoundKey[105]), .ZN(
        KeyReg_Inst_ff_SDE_105_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_105_next_state), .CK(clk), .Q(RoundKey[105]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .A(KeyExpansionOutput[106]), 
        .B(key[106]), .S(reset), .Z(KeyReg_Inst_ff_SDE_106_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_106_current_state_reg_U1 ( .A(RoundKey[106]), .ZN(
        KeyReg_Inst_ff_SDE_106_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_106_next_state), .CK(clk), .Q(RoundKey[106]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .A(KeyExpansionOutput[107]), 
        .B(key[107]), .S(reset), .Z(KeyReg_Inst_ff_SDE_107_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_107_current_state_reg_U1 ( .A(RoundKey[107]), .ZN(
        KeyReg_Inst_ff_SDE_107_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_107_next_state), .CK(clk), .Q(RoundKey[107]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .A(KeyExpansionOutput[108]), 
        .B(key[108]), .S(reset), .Z(KeyReg_Inst_ff_SDE_108_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_108_current_state_reg_U1 ( .A(RoundKey[108]), .ZN(
        KeyReg_Inst_ff_SDE_108_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_108_next_state), .CK(clk), .Q(RoundKey[108]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .A(KeyExpansionOutput[109]), 
        .B(key[109]), .S(reset), .Z(KeyReg_Inst_ff_SDE_109_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_109_current_state_reg_U1 ( .A(RoundKey[109]), .ZN(
        KeyReg_Inst_ff_SDE_109_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_109_next_state), .CK(clk), .Q(RoundKey[109]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .A(KeyExpansionOutput[110]), 
        .B(key[110]), .S(reset), .Z(KeyReg_Inst_ff_SDE_110_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_110_current_state_reg_U1 ( .A(RoundKey[110]), .ZN(
        KeyReg_Inst_ff_SDE_110_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_110_next_state), .CK(clk), .Q(RoundKey[110]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .A(KeyExpansionOutput[111]), 
        .B(key[111]), .S(reset), .Z(KeyReg_Inst_ff_SDE_111_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_111_current_state_reg_U1 ( .A(RoundKey[111]), .ZN(
        KeyReg_Inst_ff_SDE_111_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_111_next_state), .CK(clk), .Q(RoundKey[111]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .A(KeyExpansionOutput[112]), 
        .B(key[112]), .S(reset), .Z(KeyReg_Inst_ff_SDE_112_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_112_current_state_reg_U1 ( .A(RoundKey[112]), .ZN(
        KeyReg_Inst_ff_SDE_112_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_112_next_state), .CK(clk), .Q(RoundKey[112]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .A(KeyExpansionOutput[113]), 
        .B(key[113]), .S(reset), .Z(KeyReg_Inst_ff_SDE_113_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_113_current_state_reg_U1 ( .A(RoundKey[113]), .ZN(
        KeyReg_Inst_ff_SDE_113_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_113_next_state), .CK(clk), .Q(RoundKey[113]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .A(KeyExpansionOutput[114]), 
        .B(key[114]), .S(reset), .Z(KeyReg_Inst_ff_SDE_114_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_114_current_state_reg_U1 ( .A(RoundKey[114]), .ZN(
        KeyReg_Inst_ff_SDE_114_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_114_next_state), .CK(clk), .Q(RoundKey[114]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .A(KeyExpansionOutput[115]), 
        .B(key[115]), .S(reset), .Z(KeyReg_Inst_ff_SDE_115_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_115_current_state_reg_U1 ( .A(RoundKey[115]), .ZN(
        KeyReg_Inst_ff_SDE_115_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_115_next_state), .CK(clk), .Q(RoundKey[115]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .A(KeyExpansionOutput[116]), 
        .B(key[116]), .S(reset), .Z(KeyReg_Inst_ff_SDE_116_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_116_current_state_reg_U1 ( .A(RoundKey[116]), .ZN(
        KeyReg_Inst_ff_SDE_116_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_116_next_state), .CK(clk), .Q(RoundKey[116]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .A(KeyExpansionOutput[117]), 
        .B(key[117]), .S(reset), .Z(KeyReg_Inst_ff_SDE_117_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_117_current_state_reg_U1 ( .A(RoundKey[117]), .ZN(
        KeyReg_Inst_ff_SDE_117_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_117_next_state), .CK(clk), .Q(RoundKey[117]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .A(KeyExpansionOutput[118]), 
        .B(key[118]), .S(reset), .Z(KeyReg_Inst_ff_SDE_118_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_118_current_state_reg_U1 ( .A(RoundKey[118]), .ZN(
        KeyReg_Inst_ff_SDE_118_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_118_next_state), .CK(clk), .Q(RoundKey[118]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .A(KeyExpansionOutput[119]), 
        .B(key[119]), .S(reset), .Z(KeyReg_Inst_ff_SDE_119_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_119_current_state_reg_U1 ( .A(RoundKey[119]), .ZN(
        KeyReg_Inst_ff_SDE_119_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_119_next_state), .CK(clk), .Q(RoundKey[119]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .A(KeyExpansionOutput[120]), 
        .B(key[120]), .S(reset), .Z(KeyReg_Inst_ff_SDE_120_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_120_current_state_reg_U1 ( .A(RoundKey[120]), .ZN(
        KeyReg_Inst_ff_SDE_120_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_120_next_state), .CK(clk), .Q(RoundKey[120]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .A(KeyExpansionOutput[121]), 
        .B(key[121]), .S(reset), .Z(KeyReg_Inst_ff_SDE_121_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_121_current_state_reg_U1 ( .A(RoundKey[121]), .ZN(
        KeyReg_Inst_ff_SDE_121_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_121_next_state), .CK(clk), .Q(RoundKey[121]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .A(KeyExpansionOutput[122]), 
        .B(key[122]), .S(reset), .Z(KeyReg_Inst_ff_SDE_122_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_122_current_state_reg_U1 ( .A(RoundKey[122]), .ZN(
        KeyReg_Inst_ff_SDE_122_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_122_next_state), .CK(clk), .Q(RoundKey[122]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .A(KeyExpansionOutput[123]), 
        .B(key[123]), .S(reset), .Z(KeyReg_Inst_ff_SDE_123_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_123_current_state_reg_U1 ( .A(RoundKey[123]), .ZN(
        KeyReg_Inst_ff_SDE_123_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_123_next_state), .CK(clk), .Q(RoundKey[123]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .A(KeyExpansionOutput[124]), 
        .B(key[124]), .S(reset), .Z(KeyReg_Inst_ff_SDE_124_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_124_current_state_reg_U1 ( .A(RoundKey[124]), .ZN(
        KeyReg_Inst_ff_SDE_124_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_124_next_state), .CK(clk), .Q(RoundKey[124]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .A(KeyExpansionOutput[125]), 
        .B(key[125]), .S(reset), .Z(KeyReg_Inst_ff_SDE_125_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_125_current_state_reg_U1 ( .A(RoundKey[125]), .ZN(
        KeyReg_Inst_ff_SDE_125_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_125_next_state), .CK(clk), .Q(RoundKey[125]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .A(KeyExpansionOutput[126]), 
        .B(key[126]), .S(reset), .Z(KeyReg_Inst_ff_SDE_126_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_126_current_state_reg_U1 ( .A(RoundKey[126]), .ZN(
        KeyReg_Inst_ff_SDE_126_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_126_next_state), .CK(clk), .Q(RoundKey[126]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .A(KeyExpansionOutput[127]), 
        .B(key[127]), .S(reset), .Z(KeyReg_Inst_ff_SDE_127_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_127_current_state_reg_U1 ( .A(RoundKey[127]), .ZN(
        KeyReg_Inst_ff_SDE_127_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_127_next_state), .CK(clk), .Q(RoundKey[127]), .QN()
         );
  XOR2_X1 KeyExpansionIns_U128 ( .A(RoundKey[9]), .B(KeyExpansionOutput[41]), 
        .Z(KeyExpansionOutput[9]) );
  XOR2_X1 KeyExpansionIns_U127 ( .A(RoundKey[8]), .B(KeyExpansionOutput[40]), 
        .Z(KeyExpansionOutput[8]) );
  XOR2_X1 KeyExpansionIns_U126 ( .A(RoundKey[7]), .B(KeyExpansionOutput[39]), 
        .Z(KeyExpansionOutput[7]) );
  XOR2_X1 KeyExpansionIns_U125 ( .A(RoundKey[6]), .B(KeyExpansionOutput[38]), 
        .Z(KeyExpansionOutput[6]) );
  XOR2_X1 KeyExpansionIns_U124 ( .A(RoundKey[5]), .B(KeyExpansionOutput[37]), 
        .Z(KeyExpansionOutput[5]) );
  XOR2_X1 KeyExpansionIns_U123 ( .A(RoundKey[4]), .B(KeyExpansionOutput[36]), 
        .Z(KeyExpansionOutput[4]) );
  XOR2_X1 KeyExpansionIns_U122 ( .A(RoundKey[41]), .B(KeyExpansionOutput[73]), 
        .Z(KeyExpansionOutput[41]) );
  XOR2_X1 KeyExpansionIns_U121 ( .A(RoundKey[73]), .B(KeyExpansionOutput[105]), 
        .Z(KeyExpansionOutput[73]) );
  XOR2_X1 KeyExpansionIns_U120 ( .A(RoundKey[40]), .B(KeyExpansionOutput[72]), 
        .Z(KeyExpansionOutput[40]) );
  XOR2_X1 KeyExpansionIns_U119 ( .A(RoundKey[72]), .B(KeyExpansionOutput[104]), 
        .Z(KeyExpansionOutput[72]) );
  XOR2_X1 KeyExpansionIns_U118 ( .A(RoundKey[3]), .B(KeyExpansionOutput[35]), 
        .Z(KeyExpansionOutput[3]) );
  XOR2_X1 KeyExpansionIns_U117 ( .A(RoundKey[39]), .B(KeyExpansionOutput[71]), 
        .Z(KeyExpansionOutput[39]) );
  XOR2_X1 KeyExpansionIns_U116 ( .A(RoundKey[71]), .B(KeyExpansionOutput[103]), 
        .Z(KeyExpansionOutput[71]) );
  XOR2_X1 KeyExpansionIns_U115 ( .A(RoundKey[38]), .B(KeyExpansionOutput[70]), 
        .Z(KeyExpansionOutput[38]) );
  XOR2_X1 KeyExpansionIns_U114 ( .A(RoundKey[70]), .B(KeyExpansionOutput[102]), 
        .Z(KeyExpansionOutput[70]) );
  XOR2_X1 KeyExpansionIns_U113 ( .A(RoundKey[37]), .B(KeyExpansionOutput[69]), 
        .Z(KeyExpansionOutput[37]) );
  XOR2_X1 KeyExpansionIns_U112 ( .A(RoundKey[69]), .B(KeyExpansionOutput[101]), 
        .Z(KeyExpansionOutput[69]) );
  XOR2_X1 KeyExpansionIns_U111 ( .A(RoundKey[36]), .B(KeyExpansionOutput[68]), 
        .Z(KeyExpansionOutput[36]) );
  XOR2_X1 KeyExpansionIns_U110 ( .A(RoundKey[68]), .B(KeyExpansionOutput[100]), 
        .Z(KeyExpansionOutput[68]) );
  XOR2_X1 KeyExpansionIns_U109 ( .A(RoundKey[35]), .B(KeyExpansionOutput[67]), 
        .Z(KeyExpansionOutput[35]) );
  XOR2_X1 KeyExpansionIns_U108 ( .A(RoundKey[67]), .B(KeyExpansionOutput[99]), 
        .Z(KeyExpansionOutput[67]) );
  XOR2_X1 KeyExpansionIns_U107 ( .A(RoundKey[99]), .B(KeyExpansionIns_tmp[3]), 
        .Z(KeyExpansionOutput[99]) );
  XOR2_X1 KeyExpansionIns_U106 ( .A(RoundKey[31]), .B(KeyExpansionOutput[63]), 
        .Z(KeyExpansionOutput[31]) );
  XOR2_X1 KeyExpansionIns_U105 ( .A(RoundKey[63]), .B(KeyExpansionOutput[95]), 
        .Z(KeyExpansionOutput[63]) );
  XOR2_X1 KeyExpansionIns_U104 ( .A(RoundKey[95]), .B(KeyExpansionOutput[127]), 
        .Z(KeyExpansionOutput[95]) );
  XOR2_X1 KeyExpansionIns_U103 ( .A(RoundKey[30]), .B(KeyExpansionOutput[62]), 
        .Z(KeyExpansionOutput[30]) );
  XOR2_X1 KeyExpansionIns_U102 ( .A(RoundKey[62]), .B(KeyExpansionOutput[94]), 
        .Z(KeyExpansionOutput[62]) );
  XOR2_X1 KeyExpansionIns_U101 ( .A(RoundKey[94]), .B(KeyExpansionOutput[126]), 
        .Z(KeyExpansionOutput[94]) );
  XOR2_X1 KeyExpansionIns_U100 ( .A(RoundKey[2]), .B(KeyExpansionOutput[34]), 
        .Z(KeyExpansionOutput[2]) );
  XOR2_X1 KeyExpansionIns_U99 ( .A(RoundKey[34]), .B(KeyExpansionOutput[66]), 
        .Z(KeyExpansionOutput[34]) );
  XOR2_X1 KeyExpansionIns_U98 ( .A(RoundKey[66]), .B(KeyExpansionOutput[98]), 
        .Z(KeyExpansionOutput[66]) );
  XOR2_X1 KeyExpansionIns_U97 ( .A(RoundKey[98]), .B(KeyExpansionIns_tmp[2]), 
        .Z(KeyExpansionOutput[98]) );
  XOR2_X1 KeyExpansionIns_U96 ( .A(RoundKey[29]), .B(KeyExpansionOutput[61]), 
        .Z(KeyExpansionOutput[29]) );
  XOR2_X1 KeyExpansionIns_U95 ( .A(RoundKey[61]), .B(KeyExpansionOutput[93]), 
        .Z(KeyExpansionOutput[61]) );
  XOR2_X1 KeyExpansionIns_U94 ( .A(RoundKey[93]), .B(KeyExpansionOutput[125]), 
        .Z(KeyExpansionOutput[93]) );
  XOR2_X1 KeyExpansionIns_U93 ( .A(RoundKey[28]), .B(KeyExpansionOutput[60]), 
        .Z(KeyExpansionOutput[28]) );
  XOR2_X1 KeyExpansionIns_U92 ( .A(RoundKey[60]), .B(KeyExpansionOutput[92]), 
        .Z(KeyExpansionOutput[60]) );
  XOR2_X1 KeyExpansionIns_U91 ( .A(RoundKey[92]), .B(KeyExpansionOutput[124]), 
        .Z(KeyExpansionOutput[92]) );
  XOR2_X1 KeyExpansionIns_U90 ( .A(RoundKey[27]), .B(KeyExpansionOutput[59]), 
        .Z(KeyExpansionOutput[27]) );
  XOR2_X1 KeyExpansionIns_U89 ( .A(RoundKey[59]), .B(KeyExpansionOutput[91]), 
        .Z(KeyExpansionOutput[59]) );
  XOR2_X1 KeyExpansionIns_U88 ( .A(RoundKey[91]), .B(KeyExpansionOutput[123]), 
        .Z(KeyExpansionOutput[91]) );
  XOR2_X1 KeyExpansionIns_U87 ( .A(RoundKey[26]), .B(KeyExpansionOutput[58]), 
        .Z(KeyExpansionOutput[26]) );
  XOR2_X1 KeyExpansionIns_U86 ( .A(RoundKey[58]), .B(KeyExpansionOutput[90]), 
        .Z(KeyExpansionOutput[58]) );
  XOR2_X1 KeyExpansionIns_U85 ( .A(RoundKey[90]), .B(KeyExpansionOutput[122]), 
        .Z(KeyExpansionOutput[90]) );
  XOR2_X1 KeyExpansionIns_U84 ( .A(RoundKey[25]), .B(KeyExpansionOutput[57]), 
        .Z(KeyExpansionOutput[25]) );
  XOR2_X1 KeyExpansionIns_U83 ( .A(RoundKey[57]), .B(KeyExpansionOutput[89]), 
        .Z(KeyExpansionOutput[57]) );
  XOR2_X1 KeyExpansionIns_U82 ( .A(RoundKey[89]), .B(KeyExpansionOutput[121]), 
        .Z(KeyExpansionOutput[89]) );
  XOR2_X1 KeyExpansionIns_U81 ( .A(RoundKey[24]), .B(KeyExpansionOutput[56]), 
        .Z(KeyExpansionOutput[24]) );
  XOR2_X1 KeyExpansionIns_U80 ( .A(RoundKey[56]), .B(KeyExpansionOutput[88]), 
        .Z(KeyExpansionOutput[56]) );
  XOR2_X1 KeyExpansionIns_U79 ( .A(RoundKey[88]), .B(KeyExpansionOutput[120]), 
        .Z(KeyExpansionOutput[88]) );
  XOR2_X1 KeyExpansionIns_U78 ( .A(RoundKey[23]), .B(KeyExpansionOutput[55]), 
        .Z(KeyExpansionOutput[23]) );
  XOR2_X1 KeyExpansionIns_U77 ( .A(RoundKey[55]), .B(KeyExpansionOutput[87]), 
        .Z(KeyExpansionOutput[55]) );
  XOR2_X1 KeyExpansionIns_U76 ( .A(RoundKey[87]), .B(KeyExpansionOutput[119]), 
        .Z(KeyExpansionOutput[87]) );
  XOR2_X1 KeyExpansionIns_U75 ( .A(RoundKey[22]), .B(KeyExpansionOutput[54]), 
        .Z(KeyExpansionOutput[22]) );
  XOR2_X1 KeyExpansionIns_U74 ( .A(RoundKey[54]), .B(KeyExpansionOutput[86]), 
        .Z(KeyExpansionOutput[54]) );
  XOR2_X1 KeyExpansionIns_U73 ( .A(RoundKey[86]), .B(KeyExpansionOutput[118]), 
        .Z(KeyExpansionOutput[86]) );
  XOR2_X1 KeyExpansionIns_U72 ( .A(RoundKey[21]), .B(KeyExpansionOutput[53]), 
        .Z(KeyExpansionOutput[21]) );
  XOR2_X1 KeyExpansionIns_U71 ( .A(RoundKey[53]), .B(KeyExpansionOutput[85]), 
        .Z(KeyExpansionOutput[53]) );
  XOR2_X1 KeyExpansionIns_U70 ( .A(RoundKey[85]), .B(KeyExpansionOutput[117]), 
        .Z(KeyExpansionOutput[85]) );
  XOR2_X1 KeyExpansionIns_U69 ( .A(RoundKey[20]), .B(KeyExpansionOutput[52]), 
        .Z(KeyExpansionOutput[20]) );
  XOR2_X1 KeyExpansionIns_U68 ( .A(RoundKey[52]), .B(KeyExpansionOutput[84]), 
        .Z(KeyExpansionOutput[52]) );
  XOR2_X1 KeyExpansionIns_U67 ( .A(RoundKey[84]), .B(KeyExpansionOutput[116]), 
        .Z(KeyExpansionOutput[84]) );
  XOR2_X1 KeyExpansionIns_U66 ( .A(RoundKey[1]), .B(KeyExpansionOutput[33]), 
        .Z(KeyExpansionOutput[1]) );
  XOR2_X1 KeyExpansionIns_U65 ( .A(RoundKey[33]), .B(KeyExpansionOutput[65]), 
        .Z(KeyExpansionOutput[33]) );
  XOR2_X1 KeyExpansionIns_U64 ( .A(RoundKey[65]), .B(KeyExpansionOutput[97]), 
        .Z(KeyExpansionOutput[65]) );
  XOR2_X1 KeyExpansionIns_U63 ( .A(RoundKey[97]), .B(KeyExpansionIns_tmp[1]), 
        .Z(KeyExpansionOutput[97]) );
  XOR2_X1 KeyExpansionIns_U62 ( .A(RoundKey[19]), .B(KeyExpansionOutput[51]), 
        .Z(KeyExpansionOutput[19]) );
  XOR2_X1 KeyExpansionIns_U61 ( .A(RoundKey[51]), .B(KeyExpansionOutput[83]), 
        .Z(KeyExpansionOutput[51]) );
  XOR2_X1 KeyExpansionIns_U60 ( .A(RoundKey[83]), .B(KeyExpansionOutput[115]), 
        .Z(KeyExpansionOutput[83]) );
  XOR2_X1 KeyExpansionIns_U59 ( .A(RoundKey[18]), .B(KeyExpansionOutput[50]), 
        .Z(KeyExpansionOutput[18]) );
  XOR2_X1 KeyExpansionIns_U58 ( .A(RoundKey[50]), .B(KeyExpansionOutput[82]), 
        .Z(KeyExpansionOutput[50]) );
  XOR2_X1 KeyExpansionIns_U57 ( .A(RoundKey[82]), .B(KeyExpansionOutput[114]), 
        .Z(KeyExpansionOutput[82]) );
  XOR2_X1 KeyExpansionIns_U56 ( .A(RoundKey[17]), .B(KeyExpansionOutput[49]), 
        .Z(KeyExpansionOutput[17]) );
  XOR2_X1 KeyExpansionIns_U55 ( .A(RoundKey[49]), .B(KeyExpansionOutput[81]), 
        .Z(KeyExpansionOutput[49]) );
  XOR2_X1 KeyExpansionIns_U54 ( .A(RoundKey[81]), .B(KeyExpansionOutput[113]), 
        .Z(KeyExpansionOutput[81]) );
  XOR2_X1 KeyExpansionIns_U53 ( .A(RoundKey[16]), .B(KeyExpansionOutput[48]), 
        .Z(KeyExpansionOutput[16]) );
  XOR2_X1 KeyExpansionIns_U52 ( .A(RoundKey[48]), .B(KeyExpansionOutput[80]), 
        .Z(KeyExpansionOutput[48]) );
  XOR2_X1 KeyExpansionIns_U51 ( .A(RoundKey[80]), .B(KeyExpansionOutput[112]), 
        .Z(KeyExpansionOutput[80]) );
  XOR2_X1 KeyExpansionIns_U50 ( .A(RoundKey[15]), .B(KeyExpansionOutput[47]), 
        .Z(KeyExpansionOutput[15]) );
  XOR2_X1 KeyExpansionIns_U49 ( .A(RoundKey[47]), .B(KeyExpansionOutput[79]), 
        .Z(KeyExpansionOutput[47]) );
  XOR2_X1 KeyExpansionIns_U48 ( .A(RoundKey[79]), .B(KeyExpansionOutput[111]), 
        .Z(KeyExpansionOutput[79]) );
  XOR2_X1 KeyExpansionIns_U47 ( .A(RoundKey[14]), .B(KeyExpansionOutput[46]), 
        .Z(KeyExpansionOutput[14]) );
  XOR2_X1 KeyExpansionIns_U46 ( .A(RoundKey[46]), .B(KeyExpansionOutput[78]), 
        .Z(KeyExpansionOutput[46]) );
  XOR2_X1 KeyExpansionIns_U45 ( .A(RoundKey[78]), .B(KeyExpansionOutput[110]), 
        .Z(KeyExpansionOutput[78]) );
  XOR2_X1 KeyExpansionIns_U44 ( .A(RoundKey[13]), .B(KeyExpansionOutput[45]), 
        .Z(KeyExpansionOutput[13]) );
  XOR2_X1 KeyExpansionIns_U43 ( .A(RoundKey[45]), .B(KeyExpansionOutput[77]), 
        .Z(KeyExpansionOutput[45]) );
  XOR2_X1 KeyExpansionIns_U42 ( .A(RoundKey[77]), .B(KeyExpansionOutput[109]), 
        .Z(KeyExpansionOutput[77]) );
  XOR2_X1 KeyExpansionIns_U41 ( .A(RoundKey[12]), .B(KeyExpansionOutput[44]), 
        .Z(KeyExpansionOutput[12]) );
  XOR2_X1 KeyExpansionIns_U40 ( .A(RoundKey[44]), .B(KeyExpansionOutput[76]), 
        .Z(KeyExpansionOutput[44]) );
  XOR2_X1 KeyExpansionIns_U39 ( .A(RoundKey[76]), .B(KeyExpansionOutput[108]), 
        .Z(KeyExpansionOutput[76]) );
  XOR2_X1 KeyExpansionIns_U38 ( .A(RoundKey[127]), .B(KeyExpansionIns_tmp[31]), 
        .Z(KeyExpansionOutput[127]) );
  XOR2_X1 KeyExpansionIns_U37 ( .A(RoundKey[126]), .B(KeyExpansionIns_tmp[30]), 
        .Z(KeyExpansionOutput[126]) );
  XOR2_X1 KeyExpansionIns_U36 ( .A(RoundKey[125]), .B(KeyExpansionIns_tmp[29]), 
        .Z(KeyExpansionOutput[125]) );
  XOR2_X1 KeyExpansionIns_U35 ( .A(RoundKey[124]), .B(KeyExpansionIns_tmp[28]), 
        .Z(KeyExpansionOutput[124]) );
  XOR2_X1 KeyExpansionIns_U34 ( .A(RoundKey[123]), .B(KeyExpansionIns_tmp[27]), 
        .Z(KeyExpansionOutput[123]) );
  XOR2_X1 KeyExpansionIns_U33 ( .A(RoundKey[122]), .B(KeyExpansionIns_tmp[26]), 
        .Z(KeyExpansionOutput[122]) );
  XOR2_X1 KeyExpansionIns_U32 ( .A(RoundKey[121]), .B(KeyExpansionIns_tmp[25]), 
        .Z(KeyExpansionOutput[121]) );
  XOR2_X1 KeyExpansionIns_U31 ( .A(RoundKey[120]), .B(KeyExpansionIns_tmp[24]), 
        .Z(KeyExpansionOutput[120]) );
  XOR2_X1 KeyExpansionIns_U30 ( .A(RoundKey[11]), .B(KeyExpansionOutput[43]), 
        .Z(KeyExpansionOutput[11]) );
  XOR2_X1 KeyExpansionIns_U29 ( .A(RoundKey[43]), .B(KeyExpansionOutput[75]), 
        .Z(KeyExpansionOutput[43]) );
  XOR2_X1 KeyExpansionIns_U28 ( .A(RoundKey[75]), .B(KeyExpansionOutput[107]), 
        .Z(KeyExpansionOutput[75]) );
  XOR2_X1 KeyExpansionIns_U27 ( .A(RoundKey[119]), .B(KeyExpansionIns_tmp[23]), 
        .Z(KeyExpansionOutput[119]) );
  XOR2_X1 KeyExpansionIns_U26 ( .A(RoundKey[118]), .B(KeyExpansionIns_tmp[22]), 
        .Z(KeyExpansionOutput[118]) );
  XOR2_X1 KeyExpansionIns_U25 ( .A(RoundKey[117]), .B(KeyExpansionIns_tmp[21]), 
        .Z(KeyExpansionOutput[117]) );
  XOR2_X1 KeyExpansionIns_U24 ( .A(RoundKey[116]), .B(KeyExpansionIns_tmp[20]), 
        .Z(KeyExpansionOutput[116]) );
  XOR2_X1 KeyExpansionIns_U23 ( .A(RoundKey[115]), .B(KeyExpansionIns_tmp[19]), 
        .Z(KeyExpansionOutput[115]) );
  XOR2_X1 KeyExpansionIns_U22 ( .A(RoundKey[114]), .B(KeyExpansionIns_tmp[18]), 
        .Z(KeyExpansionOutput[114]) );
  XOR2_X1 KeyExpansionIns_U21 ( .A(RoundKey[113]), .B(KeyExpansionIns_tmp[17]), 
        .Z(KeyExpansionOutput[113]) );
  XOR2_X1 KeyExpansionIns_U20 ( .A(RoundKey[112]), .B(KeyExpansionIns_tmp[16]), 
        .Z(KeyExpansionOutput[112]) );
  XOR2_X1 KeyExpansionIns_U19 ( .A(RoundKey[111]), .B(KeyExpansionIns_tmp[15]), 
        .Z(KeyExpansionOutput[111]) );
  XOR2_X1 KeyExpansionIns_U18 ( .A(RoundKey[110]), .B(KeyExpansionIns_tmp[14]), 
        .Z(KeyExpansionOutput[110]) );
  XOR2_X1 KeyExpansionIns_U17 ( .A(RoundKey[10]), .B(KeyExpansionOutput[42]), 
        .Z(KeyExpansionOutput[10]) );
  XOR2_X1 KeyExpansionIns_U16 ( .A(RoundKey[42]), .B(KeyExpansionOutput[74]), 
        .Z(KeyExpansionOutput[42]) );
  XOR2_X1 KeyExpansionIns_U15 ( .A(RoundKey[74]), .B(KeyExpansionOutput[106]), 
        .Z(KeyExpansionOutput[74]) );
  XOR2_X1 KeyExpansionIns_U14 ( .A(RoundKey[109]), .B(KeyExpansionIns_tmp[13]), 
        .Z(KeyExpansionOutput[109]) );
  XOR2_X1 KeyExpansionIns_U13 ( .A(RoundKey[108]), .B(KeyExpansionIns_tmp[12]), 
        .Z(KeyExpansionOutput[108]) );
  XOR2_X1 KeyExpansionIns_U12 ( .A(RoundKey[107]), .B(KeyExpansionIns_tmp[11]), 
        .Z(KeyExpansionOutput[107]) );
  XOR2_X1 KeyExpansionIns_U11 ( .A(RoundKey[106]), .B(KeyExpansionIns_tmp[10]), 
        .Z(KeyExpansionOutput[106]) );
  XOR2_X1 KeyExpansionIns_U10 ( .A(RoundKey[105]), .B(KeyExpansionIns_tmp[9]), 
        .Z(KeyExpansionOutput[105]) );
  XOR2_X1 KeyExpansionIns_U9 ( .A(RoundKey[104]), .B(KeyExpansionIns_tmp[8]), 
        .Z(KeyExpansionOutput[104]) );
  XOR2_X1 KeyExpansionIns_U8 ( .A(RoundKey[103]), .B(KeyExpansionIns_tmp[7]), 
        .Z(KeyExpansionOutput[103]) );
  XOR2_X1 KeyExpansionIns_U7 ( .A(RoundKey[102]), .B(KeyExpansionIns_tmp[6]), 
        .Z(KeyExpansionOutput[102]) );
  XOR2_X1 KeyExpansionIns_U6 ( .A(RoundKey[101]), .B(KeyExpansionIns_tmp[5]), 
        .Z(KeyExpansionOutput[101]) );
  XOR2_X1 KeyExpansionIns_U5 ( .A(RoundKey[100]), .B(KeyExpansionIns_tmp[4]), 
        .Z(KeyExpansionOutput[100]) );
  XOR2_X1 KeyExpansionIns_U4 ( .A(RoundKey[0]), .B(KeyExpansionOutput[32]), 
        .Z(KeyExpansionOutput[0]) );
  XOR2_X1 KeyExpansionIns_U3 ( .A(RoundKey[32]), .B(KeyExpansionOutput[64]), 
        .Z(KeyExpansionOutput[32]) );
  XOR2_X1 KeyExpansionIns_U2 ( .A(RoundKey[64]), .B(KeyExpansionOutput[96]), 
        .Z(KeyExpansionOutput[64]) );
  XOR2_X1 KeyExpansionIns_U1 ( .A(RoundKey[96]), .B(KeyExpansionIns_tmp[0]), 
        .Z(KeyExpansionOutput[96]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U8 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_), .B(n283), .Z(
        KeyExpansionIns_tmp[31]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U7 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_), .B(n285), .Z(
        KeyExpansionIns_tmp[30]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U6 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_), .B(Rcon[5]), .Z(
        KeyExpansionIns_tmp[29]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U5 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_), .B(Rcon[4]), .Z(
        KeyExpansionIns_tmp[28]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U4 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_), .B(Rcon[3]), .Z(
        KeyExpansionIns_tmp[27]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U3 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_), .B(Rcon[2]), .Z(
        KeyExpansionIns_tmp[26]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U2 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_), .B(Rcon[1]), .Z(
        KeyExpansionIns_tmp[25]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_), .B(Rcon[0]), .Z(
        KeyExpansionIns_tmp[24]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T1_U1 ( .A(
        RoundKey[23]), .B(RoundKey[20]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T2_U1 ( .A(
        RoundKey[23]), .B(RoundKey[18]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T3_U1 ( .A(
        RoundKey[23]), .B(RoundKey[17]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T4_U1 ( .A(
        RoundKey[20]), .B(RoundKey[18]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T5_U1 ( .A(
        RoundKey[19]), .B(RoundKey[17]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T7_U1 ( .A(
        RoundKey[22]), .B(RoundKey[21]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T8_U1 ( .A(
        RoundKey[16]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T9_U1 ( .A(
        RoundKey[16]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T11_U1 ( .A(
        RoundKey[22]), .B(RoundKey[18]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T12_U1 ( .A(
        RoundKey[21]), .B(RoundKey[18]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T18_U1 ( .A(
        RoundKey[20]), .B(RoundKey[16]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T21_U1 ( .A(
        RoundKey[17]), .B(RoundKey[16]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M1_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M2_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M4_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .A2(RoundKey[16]), 
        .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M6_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M7_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M9_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M11_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M12_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M14_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M25_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M29_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M30_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M31_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M32_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M33_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M34_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M35_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M36_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M37_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M38_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M39_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M40_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M41_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M42_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M43_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M44_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M45_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M46_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M47_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M48_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .A2(RoundKey[16]), 
        .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M49_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M50_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M51_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M52_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M53_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M54_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M55_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M56_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M57_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M58_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M59_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M60_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M61_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M62_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M63_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L9_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L11_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L12_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L29_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24), .Z(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26), .ZN(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28), .ZN(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21), .Z(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22), .Z(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29), .Z(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T1_U1 ( .A(
        RoundKey[15]), .B(RoundKey[12]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T2_U1 ( .A(
        RoundKey[15]), .B(RoundKey[10]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T3_U1 ( .A(
        RoundKey[15]), .B(RoundKey[9]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T4_U1 ( .A(
        RoundKey[12]), .B(RoundKey[10]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T5_U1 ( .A(
        RoundKey[11]), .B(RoundKey[9]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T7_U1 ( .A(
        RoundKey[14]), .B(RoundKey[13]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T8_U1 ( .A(
        RoundKey[8]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T9_U1 ( .A(
        RoundKey[8]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T11_U1 ( .A(
        RoundKey[14]), .B(RoundKey[10]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T12_U1 ( .A(
        RoundKey[13]), .B(RoundKey[10]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T18_U1 ( .A(
        RoundKey[12]), .B(RoundKey[8]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T21_U1 ( .A(
        RoundKey[9]), .B(RoundKey[8]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M1_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M2_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M4_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .A2(RoundKey[8]), 
        .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M6_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M7_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M9_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M11_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M12_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M14_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M25_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M29_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M30_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M31_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M32_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M33_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M34_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M35_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M36_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M37_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M38_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M39_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M40_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M41_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M42_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M43_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M44_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M45_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M46_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M47_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M48_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .A2(RoundKey[8]), 
        .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M49_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M50_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M51_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M52_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M53_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M54_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M55_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M56_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M57_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M58_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M59_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M60_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M61_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M62_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M63_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L9_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L11_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L12_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L29_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24), .Z(
        KeyExpansionIns_tmp[23]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26), .ZN(
        KeyExpansionIns_tmp[22]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28), .ZN(
        KeyExpansionIns_tmp[21]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21), .Z(
        KeyExpansionIns_tmp[20]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22), .Z(
        KeyExpansionIns_tmp[19]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29), .Z(
        KeyExpansionIns_tmp[18]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27), .ZN(
        KeyExpansionIns_tmp[17]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23), .ZN(
        KeyExpansionIns_tmp[16]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T1_U1 ( .A(
        RoundKey[7]), .B(RoundKey[4]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T2_U1 ( .A(
        RoundKey[7]), .B(RoundKey[2]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T3_U1 ( .A(
        RoundKey[7]), .B(RoundKey[1]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T4_U1 ( .A(
        RoundKey[4]), .B(RoundKey[2]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T5_U1 ( .A(
        RoundKey[3]), .B(RoundKey[1]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T7_U1 ( .A(
        RoundKey[6]), .B(RoundKey[5]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T8_U1 ( .A(
        RoundKey[0]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T9_U1 ( .A(
        RoundKey[0]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T11_U1 ( .A(
        RoundKey[6]), .B(RoundKey[2]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T12_U1 ( .A(
        RoundKey[5]), .B(RoundKey[2]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T18_U1 ( .A(
        RoundKey[4]), .B(RoundKey[0]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T21_U1 ( .A(
        RoundKey[1]), .B(RoundKey[0]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M1_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M2_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M4_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .A2(RoundKey[0]), 
        .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M6_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M7_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M9_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M11_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M12_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M14_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M25_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M29_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M30_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M31_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M32_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M33_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M34_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M35_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M36_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M37_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M38_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M39_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M40_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M41_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M42_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M43_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M44_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M45_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M46_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M47_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M48_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .A2(RoundKey[0]), 
        .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M49_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M50_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M51_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M52_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M53_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M54_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M55_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M56_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M57_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M58_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M59_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M60_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M61_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M62_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M63_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L9_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L11_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L12_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L29_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24), .Z(
        KeyExpansionIns_tmp[15]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26), .ZN(
        KeyExpansionIns_tmp[14]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28), .ZN(
        KeyExpansionIns_tmp[13]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21), .Z(
        KeyExpansionIns_tmp[12]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22), .Z(
        KeyExpansionIns_tmp[11]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29), .Z(
        KeyExpansionIns_tmp[10]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27), .ZN(
        KeyExpansionIns_tmp[9]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23), .ZN(
        KeyExpansionIns_tmp[8]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T1_U1 ( .A(
        RoundKey[31]), .B(RoundKey[28]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T2_U1 ( .A(
        RoundKey[31]), .B(RoundKey[26]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T3_U1 ( .A(
        RoundKey[31]), .B(RoundKey[25]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T4_U1 ( .A(
        RoundKey[28]), .B(RoundKey[26]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T5_U1 ( .A(
        RoundKey[27]), .B(RoundKey[25]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T7_U1 ( .A(
        RoundKey[30]), .B(RoundKey[29]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T8_U1 ( .A(
        RoundKey[24]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T9_U1 ( .A(
        RoundKey[24]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T11_U1 ( .A(
        RoundKey[30]), .B(RoundKey[26]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T12_U1 ( .A(
        RoundKey[29]), .B(RoundKey[26]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T18_U1 ( .A(
        RoundKey[28]), .B(RoundKey[24]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T21_U1 ( .A(
        RoundKey[25]), .B(RoundKey[24]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M1_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M2_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M4_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .A2(RoundKey[24]), 
        .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M6_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M7_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M9_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M11_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M12_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M14_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M25_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M29_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M30_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M31_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M32_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M33_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M34_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M35_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M36_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M37_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M38_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M39_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M40_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M41_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M42_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M43_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M44_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M45_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M46_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M47_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M48_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .A2(RoundKey[24]), 
        .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M49_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M50_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M51_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M52_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M53_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M54_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M55_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M56_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M57_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M58_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M59_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M60_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M61_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M62_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M63_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L9_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L11_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L12_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L29_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24), .Z(
        KeyExpansionIns_tmp[7]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26), .ZN(
        KeyExpansionIns_tmp[6]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28), .ZN(
        KeyExpansionIns_tmp[5]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21), .Z(
        KeyExpansionIns_tmp[4]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22), .Z(
        KeyExpansionIns_tmp[3]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29), .Z(
        KeyExpansionIns_tmp[2]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27), .ZN(
        KeyExpansionIns_tmp[1]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23), .ZN(
        KeyExpansionIns_tmp[0]) );
  INV_X1 RoundCounterIns_U14 ( .A(RoundCounterIns_n13), .ZN(RoundCounterIns_n1) );
  MUX2_X1 RoundCounterIns_U13 ( .A(RoundCounterIns_n12), .B(
        RoundCounterIns_n11), .S(RoundCounterIns_n5), .Z(RoundCounterIns_n13)
         );
  NOR2_X1 RoundCounterIns_U12 ( .A1(reset), .A2(RoundCounterIns_n10), .ZN(
        RoundCounterIns_N8) );
  XNOR2_X1 RoundCounterIns_U11 ( .A(RoundCounter[0]), .B(RoundCounter[1]), 
        .ZN(RoundCounterIns_n10) );
  MUX2_X1 RoundCounterIns_U10 ( .A(RoundCounterIns_n9), .B(RoundCounterIns_n8), 
        .S(RoundCounter[3]), .Z(RoundCounterIns_N10) );
  NAND2_X1 RoundCounterIns_U9 ( .A1(RoundCounterIns_n12), .A2(
        RoundCounterIns_n7), .ZN(RoundCounterIns_n8) );
  NAND2_X1 RoundCounterIns_U8 ( .A1(RoundCounterIns_n5), .A2(
        RoundCounterIns_n2), .ZN(RoundCounterIns_n7) );
  NOR2_X1 RoundCounterIns_U7 ( .A1(RoundCounterIns_n4), .A2(RoundCounterIns_N7), .ZN(RoundCounterIns_n12) );
  NOR2_X1 RoundCounterIns_U6 ( .A1(RoundCounter[1]), .A2(reset), .ZN(
        RoundCounterIns_n4) );
  NOR2_X1 RoundCounterIns_U5 ( .A1(RoundCounterIns_n5), .A2(
        RoundCounterIns_n11), .ZN(RoundCounterIns_n9) );
  NAND2_X1 RoundCounterIns_U4 ( .A1(RoundCounter[1]), .A2(RoundCounterIns_n3), 
        .ZN(RoundCounterIns_n11) );
  NOR2_X1 RoundCounterIns_U3 ( .A1(reset), .A2(RoundCounterIns_n6), .ZN(
        RoundCounterIns_n3) );
  NOR2_X1 RoundCounterIns_U2 ( .A1(reset), .A2(RoundCounter[0]), .ZN(
        RoundCounterIns_N7) );
  INV_X1 RoundCounterIns_U1 ( .A(reset), .ZN(RoundCounterIns_n2) );
  INV_X1 RoundCounterIns_count_reg_0__U1 ( .A(RoundCounter[0]), .ZN(
        RoundCounterIns_n6) );
  DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .D(RoundCounterIns_N7), .CK(clk), 
        .Q(RoundCounter[0]), .QN() );
  INV_X1 RoundCounterIns_count_reg_1__U1 ( .A(RoundCounter[1]), .ZN(
        RoundCounterIns_count_reg_1__QN) );
  DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .D(RoundCounterIns_N8), .CK(clk), 
        .Q(RoundCounter[1]), .QN() );
  INV_X1 RoundCounterIns_count_reg_2__U1 ( .A(RoundCounter[2]), .ZN(
        RoundCounterIns_n5) );
  DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .D(RoundCounterIns_n1), .CK(clk), 
        .Q(RoundCounter[2]), .QN() );
  INV_X1 RoundCounterIns_count_reg_3__U1 ( .A(RoundCounter[3]), .ZN(
        RoundCounterIns_count_reg_3__QN) );
  DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .D(RoundCounterIns_N10), .CK(clk), .Q(RoundCounter[3]), .QN() );
endmodule

