/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 16 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 17 register stage(s) in total */

module sbox_HPC2_BDDcudd_Pipeline_d2 (X_s0, clk, X_s1, X_s2, Fresh, Y_s0, Y_s1, Y_s2);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [1232:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;

    /* cells in depth 0 */

    /* cells in depth 1 */
    buf_clk cell_547 ( .C (clk), .D (X_s0[5]), .Q (signal_2641) ) ;
    buf_clk cell_549 ( .C (clk), .D (X_s1[5]), .Q (signal_2643) ) ;
    buf_clk cell_551 ( .C (clk), .D (X_s2[5]), .Q (signal_2645) ) ;
    buf_clk cell_553 ( .C (clk), .D (X_s0[6]), .Q (signal_2647) ) ;
    buf_clk cell_555 ( .C (clk), .D (X_s1[6]), .Q (signal_2649) ) ;
    buf_clk cell_557 ( .C (clk), .D (X_s2[6]), .Q (signal_2651) ) ;
    buf_clk cell_589 ( .C (clk), .D (X_s0[3]), .Q (signal_2683) ) ;
    buf_clk cell_593 ( .C (clk), .D (X_s1[3]), .Q (signal_2687) ) ;
    buf_clk cell_597 ( .C (clk), .D (X_s2[3]), .Q (signal_2691) ) ;
    buf_clk cell_763 ( .C (clk), .D (X_s0[1]), .Q (signal_2857) ) ;
    buf_clk cell_771 ( .C (clk), .D (X_s1[1]), .Q (signal_2865) ) ;
    buf_clk cell_779 ( .C (clk), .D (X_s2[1]), .Q (signal_2873) ) ;
    buf_clk cell_823 ( .C (clk), .D (X_s0[2]), .Q (signal_2917) ) ;
    buf_clk cell_833 ( .C (clk), .D (X_s1[2]), .Q (signal_2927) ) ;
    buf_clk cell_843 ( .C (clk), .D (X_s2[2]), .Q (signal_2937) ) ;
    buf_clk cell_853 ( .C (clk), .D (X_s0[4]), .Q (signal_2947) ) ;
    buf_clk cell_865 ( .C (clk), .D (X_s1[4]), .Q (signal_2959) ) ;
    buf_clk cell_877 ( .C (clk), .D (X_s2[4]), .Q (signal_2971) ) ;
    buf_clk cell_889 ( .C (clk), .D (X_s0[7]), .Q (signal_2983) ) ;
    buf_clk cell_903 ( .C (clk), .D (X_s1[7]), .Q (signal_2997) ) ;
    buf_clk cell_917 ( .C (clk), .D (X_s2[7]), .Q (signal_3011) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_136 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_557, signal_556, signal_151}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_137 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({signal_561, signal_560, signal_152}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_138 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_563, signal_562, signal_153}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_139 ( .s ({X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({signal_567, signal_566, signal_154}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_140 ( .s ({X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_569, signal_568, signal_155}) ) ;
    buf_clk cell_548 ( .C (clk), .D (signal_2641), .Q (signal_2642) ) ;
    buf_clk cell_550 ( .C (clk), .D (signal_2643), .Q (signal_2644) ) ;
    buf_clk cell_552 ( .C (clk), .D (signal_2645), .Q (signal_2646) ) ;
    buf_clk cell_554 ( .C (clk), .D (signal_2647), .Q (signal_2648) ) ;
    buf_clk cell_556 ( .C (clk), .D (signal_2649), .Q (signal_2650) ) ;
    buf_clk cell_558 ( .C (clk), .D (signal_2651), .Q (signal_2652) ) ;
    buf_clk cell_590 ( .C (clk), .D (signal_2683), .Q (signal_2684) ) ;
    buf_clk cell_594 ( .C (clk), .D (signal_2687), .Q (signal_2688) ) ;
    buf_clk cell_598 ( .C (clk), .D (signal_2691), .Q (signal_2692) ) ;
    buf_clk cell_764 ( .C (clk), .D (signal_2857), .Q (signal_2858) ) ;
    buf_clk cell_772 ( .C (clk), .D (signal_2865), .Q (signal_2866) ) ;
    buf_clk cell_780 ( .C (clk), .D (signal_2873), .Q (signal_2874) ) ;
    buf_clk cell_824 ( .C (clk), .D (signal_2917), .Q (signal_2918) ) ;
    buf_clk cell_834 ( .C (clk), .D (signal_2927), .Q (signal_2928) ) ;
    buf_clk cell_844 ( .C (clk), .D (signal_2937), .Q (signal_2938) ) ;
    buf_clk cell_854 ( .C (clk), .D (signal_2947), .Q (signal_2948) ) ;
    buf_clk cell_866 ( .C (clk), .D (signal_2959), .Q (signal_2960) ) ;
    buf_clk cell_878 ( .C (clk), .D (signal_2971), .Q (signal_2972) ) ;
    buf_clk cell_890 ( .C (clk), .D (signal_2983), .Q (signal_2984) ) ;
    buf_clk cell_904 ( .C (clk), .D (signal_2997), .Q (signal_2998) ) ;
    buf_clk cell_918 ( .C (clk), .D (signal_3011), .Q (signal_3012) ) ;

    /* cells in depth 3 */
    buf_clk cell_559 ( .C (clk), .D (signal_2648), .Q (signal_2653) ) ;
    buf_clk cell_561 ( .C (clk), .D (signal_2650), .Q (signal_2655) ) ;
    buf_clk cell_563 ( .C (clk), .D (signal_2652), .Q (signal_2657) ) ;
    buf_clk cell_565 ( .C (clk), .D (signal_153), .Q (signal_2659) ) ;
    buf_clk cell_567 ( .C (clk), .D (signal_562), .Q (signal_2661) ) ;
    buf_clk cell_569 ( .C (clk), .D (signal_563), .Q (signal_2663) ) ;
    buf_clk cell_571 ( .C (clk), .D (signal_154), .Q (signal_2665) ) ;
    buf_clk cell_573 ( .C (clk), .D (signal_566), .Q (signal_2667) ) ;
    buf_clk cell_575 ( .C (clk), .D (signal_567), .Q (signal_2669) ) ;
    buf_clk cell_577 ( .C (clk), .D (signal_151), .Q (signal_2671) ) ;
    buf_clk cell_579 ( .C (clk), .D (signal_556), .Q (signal_2673) ) ;
    buf_clk cell_581 ( .C (clk), .D (signal_557), .Q (signal_2675) ) ;
    buf_clk cell_583 ( .C (clk), .D (signal_155), .Q (signal_2677) ) ;
    buf_clk cell_585 ( .C (clk), .D (signal_568), .Q (signal_2679) ) ;
    buf_clk cell_587 ( .C (clk), .D (signal_569), .Q (signal_2681) ) ;
    buf_clk cell_591 ( .C (clk), .D (signal_2684), .Q (signal_2685) ) ;
    buf_clk cell_595 ( .C (clk), .D (signal_2688), .Q (signal_2689) ) ;
    buf_clk cell_599 ( .C (clk), .D (signal_2692), .Q (signal_2693) ) ;
    buf_clk cell_601 ( .C (clk), .D (signal_152), .Q (signal_2695) ) ;
    buf_clk cell_603 ( .C (clk), .D (signal_560), .Q (signal_2697) ) ;
    buf_clk cell_605 ( .C (clk), .D (signal_561), .Q (signal_2699) ) ;
    buf_clk cell_765 ( .C (clk), .D (signal_2858), .Q (signal_2859) ) ;
    buf_clk cell_773 ( .C (clk), .D (signal_2866), .Q (signal_2867) ) ;
    buf_clk cell_781 ( .C (clk), .D (signal_2874), .Q (signal_2875) ) ;
    buf_clk cell_825 ( .C (clk), .D (signal_2918), .Q (signal_2919) ) ;
    buf_clk cell_835 ( .C (clk), .D (signal_2928), .Q (signal_2929) ) ;
    buf_clk cell_845 ( .C (clk), .D (signal_2938), .Q (signal_2939) ) ;
    buf_clk cell_855 ( .C (clk), .D (signal_2948), .Q (signal_2949) ) ;
    buf_clk cell_867 ( .C (clk), .D (signal_2960), .Q (signal_2961) ) ;
    buf_clk cell_879 ( .C (clk), .D (signal_2972), .Q (signal_2973) ) ;
    buf_clk cell_891 ( .C (clk), .D (signal_2984), .Q (signal_2985) ) ;
    buf_clk cell_905 ( .C (clk), .D (signal_2998), .Q (signal_2999) ) ;
    buf_clk cell_919 ( .C (clk), .D (signal_3012), .Q (signal_3013) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_141 ( .s ({signal_2646, signal_2644, signal_2642}), .b ({signal_569, signal_568, signal_155}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({signal_571, signal_570, signal_156}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_142 ( .s ({signal_2646, signal_2644, signal_2642}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_569, signal_568, signal_155}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_573, signal_572, signal_157}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_143 ( .s ({signal_2646, signal_2644, signal_2642}), .b ({signal_567, signal_566, signal_154}), .a ({signal_569, signal_568, signal_155}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({signal_575, signal_574, signal_158}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_144 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_563, signal_562, signal_153}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_577, signal_576, signal_159}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_145 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_569, signal_568, signal_155}), .a ({signal_567, signal_566, signal_154}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({signal_579, signal_578, signal_160}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_146 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_563, signal_562, signal_153}), .a ({signal_567, signal_566, signal_154}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_581, signal_580, signal_161}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_147 ( .s ({signal_2646, signal_2644, signal_2642}), .b ({signal_569, signal_568, signal_155}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({signal_583, signal_582, signal_162}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_148 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_557, signal_556, signal_151}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_585, signal_584, signal_163}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_149 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_563, signal_562, signal_153}), .a ({signal_569, signal_568, signal_155}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({signal_587, signal_586, signal_164}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_150 ( .s ({signal_2646, signal_2644, signal_2642}), .b ({signal_567, signal_566, signal_154}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_589, signal_588, signal_165}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_151 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_557, signal_556, signal_151}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({signal_591, signal_590, signal_166}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_152 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_567, signal_566, signal_154}), .a ({signal_557, signal_556, signal_151}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_593, signal_592, signal_167}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_153 ( .s ({signal_2646, signal_2644, signal_2642}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_567, signal_566, signal_154}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({signal_595, signal_594, signal_168}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_154 ( .s ({signal_2646, signal_2644, signal_2642}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_567, signal_566, signal_154}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_597, signal_596, signal_169}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_155 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_567, signal_566, signal_154}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({signal_599, signal_598, signal_170}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_156 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_557, signal_556, signal_151}), .a ({signal_567, signal_566, signal_154}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_601, signal_600, signal_171}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_157 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_567, signal_566, signal_154}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({signal_603, signal_602, signal_172}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_158 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_563, signal_562, signal_153}), .a ({signal_557, signal_556, signal_151}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_605, signal_604, signal_173}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_159 ( .s ({signal_2646, signal_2644, signal_2642}), .b ({signal_567, signal_566, signal_154}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({signal_607, signal_606, signal_174}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_160 ( .s ({signal_2646, signal_2644, signal_2642}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_569, signal_568, signal_155}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_609, signal_608, signal_175}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_161 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_563, signal_562, signal_153}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({signal_611, signal_610, signal_176}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_162 ( .s ({signal_2646, signal_2644, signal_2642}), .b ({signal_569, signal_568, signal_155}), .a ({signal_567, signal_566, signal_154}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_613, signal_612, signal_177}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_163 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_557, signal_556, signal_151}), .a ({signal_563, signal_562, signal_153}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({signal_615, signal_614, signal_178}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_164 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_567, signal_566, signal_154}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_617, signal_616, signal_179}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_165 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_569, signal_568, signal_155}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({signal_619, signal_618, signal_180}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_166 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_569, signal_568, signal_155}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_621, signal_620, signal_181}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_167 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_569, signal_568, signal_155}), .a ({signal_557, signal_556, signal_151}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({signal_623, signal_622, signal_182}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_168 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({signal_563, signal_562, signal_153}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_625, signal_624, signal_183}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_169 ( .s ({signal_2652, signal_2650, signal_2648}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_557, signal_556, signal_151}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({signal_627, signal_626, signal_184}) ) ;
    buf_clk cell_560 ( .C (clk), .D (signal_2653), .Q (signal_2654) ) ;
    buf_clk cell_562 ( .C (clk), .D (signal_2655), .Q (signal_2656) ) ;
    buf_clk cell_564 ( .C (clk), .D (signal_2657), .Q (signal_2658) ) ;
    buf_clk cell_566 ( .C (clk), .D (signal_2659), .Q (signal_2660) ) ;
    buf_clk cell_568 ( .C (clk), .D (signal_2661), .Q (signal_2662) ) ;
    buf_clk cell_570 ( .C (clk), .D (signal_2663), .Q (signal_2664) ) ;
    buf_clk cell_572 ( .C (clk), .D (signal_2665), .Q (signal_2666) ) ;
    buf_clk cell_574 ( .C (clk), .D (signal_2667), .Q (signal_2668) ) ;
    buf_clk cell_576 ( .C (clk), .D (signal_2669), .Q (signal_2670) ) ;
    buf_clk cell_578 ( .C (clk), .D (signal_2671), .Q (signal_2672) ) ;
    buf_clk cell_580 ( .C (clk), .D (signal_2673), .Q (signal_2674) ) ;
    buf_clk cell_582 ( .C (clk), .D (signal_2675), .Q (signal_2676) ) ;
    buf_clk cell_584 ( .C (clk), .D (signal_2677), .Q (signal_2678) ) ;
    buf_clk cell_586 ( .C (clk), .D (signal_2679), .Q (signal_2680) ) ;
    buf_clk cell_588 ( .C (clk), .D (signal_2681), .Q (signal_2682) ) ;
    buf_clk cell_592 ( .C (clk), .D (signal_2685), .Q (signal_2686) ) ;
    buf_clk cell_596 ( .C (clk), .D (signal_2689), .Q (signal_2690) ) ;
    buf_clk cell_600 ( .C (clk), .D (signal_2693), .Q (signal_2694) ) ;
    buf_clk cell_602 ( .C (clk), .D (signal_2695), .Q (signal_2696) ) ;
    buf_clk cell_604 ( .C (clk), .D (signal_2697), .Q (signal_2698) ) ;
    buf_clk cell_606 ( .C (clk), .D (signal_2699), .Q (signal_2700) ) ;
    buf_clk cell_766 ( .C (clk), .D (signal_2859), .Q (signal_2860) ) ;
    buf_clk cell_774 ( .C (clk), .D (signal_2867), .Q (signal_2868) ) ;
    buf_clk cell_782 ( .C (clk), .D (signal_2875), .Q (signal_2876) ) ;
    buf_clk cell_826 ( .C (clk), .D (signal_2919), .Q (signal_2920) ) ;
    buf_clk cell_836 ( .C (clk), .D (signal_2929), .Q (signal_2930) ) ;
    buf_clk cell_846 ( .C (clk), .D (signal_2939), .Q (signal_2940) ) ;
    buf_clk cell_856 ( .C (clk), .D (signal_2949), .Q (signal_2950) ) ;
    buf_clk cell_868 ( .C (clk), .D (signal_2961), .Q (signal_2962) ) ;
    buf_clk cell_880 ( .C (clk), .D (signal_2973), .Q (signal_2974) ) ;
    buf_clk cell_892 ( .C (clk), .D (signal_2985), .Q (signal_2986) ) ;
    buf_clk cell_906 ( .C (clk), .D (signal_2999), .Q (signal_3000) ) ;
    buf_clk cell_920 ( .C (clk), .D (signal_3013), .Q (signal_3014) ) ;

    /* cells in depth 5 */
    buf_clk cell_607 ( .C (clk), .D (signal_2686), .Q (signal_2701) ) ;
    buf_clk cell_609 ( .C (clk), .D (signal_2690), .Q (signal_2703) ) ;
    buf_clk cell_611 ( .C (clk), .D (signal_2694), .Q (signal_2705) ) ;
    buf_clk cell_613 ( .C (clk), .D (signal_2672), .Q (signal_2707) ) ;
    buf_clk cell_615 ( .C (clk), .D (signal_2674), .Q (signal_2709) ) ;
    buf_clk cell_617 ( .C (clk), .D (signal_2676), .Q (signal_2711) ) ;
    buf_clk cell_619 ( .C (clk), .D (signal_2696), .Q (signal_2713) ) ;
    buf_clk cell_621 ( .C (clk), .D (signal_2698), .Q (signal_2715) ) ;
    buf_clk cell_623 ( .C (clk), .D (signal_2700), .Q (signal_2717) ) ;
    buf_clk cell_625 ( .C (clk), .D (signal_182), .Q (signal_2719) ) ;
    buf_clk cell_627 ( .C (clk), .D (signal_622), .Q (signal_2721) ) ;
    buf_clk cell_629 ( .C (clk), .D (signal_623), .Q (signal_2723) ) ;
    buf_clk cell_631 ( .C (clk), .D (signal_175), .Q (signal_2725) ) ;
    buf_clk cell_633 ( .C (clk), .D (signal_608), .Q (signal_2727) ) ;
    buf_clk cell_635 ( .C (clk), .D (signal_609), .Q (signal_2729) ) ;
    buf_clk cell_637 ( .C (clk), .D (signal_177), .Q (signal_2731) ) ;
    buf_clk cell_639 ( .C (clk), .D (signal_612), .Q (signal_2733) ) ;
    buf_clk cell_641 ( .C (clk), .D (signal_613), .Q (signal_2735) ) ;
    buf_clk cell_643 ( .C (clk), .D (signal_169), .Q (signal_2737) ) ;
    buf_clk cell_645 ( .C (clk), .D (signal_596), .Q (signal_2739) ) ;
    buf_clk cell_647 ( .C (clk), .D (signal_597), .Q (signal_2741) ) ;
    buf_clk cell_649 ( .C (clk), .D (signal_178), .Q (signal_2743) ) ;
    buf_clk cell_651 ( .C (clk), .D (signal_614), .Q (signal_2745) ) ;
    buf_clk cell_653 ( .C (clk), .D (signal_615), .Q (signal_2747) ) ;
    buf_clk cell_655 ( .C (clk), .D (signal_167), .Q (signal_2749) ) ;
    buf_clk cell_657 ( .C (clk), .D (signal_592), .Q (signal_2751) ) ;
    buf_clk cell_659 ( .C (clk), .D (signal_593), .Q (signal_2753) ) ;
    buf_clk cell_661 ( .C (clk), .D (signal_171), .Q (signal_2755) ) ;
    buf_clk cell_663 ( .C (clk), .D (signal_600), .Q (signal_2757) ) ;
    buf_clk cell_665 ( .C (clk), .D (signal_601), .Q (signal_2759) ) ;
    buf_clk cell_667 ( .C (clk), .D (signal_183), .Q (signal_2761) ) ;
    buf_clk cell_669 ( .C (clk), .D (signal_624), .Q (signal_2763) ) ;
    buf_clk cell_671 ( .C (clk), .D (signal_625), .Q (signal_2765) ) ;
    buf_clk cell_673 ( .C (clk), .D (signal_184), .Q (signal_2767) ) ;
    buf_clk cell_675 ( .C (clk), .D (signal_626), .Q (signal_2769) ) ;
    buf_clk cell_677 ( .C (clk), .D (signal_627), .Q (signal_2771) ) ;
    buf_clk cell_679 ( .C (clk), .D (signal_180), .Q (signal_2773) ) ;
    buf_clk cell_681 ( .C (clk), .D (signal_618), .Q (signal_2775) ) ;
    buf_clk cell_683 ( .C (clk), .D (signal_619), .Q (signal_2777) ) ;
    buf_clk cell_685 ( .C (clk), .D (signal_172), .Q (signal_2779) ) ;
    buf_clk cell_687 ( .C (clk), .D (signal_602), .Q (signal_2781) ) ;
    buf_clk cell_689 ( .C (clk), .D (signal_603), .Q (signal_2783) ) ;
    buf_clk cell_691 ( .C (clk), .D (signal_163), .Q (signal_2785) ) ;
    buf_clk cell_693 ( .C (clk), .D (signal_584), .Q (signal_2787) ) ;
    buf_clk cell_695 ( .C (clk), .D (signal_585), .Q (signal_2789) ) ;
    buf_clk cell_697 ( .C (clk), .D (signal_168), .Q (signal_2791) ) ;
    buf_clk cell_699 ( .C (clk), .D (signal_594), .Q (signal_2793) ) ;
    buf_clk cell_701 ( .C (clk), .D (signal_595), .Q (signal_2795) ) ;
    buf_clk cell_703 ( .C (clk), .D (signal_170), .Q (signal_2797) ) ;
    buf_clk cell_705 ( .C (clk), .D (signal_598), .Q (signal_2799) ) ;
    buf_clk cell_707 ( .C (clk), .D (signal_599), .Q (signal_2801) ) ;
    buf_clk cell_709 ( .C (clk), .D (signal_161), .Q (signal_2803) ) ;
    buf_clk cell_711 ( .C (clk), .D (signal_580), .Q (signal_2805) ) ;
    buf_clk cell_713 ( .C (clk), .D (signal_581), .Q (signal_2807) ) ;
    buf_clk cell_715 ( .C (clk), .D (signal_164), .Q (signal_2809) ) ;
    buf_clk cell_717 ( .C (clk), .D (signal_586), .Q (signal_2811) ) ;
    buf_clk cell_719 ( .C (clk), .D (signal_587), .Q (signal_2813) ) ;
    buf_clk cell_721 ( .C (clk), .D (signal_162), .Q (signal_2815) ) ;
    buf_clk cell_723 ( .C (clk), .D (signal_582), .Q (signal_2817) ) ;
    buf_clk cell_725 ( .C (clk), .D (signal_583), .Q (signal_2819) ) ;
    buf_clk cell_727 ( .C (clk), .D (signal_173), .Q (signal_2821) ) ;
    buf_clk cell_729 ( .C (clk), .D (signal_604), .Q (signal_2823) ) ;
    buf_clk cell_731 ( .C (clk), .D (signal_605), .Q (signal_2825) ) ;
    buf_clk cell_733 ( .C (clk), .D (signal_158), .Q (signal_2827) ) ;
    buf_clk cell_735 ( .C (clk), .D (signal_574), .Q (signal_2829) ) ;
    buf_clk cell_737 ( .C (clk), .D (signal_575), .Q (signal_2831) ) ;
    buf_clk cell_739 ( .C (clk), .D (signal_181), .Q (signal_2833) ) ;
    buf_clk cell_741 ( .C (clk), .D (signal_620), .Q (signal_2835) ) ;
    buf_clk cell_743 ( .C (clk), .D (signal_621), .Q (signal_2837) ) ;
    buf_clk cell_745 ( .C (clk), .D (signal_176), .Q (signal_2839) ) ;
    buf_clk cell_747 ( .C (clk), .D (signal_610), .Q (signal_2841) ) ;
    buf_clk cell_749 ( .C (clk), .D (signal_611), .Q (signal_2843) ) ;
    buf_clk cell_751 ( .C (clk), .D (signal_157), .Q (signal_2845) ) ;
    buf_clk cell_753 ( .C (clk), .D (signal_572), .Q (signal_2847) ) ;
    buf_clk cell_755 ( .C (clk), .D (signal_573), .Q (signal_2849) ) ;
    buf_clk cell_757 ( .C (clk), .D (signal_166), .Q (signal_2851) ) ;
    buf_clk cell_759 ( .C (clk), .D (signal_590), .Q (signal_2853) ) ;
    buf_clk cell_761 ( .C (clk), .D (signal_591), .Q (signal_2855) ) ;
    buf_clk cell_767 ( .C (clk), .D (signal_2860), .Q (signal_2861) ) ;
    buf_clk cell_775 ( .C (clk), .D (signal_2868), .Q (signal_2869) ) ;
    buf_clk cell_783 ( .C (clk), .D (signal_2876), .Q (signal_2877) ) ;
    buf_clk cell_827 ( .C (clk), .D (signal_2920), .Q (signal_2921) ) ;
    buf_clk cell_837 ( .C (clk), .D (signal_2930), .Q (signal_2931) ) ;
    buf_clk cell_847 ( .C (clk), .D (signal_2940), .Q (signal_2941) ) ;
    buf_clk cell_857 ( .C (clk), .D (signal_2950), .Q (signal_2951) ) ;
    buf_clk cell_869 ( .C (clk), .D (signal_2962), .Q (signal_2963) ) ;
    buf_clk cell_881 ( .C (clk), .D (signal_2974), .Q (signal_2975) ) ;
    buf_clk cell_893 ( .C (clk), .D (signal_2986), .Q (signal_2987) ) ;
    buf_clk cell_907 ( .C (clk), .D (signal_3000), .Q (signal_3001) ) ;
    buf_clk cell_921 ( .C (clk), .D (signal_3014), .Q (signal_3015) ) ;

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_170 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_571, signal_570, signal_156}), .a ({signal_2664, signal_2662, signal_2660}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_629, signal_628, signal_185}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_171 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_609, signal_608, signal_175}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({signal_631, signal_630, signal_186}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_172 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_595, signal_594, signal_168}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_633, signal_632, signal_187}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_173 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({signal_635, signal_634, signal_188}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_174 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_595, signal_594, signal_168}), .a ({signal_597, signal_596, signal_169}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_637, signal_636, signal_189}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_175 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2670, signal_2668, signal_2666}), .a ({signal_613, signal_612, signal_177}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({signal_639, signal_638, signal_190}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_176 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2664, signal_2662, signal_2660}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_641, signal_640, signal_191}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_177 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2664, signal_2662, signal_2660}), .a ({signal_607, signal_606, signal_174}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({signal_643, signal_642, signal_192}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_178 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2676, signal_2674, signal_2672}), .a ({signal_609, signal_608, signal_175}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_645, signal_644, signal_193}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_179 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({signal_647, signal_646, signal_194}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_180 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_2682, signal_2680, signal_2678}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_649, signal_648, signal_195}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_181 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({signal_651, signal_650, signal_196}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_182 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_573, signal_572, signal_157}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_653, signal_652, signal_197}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_183 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_609, signal_608, signal_175}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({signal_655, signal_654, signal_198}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_184 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_571, signal_570, signal_156}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_657, signal_656, signal_199}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_185 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_595, signal_594, signal_168}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({signal_659, signal_658, signal_200}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_186 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2670, signal_2668, signal_2666}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_661, signal_660, signal_201}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_187 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_573, signal_572, signal_157}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({signal_663, signal_662, signal_202}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_188 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_583, signal_582, signal_162}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_665, signal_664, signal_203}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_189 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_571, signal_570, signal_156}), .a ({signal_2682, signal_2680, signal_2678}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({signal_667, signal_666, signal_204}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_190 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2670, signal_2668, signal_2666}), .a ({signal_597, signal_596, signal_169}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_669, signal_668, signal_205}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_191 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_583, signal_582, signal_162}), .a ({signal_2676, signal_2674, signal_2672}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({signal_671, signal_670, signal_206}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_192 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_609, signal_608, signal_175}), .a ({signal_2676, signal_2674, signal_2672}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_673, signal_672, signal_207}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_193 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_597, signal_596, signal_169}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({signal_675, signal_674, signal_208}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_194 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_583, signal_582, signal_162}), .a ({signal_613, signal_612, signal_177}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_677, signal_676, signal_209}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_195 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_573, signal_572, signal_157}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({signal_679, signal_678, signal_210}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_196 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_681, signal_680, signal_211}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_197 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2682, signal_2680, signal_2678}), .a ({signal_607, signal_606, signal_174}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({signal_683, signal_682, signal_212}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_198 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_575, signal_574, signal_158}), .a ({signal_2664, signal_2662, signal_2660}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_685, signal_684, signal_213}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_199 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_575, signal_574, signal_158}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({signal_687, signal_686, signal_214}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_200 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_595, signal_594, signal_168}), .a ({signal_613, signal_612, signal_177}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_689, signal_688, signal_215}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_201 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_609, signal_608, signal_175}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({signal_691, signal_690, signal_216}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_202 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_589, signal_588, signal_165}), .a ({signal_609, signal_608, signal_175}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_693, signal_692, signal_217}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_203 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_2664, signal_2662, signal_2660}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({signal_695, signal_694, signal_218}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_204 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2682, signal_2680, signal_2678}), .a ({signal_597, signal_596, signal_169}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({signal_697, signal_696, signal_219}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_205 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2682, signal_2680, signal_2678}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({signal_699, signal_698, signal_220}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_206 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_595, signal_594, signal_168}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_701, signal_700, signal_221}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_207 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_571, signal_570, signal_156}), .a ({signal_607, signal_606, signal_174}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({signal_703, signal_702, signal_222}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_208 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_575, signal_574, signal_158}), .a ({signal_2682, signal_2680, signal_2678}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({signal_705, signal_704, signal_223}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_209 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_613, signal_612, signal_177}), .a ({signal_2670, signal_2668, signal_2666}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({signal_707, signal_706, signal_224}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_210 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_571, signal_570, signal_156}), .a ({signal_583, signal_582, signal_162}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({signal_709, signal_708, signal_225}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_211 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_571, signal_570, signal_156}), .a ({signal_609, signal_608, signal_175}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({signal_711, signal_710, signal_226}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_212 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_575, signal_574, signal_158}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({signal_713, signal_712, signal_227}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_213 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2664, signal_2662, signal_2660}), .a ({signal_613, signal_612, signal_177}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({signal_715, signal_714, signal_228}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_214 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_573, signal_572, signal_157}), .a ({signal_613, signal_612, signal_177}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({signal_717, signal_716, signal_229}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_215 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({signal_719, signal_718, signal_230}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_216 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_571, signal_570, signal_156}), .a ({signal_2670, signal_2668, signal_2666}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_721, signal_720, signal_231}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_217 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_2670, signal_2668, signal_2666}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({signal_723, signal_722, signal_232}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_218 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({signal_725, signal_724, signal_233}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_219 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_607, signal_606, signal_174}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({signal_727, signal_726, signal_234}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_220 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2676, signal_2674, signal_2672}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({signal_729, signal_728, signal_235}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_221 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_573, signal_572, signal_157}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({signal_731, signal_730, signal_236}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_222 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_613, signal_612, signal_177}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({signal_733, signal_732, signal_237}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_223 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_583, signal_582, signal_162}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({signal_735, signal_734, signal_238}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_224 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_583, signal_582, signal_162}), .a ({signal_571, signal_570, signal_156}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({signal_737, signal_736, signal_239}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_225 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2682, signal_2680, signal_2678}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({signal_739, signal_738, signal_240}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_226 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_571, signal_570, signal_156}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_741, signal_740, signal_241}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_227 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_589, signal_588, signal_165}), .a ({signal_2670, signal_2668, signal_2666}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({signal_743, signal_742, signal_242}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_228 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_2676, signal_2674, signal_2672}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({signal_745, signal_744, signal_243}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_229 ( .s ({signal_2694, signal_2690, signal_2686}), .b ({signal_579, signal_578, signal_160}), .a ({signal_611, signal_610, signal_176}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({signal_749, signal_748, signal_244}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_230 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_583, signal_582, signal_162}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({signal_751, signal_750, signal_245}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_231 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_595, signal_594, signal_168}), .a ({signal_607, signal_606, signal_174}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({signal_753, signal_752, signal_246}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_232 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_613, signal_612, signal_177}), .a ({signal_573, signal_572, signal_157}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({signal_755, signal_754, signal_247}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_233 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({signal_757, signal_756, signal_248}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_234 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_609, signal_608, signal_175}), .a ({signal_597, signal_596, signal_169}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({signal_759, signal_758, signal_249}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_235 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_583, signal_582, signal_162}), .a ({signal_573, signal_572, signal_157}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({signal_761, signal_760, signal_250}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_236 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_609, signal_608, signal_175}), .a ({signal_571, signal_570, signal_156}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_763, signal_762, signal_251}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_237 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({signal_765, signal_764, signal_252}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_238 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_613, signal_612, signal_177}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({signal_767, signal_766, signal_253}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_239 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_573, signal_572, signal_157}), .a ({signal_2670, signal_2668, signal_2666}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({signal_769, signal_768, signal_254}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_240 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_595, signal_594, signal_168}), .a ({signal_609, signal_608, signal_175}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({signal_771, signal_770, signal_255}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_241 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2670, signal_2668, signal_2666}), .a ({signal_573, signal_572, signal_157}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({signal_773, signal_772, signal_256}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_242 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2682, signal_2680, signal_2678}), .a ({signal_571, signal_570, signal_156}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({signal_775, signal_774, signal_257}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_243 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_613, signal_612, signal_177}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({signal_777, signal_776, signal_258}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_244 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_571, signal_570, signal_156}), .a ({signal_597, signal_596, signal_169}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({signal_779, signal_778, signal_259}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_245 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_609, signal_608, signal_175}), .a ({signal_2682, signal_2680, signal_2678}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({signal_781, signal_780, signal_260}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_246 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_2670, signal_2668, signal_2666}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_783, signal_782, signal_261}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_247 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2676, signal_2674, signal_2672}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({signal_785, signal_784, signal_262}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_248 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_589, signal_588, signal_165}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({signal_787, signal_786, signal_263}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_249 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_573, signal_572, signal_157}), .a ({signal_2676, signal_2674, signal_2672}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({signal_789, signal_788, signal_264}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_250 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_583, signal_582, signal_162}), .a ({signal_2664, signal_2662, signal_2660}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({signal_791, signal_790, signal_265}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_251 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2664, signal_2662, signal_2660}), .a ({signal_571, signal_570, signal_156}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({signal_793, signal_792, signal_266}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_252 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2682, signal_2680, signal_2678}), .a ({signal_613, signal_612, signal_177}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({signal_795, signal_794, signal_267}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_253 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2676, signal_2674, signal_2672}), .a ({signal_583, signal_582, signal_162}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({signal_797, signal_796, signal_268}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_254 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2676, signal_2674, signal_2672}), .a ({signal_597, signal_596, signal_169}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({signal_799, signal_798, signal_269}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_255 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_589, signal_588, signal_165}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({signal_801, signal_800, signal_270}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_256 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_575, signal_574, signal_158}), .a ({signal_571, signal_570, signal_156}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_803, signal_802, signal_271}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_257 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_595, signal_594, signal_168}), .a ({signal_2670, signal_2668, signal_2666}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({signal_805, signal_804, signal_272}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_258 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({signal_807, signal_806, signal_273}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_259 ( .s ({signal_2694, signal_2690, signal_2686}), .b ({signal_2682, signal_2680, signal_2678}), .a ({signal_587, signal_586, signal_164}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({signal_809, signal_808, signal_274}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_260 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_573, signal_572, signal_157}), .a ({signal_2664, signal_2662, signal_2660}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({signal_811, signal_810, signal_275}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_261 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_2664, signal_2662, signal_2660}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({signal_813, signal_812, signal_276}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_262 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_609, signal_608, signal_175}), .a ({signal_583, signal_582, signal_162}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({signal_815, signal_814, signal_277}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_263 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_613, signal_612, signal_177}), .a ({signal_583, signal_582, signal_162}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({signal_817, signal_816, signal_278}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_264 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({signal_819, signal_818, signal_279}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_265 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_613, signal_612, signal_177}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({signal_821, signal_820, signal_280}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_266 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_609, signal_608, signal_175}), .a ({signal_607, signal_606, signal_174}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_823, signal_822, signal_281}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_267 ( .s ({signal_2694, signal_2690, signal_2686}), .b ({signal_571, signal_570, signal_156}), .a ({signal_2700, signal_2698, signal_2696}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({signal_825, signal_824, signal_282}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_268 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_573, signal_572, signal_157}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({signal_827, signal_826, signal_283}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_269 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_583, signal_582, signal_162}), .a ({signal_609, signal_608, signal_175}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({signal_829, signal_828, signal_284}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_270 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({signal_831, signal_830, signal_285}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_271 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_571, signal_570, signal_156}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({signal_833, signal_832, signal_286}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_272 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_571, signal_570, signal_156}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({signal_835, signal_834, signal_287}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_273 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2670, signal_2668, signal_2666}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({signal_837, signal_836, signal_288}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_274 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_583, signal_582, signal_162}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({signal_839, signal_838, signal_289}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_275 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_613, signal_612, signal_177}), .a ({signal_607, signal_606, signal_174}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({signal_841, signal_840, signal_290}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_276 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_571, signal_570, signal_156}), .a ({signal_613, signal_612, signal_177}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_843, signal_842, signal_291}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_277 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_589, signal_588, signal_165}), .a ({signal_2676, signal_2674, signal_2672}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({signal_845, signal_844, signal_292}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_278 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_609, signal_608, signal_175}), .a ({signal_573, signal_572, signal_157}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({signal_847, signal_846, signal_293}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_279 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({signal_849, signal_848, signal_294}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_280 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_583, signal_582, signal_162}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({signal_851, signal_850, signal_295}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_281 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_597, signal_596, signal_169}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({signal_853, signal_852, signal_296}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_282 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({signal_855, signal_854, signal_297}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_283 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({signal_857, signal_856, signal_298}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_284 ( .s ({signal_2694, signal_2690, signal_2686}), .b ({signal_623, signal_622, signal_182}), .a ({signal_2664, signal_2662, signal_2660}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({signal_859, signal_858, signal_299}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_285 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_613, signal_612, signal_177}), .a ({signal_609, signal_608, signal_175}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({signal_861, signal_860, signal_300}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_286 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_575, signal_574, signal_158}), .a ({signal_583, signal_582, signal_162}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_863, signal_862, signal_301}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_287 ( .s ({signal_2694, signal_2690, signal_2686}), .b ({signal_577, signal_576, signal_159}), .a ({signal_581, signal_580, signal_161}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({signal_865, signal_864, signal_302}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_288 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_613, signal_612, signal_177}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({signal_867, signal_866, signal_303}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_289 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2664, signal_2662, signal_2660}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({signal_869, signal_868, signal_304}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_290 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_597, signal_596, signal_169}), .a ({signal_2682, signal_2680, signal_2678}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({signal_871, signal_870, signal_305}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_291 ( .s ({signal_2694, signal_2690, signal_2686}), .b ({signal_617, signal_616, signal_179}), .a ({signal_571, signal_570, signal_156}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({signal_873, signal_872, signal_306}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_292 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2682, signal_2680, signal_2678}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({signal_875, signal_874, signal_307}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_293 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_595, signal_594, signal_168}), .a ({signal_589, signal_588, signal_165}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({signal_877, signal_876, signal_308}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_294 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2676, signal_2674, signal_2672}), .a ({signal_613, signal_612, signal_177}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({signal_879, signal_878, signal_309}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_295 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_595, signal_594, signal_168}), .a ({signal_583, signal_582, signal_162}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({signal_881, signal_880, signal_310}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_296 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2664, signal_2662, signal_2660}), .a ({signal_597, signal_596, signal_169}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_883, signal_882, signal_311}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_297 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_583, signal_582, signal_162}), .a ({signal_607, signal_606, signal_174}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({signal_885, signal_884, signal_312}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_298 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_575, signal_574, signal_158}), .a ({signal_607, signal_606, signal_174}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({signal_887, signal_886, signal_313}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_299 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2670, signal_2668, signal_2666}), .a ({signal_571, signal_570, signal_156}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({signal_889, signal_888, signal_314}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_300 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_2676, signal_2674, signal_2672}), .a ({signal_575, signal_574, signal_158}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({signal_891, signal_890, signal_315}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_301 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_607, signal_606, signal_174}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({signal_893, signal_892, signal_316}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_302 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_607, signal_606, signal_174}), .a ({signal_595, signal_594, signal_168}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({signal_895, signal_894, signal_317}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_303 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_589, signal_588, signal_165}), .a ({signal_597, signal_596, signal_169}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({signal_897, signal_896, signal_318}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_304 ( .s ({signal_2658, signal_2656, signal_2654}), .b ({signal_609, signal_608, signal_175}), .a ({signal_2664, signal_2662, signal_2660}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({signal_899, signal_898, signal_319}) ) ;
    buf_clk cell_608 ( .C (clk), .D (signal_2701), .Q (signal_2702) ) ;
    buf_clk cell_610 ( .C (clk), .D (signal_2703), .Q (signal_2704) ) ;
    buf_clk cell_612 ( .C (clk), .D (signal_2705), .Q (signal_2706) ) ;
    buf_clk cell_614 ( .C (clk), .D (signal_2707), .Q (signal_2708) ) ;
    buf_clk cell_616 ( .C (clk), .D (signal_2709), .Q (signal_2710) ) ;
    buf_clk cell_618 ( .C (clk), .D (signal_2711), .Q (signal_2712) ) ;
    buf_clk cell_620 ( .C (clk), .D (signal_2713), .Q (signal_2714) ) ;
    buf_clk cell_622 ( .C (clk), .D (signal_2715), .Q (signal_2716) ) ;
    buf_clk cell_624 ( .C (clk), .D (signal_2717), .Q (signal_2718) ) ;
    buf_clk cell_626 ( .C (clk), .D (signal_2719), .Q (signal_2720) ) ;
    buf_clk cell_628 ( .C (clk), .D (signal_2721), .Q (signal_2722) ) ;
    buf_clk cell_630 ( .C (clk), .D (signal_2723), .Q (signal_2724) ) ;
    buf_clk cell_632 ( .C (clk), .D (signal_2725), .Q (signal_2726) ) ;
    buf_clk cell_634 ( .C (clk), .D (signal_2727), .Q (signal_2728) ) ;
    buf_clk cell_636 ( .C (clk), .D (signal_2729), .Q (signal_2730) ) ;
    buf_clk cell_638 ( .C (clk), .D (signal_2731), .Q (signal_2732) ) ;
    buf_clk cell_640 ( .C (clk), .D (signal_2733), .Q (signal_2734) ) ;
    buf_clk cell_642 ( .C (clk), .D (signal_2735), .Q (signal_2736) ) ;
    buf_clk cell_644 ( .C (clk), .D (signal_2737), .Q (signal_2738) ) ;
    buf_clk cell_646 ( .C (clk), .D (signal_2739), .Q (signal_2740) ) ;
    buf_clk cell_648 ( .C (clk), .D (signal_2741), .Q (signal_2742) ) ;
    buf_clk cell_650 ( .C (clk), .D (signal_2743), .Q (signal_2744) ) ;
    buf_clk cell_652 ( .C (clk), .D (signal_2745), .Q (signal_2746) ) ;
    buf_clk cell_654 ( .C (clk), .D (signal_2747), .Q (signal_2748) ) ;
    buf_clk cell_656 ( .C (clk), .D (signal_2749), .Q (signal_2750) ) ;
    buf_clk cell_658 ( .C (clk), .D (signal_2751), .Q (signal_2752) ) ;
    buf_clk cell_660 ( .C (clk), .D (signal_2753), .Q (signal_2754) ) ;
    buf_clk cell_662 ( .C (clk), .D (signal_2755), .Q (signal_2756) ) ;
    buf_clk cell_664 ( .C (clk), .D (signal_2757), .Q (signal_2758) ) ;
    buf_clk cell_666 ( .C (clk), .D (signal_2759), .Q (signal_2760) ) ;
    buf_clk cell_668 ( .C (clk), .D (signal_2761), .Q (signal_2762) ) ;
    buf_clk cell_670 ( .C (clk), .D (signal_2763), .Q (signal_2764) ) ;
    buf_clk cell_672 ( .C (clk), .D (signal_2765), .Q (signal_2766) ) ;
    buf_clk cell_674 ( .C (clk), .D (signal_2767), .Q (signal_2768) ) ;
    buf_clk cell_676 ( .C (clk), .D (signal_2769), .Q (signal_2770) ) ;
    buf_clk cell_678 ( .C (clk), .D (signal_2771), .Q (signal_2772) ) ;
    buf_clk cell_680 ( .C (clk), .D (signal_2773), .Q (signal_2774) ) ;
    buf_clk cell_682 ( .C (clk), .D (signal_2775), .Q (signal_2776) ) ;
    buf_clk cell_684 ( .C (clk), .D (signal_2777), .Q (signal_2778) ) ;
    buf_clk cell_686 ( .C (clk), .D (signal_2779), .Q (signal_2780) ) ;
    buf_clk cell_688 ( .C (clk), .D (signal_2781), .Q (signal_2782) ) ;
    buf_clk cell_690 ( .C (clk), .D (signal_2783), .Q (signal_2784) ) ;
    buf_clk cell_692 ( .C (clk), .D (signal_2785), .Q (signal_2786) ) ;
    buf_clk cell_694 ( .C (clk), .D (signal_2787), .Q (signal_2788) ) ;
    buf_clk cell_696 ( .C (clk), .D (signal_2789), .Q (signal_2790) ) ;
    buf_clk cell_698 ( .C (clk), .D (signal_2791), .Q (signal_2792) ) ;
    buf_clk cell_700 ( .C (clk), .D (signal_2793), .Q (signal_2794) ) ;
    buf_clk cell_702 ( .C (clk), .D (signal_2795), .Q (signal_2796) ) ;
    buf_clk cell_704 ( .C (clk), .D (signal_2797), .Q (signal_2798) ) ;
    buf_clk cell_706 ( .C (clk), .D (signal_2799), .Q (signal_2800) ) ;
    buf_clk cell_708 ( .C (clk), .D (signal_2801), .Q (signal_2802) ) ;
    buf_clk cell_710 ( .C (clk), .D (signal_2803), .Q (signal_2804) ) ;
    buf_clk cell_712 ( .C (clk), .D (signal_2805), .Q (signal_2806) ) ;
    buf_clk cell_714 ( .C (clk), .D (signal_2807), .Q (signal_2808) ) ;
    buf_clk cell_716 ( .C (clk), .D (signal_2809), .Q (signal_2810) ) ;
    buf_clk cell_718 ( .C (clk), .D (signal_2811), .Q (signal_2812) ) ;
    buf_clk cell_720 ( .C (clk), .D (signal_2813), .Q (signal_2814) ) ;
    buf_clk cell_722 ( .C (clk), .D (signal_2815), .Q (signal_2816) ) ;
    buf_clk cell_724 ( .C (clk), .D (signal_2817), .Q (signal_2818) ) ;
    buf_clk cell_726 ( .C (clk), .D (signal_2819), .Q (signal_2820) ) ;
    buf_clk cell_728 ( .C (clk), .D (signal_2821), .Q (signal_2822) ) ;
    buf_clk cell_730 ( .C (clk), .D (signal_2823), .Q (signal_2824) ) ;
    buf_clk cell_732 ( .C (clk), .D (signal_2825), .Q (signal_2826) ) ;
    buf_clk cell_734 ( .C (clk), .D (signal_2827), .Q (signal_2828) ) ;
    buf_clk cell_736 ( .C (clk), .D (signal_2829), .Q (signal_2830) ) ;
    buf_clk cell_738 ( .C (clk), .D (signal_2831), .Q (signal_2832) ) ;
    buf_clk cell_740 ( .C (clk), .D (signal_2833), .Q (signal_2834) ) ;
    buf_clk cell_742 ( .C (clk), .D (signal_2835), .Q (signal_2836) ) ;
    buf_clk cell_744 ( .C (clk), .D (signal_2837), .Q (signal_2838) ) ;
    buf_clk cell_746 ( .C (clk), .D (signal_2839), .Q (signal_2840) ) ;
    buf_clk cell_748 ( .C (clk), .D (signal_2841), .Q (signal_2842) ) ;
    buf_clk cell_750 ( .C (clk), .D (signal_2843), .Q (signal_2844) ) ;
    buf_clk cell_752 ( .C (clk), .D (signal_2845), .Q (signal_2846) ) ;
    buf_clk cell_754 ( .C (clk), .D (signal_2847), .Q (signal_2848) ) ;
    buf_clk cell_756 ( .C (clk), .D (signal_2849), .Q (signal_2850) ) ;
    buf_clk cell_758 ( .C (clk), .D (signal_2851), .Q (signal_2852) ) ;
    buf_clk cell_760 ( .C (clk), .D (signal_2853), .Q (signal_2854) ) ;
    buf_clk cell_762 ( .C (clk), .D (signal_2855), .Q (signal_2856) ) ;
    buf_clk cell_768 ( .C (clk), .D (signal_2861), .Q (signal_2862) ) ;
    buf_clk cell_776 ( .C (clk), .D (signal_2869), .Q (signal_2870) ) ;
    buf_clk cell_784 ( .C (clk), .D (signal_2877), .Q (signal_2878) ) ;
    buf_clk cell_828 ( .C (clk), .D (signal_2921), .Q (signal_2922) ) ;
    buf_clk cell_838 ( .C (clk), .D (signal_2931), .Q (signal_2932) ) ;
    buf_clk cell_848 ( .C (clk), .D (signal_2941), .Q (signal_2942) ) ;
    buf_clk cell_858 ( .C (clk), .D (signal_2951), .Q (signal_2952) ) ;
    buf_clk cell_870 ( .C (clk), .D (signal_2963), .Q (signal_2964) ) ;
    buf_clk cell_882 ( .C (clk), .D (signal_2975), .Q (signal_2976) ) ;
    buf_clk cell_894 ( .C (clk), .D (signal_2987), .Q (signal_2988) ) ;
    buf_clk cell_908 ( .C (clk), .D (signal_3001), .Q (signal_3002) ) ;
    buf_clk cell_922 ( .C (clk), .D (signal_3015), .Q (signal_3016) ) ;

    /* cells in depth 7 */
    buf_clk cell_769 ( .C (clk), .D (signal_2862), .Q (signal_2863) ) ;
    buf_clk cell_777 ( .C (clk), .D (signal_2870), .Q (signal_2871) ) ;
    buf_clk cell_785 ( .C (clk), .D (signal_2878), .Q (signal_2879) ) ;
    buf_clk cell_787 ( .C (clk), .D (signal_282), .Q (signal_2881) ) ;
    buf_clk cell_789 ( .C (clk), .D (signal_824), .Q (signal_2883) ) ;
    buf_clk cell_791 ( .C (clk), .D (signal_825), .Q (signal_2885) ) ;
    buf_clk cell_793 ( .C (clk), .D (signal_274), .Q (signal_2887) ) ;
    buf_clk cell_795 ( .C (clk), .D (signal_808), .Q (signal_2889) ) ;
    buf_clk cell_797 ( .C (clk), .D (signal_809), .Q (signal_2891) ) ;
    buf_clk cell_799 ( .C (clk), .D (signal_306), .Q (signal_2893) ) ;
    buf_clk cell_801 ( .C (clk), .D (signal_872), .Q (signal_2895) ) ;
    buf_clk cell_803 ( .C (clk), .D (signal_873), .Q (signal_2897) ) ;
    buf_clk cell_805 ( .C (clk), .D (signal_299), .Q (signal_2899) ) ;
    buf_clk cell_807 ( .C (clk), .D (signal_858), .Q (signal_2901) ) ;
    buf_clk cell_809 ( .C (clk), .D (signal_859), .Q (signal_2903) ) ;
    buf_clk cell_811 ( .C (clk), .D (signal_244), .Q (signal_2905) ) ;
    buf_clk cell_813 ( .C (clk), .D (signal_748), .Q (signal_2907) ) ;
    buf_clk cell_815 ( .C (clk), .D (signal_749), .Q (signal_2909) ) ;
    buf_clk cell_817 ( .C (clk), .D (signal_302), .Q (signal_2911) ) ;
    buf_clk cell_819 ( .C (clk), .D (signal_864), .Q (signal_2913) ) ;
    buf_clk cell_821 ( .C (clk), .D (signal_865), .Q (signal_2915) ) ;
    buf_clk cell_829 ( .C (clk), .D (signal_2922), .Q (signal_2923) ) ;
    buf_clk cell_839 ( .C (clk), .D (signal_2932), .Q (signal_2933) ) ;
    buf_clk cell_849 ( .C (clk), .D (signal_2942), .Q (signal_2943) ) ;
    buf_clk cell_859 ( .C (clk), .D (signal_2952), .Q (signal_2953) ) ;
    buf_clk cell_871 ( .C (clk), .D (signal_2964), .Q (signal_2965) ) ;
    buf_clk cell_883 ( .C (clk), .D (signal_2976), .Q (signal_2977) ) ;
    buf_clk cell_895 ( .C (clk), .D (signal_2988), .Q (signal_2989) ) ;
    buf_clk cell_909 ( .C (clk), .D (signal_3002), .Q (signal_3003) ) ;
    buf_clk cell_923 ( .C (clk), .D (signal_3016), .Q (signal_3017) ) ;

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_305 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2712, signal_2710, signal_2708}), .a ({signal_717, signal_716, signal_229}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({signal_901, signal_900, signal_320}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_306 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_895, signal_894, signal_317}), .a ({signal_729, signal_728, signal_235}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_903, signal_902, signal_321}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_307 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_869, signal_868, signal_304}), .a ({signal_843, signal_842, signal_291}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({signal_905, signal_904, signal_322}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_308 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_883, signal_882, signal_311}), .a ({signal_2718, signal_2716, signal_2714}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({signal_907, signal_906, signal_323}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_309 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_685, signal_684, signal_213}), .a ({signal_767, signal_766, signal_253}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({signal_909, signal_908, signal_324}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_310 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_751, signal_750, signal_245}), .a ({signal_855, signal_854, signal_297}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({signal_911, signal_910, signal_325}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_311 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_631, signal_630, signal_186}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({signal_913, signal_912, signal_326}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_312 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2724, signal_2722, signal_2720}), .a ({signal_793, signal_792, signal_266}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({signal_915, signal_914, signal_327}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_313 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_657, signal_656, signal_199}), .a ({signal_711, signal_710, signal_226}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({signal_917, signal_916, signal_328}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_314 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_779, signal_778, signal_259}), .a ({signal_837, signal_836, signal_288}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({signal_919, signal_918, signal_329}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_315 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_841, signal_840, signal_290}), .a ({signal_787, signal_786, signal_263}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({signal_921, signal_920, signal_330}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_316 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_845, signal_844, signal_292}), .a ({signal_895, signal_894, signal_317}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_923, signal_922, signal_331}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_317 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_689, signal_688, signal_215}), .a ({signal_2730, signal_2728, signal_2726}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({signal_925, signal_924, signal_332}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_318 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_703, signal_702, signal_222}), .a ({signal_777, signal_776, signal_258}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({signal_927, signal_926, signal_333}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_319 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_669, signal_668, signal_205}), .a ({signal_2736, signal_2734, signal_2732}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({signal_929, signal_928, signal_334}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_320 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_735, signal_734, signal_238}), .a ({signal_727, signal_726, signal_234}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({signal_931, signal_930, signal_335}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_321 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_697, signal_696, signal_219}), .a ({signal_685, signal_684, signal_213}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({signal_933, signal_932, signal_336}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_322 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_891, signal_890, signal_315}), .a ({signal_823, signal_822, signal_281}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({signal_935, signal_934, signal_337}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_323 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_847, signal_846, signal_293}), .a ({signal_663, signal_662, signal_202}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({signal_937, signal_936, signal_338}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_324 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_887, signal_886, signal_313}), .a ({signal_2742, signal_2740, signal_2738}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({signal_939, signal_938, signal_339}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_325 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_699, signal_698, signal_220}), .a ({signal_717, signal_716, signal_229}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({signal_941, signal_940, signal_340}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_326 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_745, signal_744, signal_243}), .a ({signal_733, signal_732, signal_237}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_943, signal_942, signal_341}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_327 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_743, signal_742, signal_242}), .a ({signal_839, signal_838, signal_289}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({signal_945, signal_944, signal_342}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_328 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_691, signal_690, signal_216}), .a ({signal_893, signal_892, signal_316}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({signal_947, signal_946, signal_343}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_329 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_733, signal_732, signal_237}), .a ({signal_827, signal_826, signal_283}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({signal_949, signal_948, signal_344}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_330 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_899, signal_898, signal_319}), .a ({signal_759, signal_758, signal_249}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({signal_951, signal_950, signal_345}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_331 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_771, signal_770, signal_255}), .a ({signal_745, signal_744, signal_243}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({signal_953, signal_952, signal_346}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_332 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_673, signal_672, signal_207}), .a ({signal_2748, signal_2746, signal_2744}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({signal_955, signal_954, signal_347}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_333 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_801, signal_800, signal_270}), .a ({signal_769, signal_768, signal_254}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({signal_957, signal_956, signal_348}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_334 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_783, signal_782, signal_261}), .a ({signal_891, signal_890, signal_315}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({signal_959, signal_958, signal_349}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_335 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2718, signal_2716, signal_2714}), .a ({signal_759, signal_758, signal_249}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({signal_961, signal_960, signal_350}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_336 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_771, signal_770, signal_255}), .a ({signal_821, signal_820, signal_280}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_963, signal_962, signal_351}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_337 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_723, signal_722, signal_232}), .a ({signal_641, signal_640, signal_191}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({signal_965, signal_964, signal_352}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_338 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_881, signal_880, signal_310}), .a ({signal_845, signal_844, signal_292}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({signal_967, signal_966, signal_353}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_339 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_757, signal_756, signal_248}), .a ({signal_721, signal_720, signal_231}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({signal_969, signal_968, signal_354}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_340 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_861, signal_860, signal_300}), .a ({signal_879, signal_878, signal_309}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({signal_971, signal_970, signal_355}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_341 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_705, signal_704, signal_223}), .a ({signal_831, signal_830, signal_285}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({signal_973, signal_972, signal_356}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_342 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_735, signal_734, signal_238}), .a ({signal_761, signal_760, signal_250}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({signal_975, signal_974, signal_357}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_343 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_731, signal_730, signal_236}), .a ({signal_2754, signal_2752, signal_2750}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({signal_977, signal_976, signal_358}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_344 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_805, signal_804, signal_272}), .a ({signal_723, signal_722, signal_232}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({signal_979, signal_978, signal_359}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_345 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2760, signal_2758, signal_2756}), .a ({signal_869, signal_868, signal_304}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({signal_981, signal_980, signal_360}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_346 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_823, signal_822, signal_281}), .a ({signal_831, signal_830, signal_285}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_983, signal_982, signal_361}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_347 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_643, signal_642, signal_192}), .a ({signal_759, signal_758, signal_249}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({signal_985, signal_984, signal_362}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_348 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_857, signal_856, signal_298}), .a ({signal_2766, signal_2764, signal_2762}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({signal_987, signal_986, signal_363}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_349 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_709, signal_708, signal_225}), .a ({signal_2772, signal_2770, signal_2768}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({signal_989, signal_988, signal_364}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_350 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2748, signal_2746, signal_2744}), .a ({signal_835, signal_834, signal_287}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({signal_991, signal_990, signal_365}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_351 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_707, signal_706, signal_224}), .a ({signal_2778, signal_2776, signal_2774}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({signal_993, signal_992, signal_366}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_352 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_639, signal_638, signal_190}), .a ({signal_2784, signal_2782, signal_2780}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({signal_995, signal_994, signal_367}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_353 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_775, signal_774, signal_257}), .a ({signal_653, signal_652, signal_197}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({signal_997, signal_996, signal_368}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_354 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2790, signal_2788, signal_2786}), .a ({signal_789, signal_788, signal_264}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({signal_999, signal_998, signal_369}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_355 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_785, signal_784, signal_262}), .a ({signal_2796, signal_2794, signal_2792}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({signal_1001, signal_1000, signal_370}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_356 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_637, signal_636, signal_189}), .a ({signal_877, signal_876, signal_308}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_1003, signal_1002, signal_371}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_357 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2712, signal_2710, signal_2708}), .a ({signal_761, signal_760, signal_250}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({signal_1005, signal_1004, signal_372}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_358 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_791, signal_790, signal_265}), .a ({signal_787, signal_786, signal_263}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({signal_1007, signal_1006, signal_373}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_359 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_817, signal_816, signal_278}), .a ({signal_737, signal_736, signal_239}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({signal_1009, signal_1008, signal_374}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_360 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_633, signal_632, signal_187}), .a ({signal_687, signal_686, signal_214}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({signal_1011, signal_1010, signal_375}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_361 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_639, signal_638, signal_190}), .a ({signal_651, signal_650, signal_196}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({signal_1013, signal_1012, signal_376}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_362 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_827, signal_826, signal_283}), .a ({signal_2802, signal_2800, signal_2798}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({signal_1015, signal_1014, signal_377}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_363 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_783, signal_782, signal_261}), .a ({signal_851, signal_850, signal_295}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({signal_1017, signal_1016, signal_378}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_364 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_695, signal_694, signal_218}), .a ({signal_635, signal_634, signal_188}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({signal_1019, signal_1018, signal_379}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_365 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_829, signal_828, signal_284}), .a ({signal_661, signal_660, signal_201}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({signal_1021, signal_1020, signal_380}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_366 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2808, signal_2806, signal_2804}), .a ({signal_807, signal_806, signal_273}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_1023, signal_1022, signal_381}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_367 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2808, signal_2806, signal_2804}), .a ({signal_653, signal_652, signal_197}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({signal_1025, signal_1024, signal_382}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_368 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_659, signal_658, signal_200}), .a ({signal_2814, signal_2812, signal_2810}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({signal_1027, signal_1026, signal_383}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_369 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_867, signal_866, signal_303}), .a ({signal_799, signal_798, signal_269}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({signal_1029, signal_1028, signal_384}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_370 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_757, signal_756, signal_248}), .a ({signal_773, signal_772, signal_256}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({signal_1031, signal_1030, signal_385}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_371 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2802, signal_2800, signal_2798}), .a ({signal_783, signal_782, signal_261}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({signal_1033, signal_1032, signal_386}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_372 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_729, signal_728, signal_235}), .a ({signal_871, signal_870, signal_305}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({signal_1035, signal_1034, signal_387}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_373 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_709, signal_708, signal_225}), .a ({signal_2778, signal_2776, signal_2774}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({signal_1037, signal_1036, signal_388}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_374 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_689, signal_688, signal_215}), .a ({signal_2802, signal_2800, signal_2798}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({signal_1039, signal_1038, signal_389}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_375 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_755, signal_754, signal_247}), .a ({signal_813, signal_812, signal_276}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({signal_1041, signal_1040, signal_390}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_376 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_693, signal_692, signal_217}), .a ({signal_697, signal_696, signal_219}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_1043, signal_1042, signal_391}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_377 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_701, signal_700, signal_221}), .a ({signal_683, signal_682, signal_212}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({signal_1045, signal_1044, signal_392}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_378 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2820, signal_2818, signal_2816}), .a ({signal_765, signal_764, signal_252}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({signal_1047, signal_1046, signal_393}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_379 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_641, signal_640, signal_191}), .a ({signal_665, signal_664, signal_203}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({signal_1049, signal_1048, signal_394}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_380 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_855, signal_854, signal_297}), .a ({signal_731, signal_730, signal_236}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({signal_1051, signal_1050, signal_395}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_381 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_687, signal_686, signal_214}), .a ({signal_2718, signal_2716, signal_2714}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({signal_1053, signal_1052, signal_396}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_382 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_769, signal_768, signal_254}), .a ({signal_637, signal_636, signal_189}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({signal_1055, signal_1054, signal_397}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_383 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_769, signal_768, signal_254}), .a ({signal_697, signal_696, signal_219}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({signal_1057, signal_1056, signal_398}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_384 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_679, signal_678, signal_210}), .a ({signal_643, signal_642, signal_192}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({signal_1059, signal_1058, signal_399}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_385 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_817, signal_816, signal_278}), .a ({signal_795, signal_794, signal_267}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({signal_1061, signal_1060, signal_400}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_386 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_683, signal_682, signal_212}), .a ({signal_689, signal_688, signal_215}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_1063, signal_1062, signal_401}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_387 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_853, signal_852, signal_296}), .a ({signal_803, signal_802, signal_271}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({signal_1065, signal_1064, signal_402}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_388 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2826, signal_2824, signal_2822}), .a ({signal_645, signal_644, signal_193}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({signal_1067, signal_1066, signal_403}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_389 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_677, signal_676, signal_209}), .a ({signal_819, signal_818, signal_279}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({signal_1069, signal_1068, signal_404}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_390 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_763, signal_762, signal_251}), .a ({signal_855, signal_854, signal_297}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({signal_1071, signal_1070, signal_405}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_391 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_665, signal_664, signal_203}), .a ({signal_2832, signal_2830, signal_2828}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({signal_1073, signal_1072, signal_406}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_392 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_745, signal_744, signal_243}), .a ({signal_833, signal_832, signal_286}), .clk (clk), .r ({Fresh[770], Fresh[769], Fresh[768]}), .c ({signal_1075, signal_1074, signal_407}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_393 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_727, signal_726, signal_234}), .a ({signal_2838, signal_2836, signal_2834}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771]}), .c ({signal_1077, signal_1076, signal_408}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_394 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_849, signal_848, signal_294}), .a ({signal_771, signal_770, signal_255}), .clk (clk), .r ({Fresh[776], Fresh[775], Fresh[774]}), .c ({signal_1079, signal_1078, signal_409}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_395 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_727, signal_726, signal_234}), .a ({signal_797, signal_796, signal_268}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777]}), .c ({signal_1081, signal_1080, signal_410}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_396 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_741, signal_740, signal_241}), .a ({signal_2802, signal_2800, signal_2798}), .clk (clk), .r ({Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_1083, signal_1082, signal_411}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_397 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_641, signal_640, signal_191}), .a ({signal_725, signal_724, signal_233}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783]}), .c ({signal_1085, signal_1084, signal_412}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_398 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_787, signal_786, signal_263}), .a ({signal_645, signal_644, signal_193}), .clk (clk), .r ({Fresh[788], Fresh[787], Fresh[786]}), .c ({signal_1087, signal_1086, signal_413}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_399 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_893, signal_892, signal_316}), .a ({signal_697, signal_696, signal_219}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789]}), .c ({signal_1089, signal_1088, signal_414}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_400 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_719, signal_718, signal_230}), .a ({signal_885, signal_884, signal_312}), .clk (clk), .r ({Fresh[794], Fresh[793], Fresh[792]}), .c ({signal_1091, signal_1090, signal_415}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_401 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_815, signal_814, signal_277}), .a ({signal_693, signal_692, signal_217}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795]}), .c ({signal_1093, signal_1092, signal_416}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_402 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_855, signal_854, signal_297}), .a ({signal_867, signal_866, signal_303}), .clk (clk), .r ({Fresh[800], Fresh[799], Fresh[798]}), .c ({signal_1095, signal_1094, signal_417}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_403 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_863, signal_862, signal_301}), .a ({signal_811, signal_810, signal_275}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801]}), .c ({signal_1097, signal_1096, signal_418}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_404 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_789, signal_788, signal_264}), .a ({signal_667, signal_666, signal_204}), .clk (clk), .r ({Fresh[806], Fresh[805], Fresh[804]}), .c ({signal_1099, signal_1098, signal_419}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_405 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_649, signal_648, signal_195}), .a ({signal_703, signal_702, signal_222}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807]}), .c ({signal_1101, signal_1100, signal_420}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_406 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_715, signal_714, signal_228}), .a ({signal_743, signal_742, signal_242}), .clk (clk), .r ({Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_1103, signal_1102, signal_421}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_407 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_765, signal_764, signal_252}), .a ({signal_895, signal_894, signal_317}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813]}), .c ({signal_1105, signal_1104, signal_422}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_408 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_697, signal_696, signal_219}), .a ({signal_633, signal_632, signal_187}), .clk (clk), .r ({Fresh[818], Fresh[817], Fresh[816]}), .c ({signal_1107, signal_1106, signal_423}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_409 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_855, signal_854, signal_297}), .a ({signal_2736, signal_2734, signal_2732}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819]}), .c ({signal_1109, signal_1108, signal_424}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_410 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_633, signal_632, signal_187}), .a ({signal_2844, signal_2842, signal_2840}), .clk (clk), .r ({Fresh[824], Fresh[823], Fresh[822]}), .c ({signal_1111, signal_1110, signal_425}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_411 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_639, signal_638, signal_190}), .a ({signal_713, signal_712, signal_227}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825]}), .c ({signal_1113, signal_1112, signal_426}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_412 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_813, signal_812, signal_276}), .a ({signal_2850, signal_2848, signal_2846}), .clk (clk), .r ({Fresh[830], Fresh[829], Fresh[828]}), .c ({signal_1115, signal_1114, signal_427}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_413 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_743, signal_742, signal_242}), .a ({signal_679, signal_678, signal_210}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831]}), .c ({signal_1117, signal_1116, signal_428}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_414 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_655, signal_654, signal_198}), .a ({signal_673, signal_672, signal_207}), .clk (clk), .r ({Fresh[836], Fresh[835], Fresh[834]}), .c ({signal_1119, signal_1118, signal_429}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_415 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_789, signal_788, signal_264}), .a ({signal_897, signal_896, signal_318}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837]}), .c ({signal_1121, signal_1120, signal_430}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_416 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2844, signal_2842, signal_2840}), .a ({signal_805, signal_804, signal_272}), .clk (clk), .r ({Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_1123, signal_1122, signal_431}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_417 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_857, signal_856, signal_298}), .a ({signal_671, signal_670, signal_206}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843]}), .c ({signal_1125, signal_1124, signal_432}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_418 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_739, signal_738, signal_240}), .a ({signal_629, signal_628, signal_185}), .clk (clk), .r ({Fresh[848], Fresh[847], Fresh[846]}), .c ({signal_1127, signal_1126, signal_433}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_419 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_841, signal_840, signal_290}), .a ({signal_739, signal_738, signal_240}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849]}), .c ({signal_1129, signal_1128, signal_434}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_420 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_889, signal_888, signal_314}), .a ({signal_685, signal_684, signal_213}), .clk (clk), .r ({Fresh[854], Fresh[853], Fresh[852]}), .c ({signal_1131, signal_1130, signal_435}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_421 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_781, signal_780, signal_260}), .a ({signal_693, signal_692, signal_217}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855]}), .c ({signal_1133, signal_1132, signal_436}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_422 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_647, signal_646, signal_194}), .a ({signal_737, signal_736, signal_239}), .clk (clk), .r ({Fresh[860], Fresh[859], Fresh[858]}), .c ({signal_1135, signal_1134, signal_437}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_423 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_681, signal_680, signal_211}), .a ({signal_675, signal_674, signal_208}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861]}), .c ({signal_1137, signal_1136, signal_438}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_424 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_775, signal_774, signal_257}), .a ({signal_679, signal_678, signal_210}), .clk (clk), .r ({Fresh[866], Fresh[865], Fresh[864]}), .c ({signal_1139, signal_1138, signal_439}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_425 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_2856, signal_2854, signal_2852}), .a ({signal_851, signal_850, signal_295}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867]}), .c ({signal_1141, signal_1140, signal_440}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_426 ( .s ({signal_2706, signal_2704, signal_2702}), .b ({signal_875, signal_874, signal_307}), .a ({signal_753, signal_752, signal_246}), .clk (clk), .r ({Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_1143, signal_1142, signal_441}) ) ;
    buf_clk cell_770 ( .C (clk), .D (signal_2863), .Q (signal_2864) ) ;
    buf_clk cell_778 ( .C (clk), .D (signal_2871), .Q (signal_2872) ) ;
    buf_clk cell_786 ( .C (clk), .D (signal_2879), .Q (signal_2880) ) ;
    buf_clk cell_788 ( .C (clk), .D (signal_2881), .Q (signal_2882) ) ;
    buf_clk cell_790 ( .C (clk), .D (signal_2883), .Q (signal_2884) ) ;
    buf_clk cell_792 ( .C (clk), .D (signal_2885), .Q (signal_2886) ) ;
    buf_clk cell_794 ( .C (clk), .D (signal_2887), .Q (signal_2888) ) ;
    buf_clk cell_796 ( .C (clk), .D (signal_2889), .Q (signal_2890) ) ;
    buf_clk cell_798 ( .C (clk), .D (signal_2891), .Q (signal_2892) ) ;
    buf_clk cell_800 ( .C (clk), .D (signal_2893), .Q (signal_2894) ) ;
    buf_clk cell_802 ( .C (clk), .D (signal_2895), .Q (signal_2896) ) ;
    buf_clk cell_804 ( .C (clk), .D (signal_2897), .Q (signal_2898) ) ;
    buf_clk cell_806 ( .C (clk), .D (signal_2899), .Q (signal_2900) ) ;
    buf_clk cell_808 ( .C (clk), .D (signal_2901), .Q (signal_2902) ) ;
    buf_clk cell_810 ( .C (clk), .D (signal_2903), .Q (signal_2904) ) ;
    buf_clk cell_812 ( .C (clk), .D (signal_2905), .Q (signal_2906) ) ;
    buf_clk cell_814 ( .C (clk), .D (signal_2907), .Q (signal_2908) ) ;
    buf_clk cell_816 ( .C (clk), .D (signal_2909), .Q (signal_2910) ) ;
    buf_clk cell_818 ( .C (clk), .D (signal_2911), .Q (signal_2912) ) ;
    buf_clk cell_820 ( .C (clk), .D (signal_2913), .Q (signal_2914) ) ;
    buf_clk cell_822 ( .C (clk), .D (signal_2915), .Q (signal_2916) ) ;
    buf_clk cell_830 ( .C (clk), .D (signal_2923), .Q (signal_2924) ) ;
    buf_clk cell_840 ( .C (clk), .D (signal_2933), .Q (signal_2934) ) ;
    buf_clk cell_850 ( .C (clk), .D (signal_2943), .Q (signal_2944) ) ;
    buf_clk cell_860 ( .C (clk), .D (signal_2953), .Q (signal_2954) ) ;
    buf_clk cell_872 ( .C (clk), .D (signal_2965), .Q (signal_2966) ) ;
    buf_clk cell_884 ( .C (clk), .D (signal_2977), .Q (signal_2978) ) ;
    buf_clk cell_896 ( .C (clk), .D (signal_2989), .Q (signal_2990) ) ;
    buf_clk cell_910 ( .C (clk), .D (signal_3003), .Q (signal_3004) ) ;
    buf_clk cell_924 ( .C (clk), .D (signal_3017), .Q (signal_3018) ) ;

    /* cells in depth 9 */
    buf_clk cell_831 ( .C (clk), .D (signal_2924), .Q (signal_2925) ) ;
    buf_clk cell_841 ( .C (clk), .D (signal_2934), .Q (signal_2935) ) ;
    buf_clk cell_851 ( .C (clk), .D (signal_2944), .Q (signal_2945) ) ;
    buf_clk cell_861 ( .C (clk), .D (signal_2954), .Q (signal_2955) ) ;
    buf_clk cell_873 ( .C (clk), .D (signal_2966), .Q (signal_2967) ) ;
    buf_clk cell_885 ( .C (clk), .D (signal_2978), .Q (signal_2979) ) ;
    buf_clk cell_897 ( .C (clk), .D (signal_2990), .Q (signal_2991) ) ;
    buf_clk cell_911 ( .C (clk), .D (signal_3004), .Q (signal_3005) ) ;
    buf_clk cell_925 ( .C (clk), .D (signal_3018), .Q (signal_3019) ) ;

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_427 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_953, signal_952, signal_346}), .a ({signal_1047, signal_1046, signal_393}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873]}), .c ({signal_1147, signal_1146, signal_442}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_428 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_949, signal_948, signal_344}), .a ({signal_1113, signal_1112, signal_426}), .clk (clk), .r ({Fresh[878], Fresh[877], Fresh[876]}), .c ({signal_1149, signal_1148, signal_443}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_429 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1039, signal_1038, signal_389}), .a ({signal_1071, signal_1070, signal_405}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879]}), .c ({signal_1151, signal_1150, signal_444}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_430 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_989, signal_988, signal_364}), .a ({signal_1133, signal_1132, signal_436}), .clk (clk), .r ({Fresh[884], Fresh[883], Fresh[882]}), .c ({signal_1153, signal_1152, signal_445}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_431 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1127, signal_1126, signal_433}), .a ({signal_1109, signal_1108, signal_424}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885]}), .c ({signal_1155, signal_1154, signal_446}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_432 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_935, signal_934, signal_337}), .a ({signal_1027, signal_1026, signal_383}), .clk (clk), .r ({Fresh[890], Fresh[889], Fresh[888]}), .c ({signal_1157, signal_1156, signal_447}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_433 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_995, signal_994, signal_367}), .a ({signal_1105, signal_1104, signal_422}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891]}), .c ({signal_1159, signal_1158, signal_448}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_434 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_947, signal_946, signal_343}), .a ({signal_1065, signal_1064, signal_402}), .clk (clk), .r ({Fresh[896], Fresh[895], Fresh[894]}), .c ({signal_1161, signal_1160, signal_449}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_435 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1141, signal_1140, signal_440}), .a ({signal_909, signal_908, signal_324}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897]}), .c ({signal_1163, signal_1162, signal_450}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_436 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_979, signal_978, signal_359}), .a ({signal_1143, signal_1142, signal_441}), .clk (clk), .r ({Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_1165, signal_1164, signal_451}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_437 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_975, signal_974, signal_357}), .a ({signal_1025, signal_1024, signal_382}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903]}), .c ({signal_1167, signal_1166, signal_452}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_438 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1045, signal_1044, signal_392}), .a ({signal_1033, signal_1032, signal_386}), .clk (clk), .r ({Fresh[908], Fresh[907], Fresh[906]}), .c ({signal_1169, signal_1168, signal_453}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_439 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_923, signal_922, signal_331}), .a ({signal_1101, signal_1100, signal_420}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909]}), .c ({signal_1171, signal_1170, signal_454}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_440 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1091, signal_1090, signal_415}), .a ({signal_1093, signal_1092, signal_416}), .clk (clk), .r ({Fresh[914], Fresh[913], Fresh[912]}), .c ({signal_1173, signal_1172, signal_455}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_441 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1053, signal_1052, signal_396}), .a ({signal_2886, signal_2884, signal_2882}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915]}), .c ({signal_1175, signal_1174, signal_456}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_442 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1131, signal_1130, signal_435}), .a ({signal_1099, signal_1098, signal_419}), .clk (clk), .r ({Fresh[920], Fresh[919], Fresh[918]}), .c ({signal_1177, signal_1176, signal_457}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_443 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_907, signal_906, signal_323}), .a ({signal_957, signal_956, signal_348}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921]}), .c ({signal_1179, signal_1178, signal_458}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_444 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1059, signal_1058, signal_399}), .a ({signal_2892, signal_2890, signal_2888}), .clk (clk), .r ({Fresh[926], Fresh[925], Fresh[924]}), .c ({signal_1181, signal_1180, signal_459}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_445 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1125, signal_1124, signal_432}), .a ({signal_2898, signal_2896, signal_2894}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927]}), .c ({signal_1183, signal_1182, signal_460}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_446 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1019, signal_1018, signal_379}), .a ({signal_913, signal_912, signal_326}), .clk (clk), .r ({Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_1185, signal_1184, signal_461}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_447 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_997, signal_996, signal_368}), .a ({signal_963, signal_962, signal_351}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933]}), .c ({signal_1187, signal_1186, signal_462}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_448 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_929, signal_928, signal_334}), .a ({signal_1009, signal_1008, signal_374}), .clk (clk), .r ({Fresh[938], Fresh[937], Fresh[936]}), .c ({signal_1189, signal_1188, signal_463}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_449 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1085, signal_1084, signal_412}), .a ({signal_911, signal_910, signal_325}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939]}), .c ({signal_1191, signal_1190, signal_464}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_450 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_983, signal_982, signal_361}), .a ({signal_1063, signal_1062, signal_401}), .clk (clk), .r ({Fresh[944], Fresh[943], Fresh[942]}), .c ({signal_1193, signal_1192, signal_465}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_451 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_915, signal_914, signal_327}), .a ({signal_921, signal_920, signal_330}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945]}), .c ({signal_1195, signal_1194, signal_466}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_452 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_901, signal_900, signal_320}), .a ({signal_951, signal_950, signal_345}), .clk (clk), .r ({Fresh[950], Fresh[949], Fresh[948]}), .c ({signal_1197, signal_1196, signal_467}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_453 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1077, signal_1076, signal_408}), .a ({signal_1137, signal_1136, signal_438}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951]}), .c ({signal_1199, signal_1198, signal_468}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_454 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1121, signal_1120, signal_430}), .a ({signal_1095, signal_1094, signal_417}), .clk (clk), .r ({Fresh[956], Fresh[955], Fresh[954]}), .c ({signal_1201, signal_1200, signal_469}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_455 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1089, signal_1088, signal_414}), .a ({signal_941, signal_940, signal_340}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957]}), .c ({signal_1203, signal_1202, signal_470}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_456 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1003, signal_1002, signal_371}), .a ({signal_2904, signal_2902, signal_2900}), .clk (clk), .r ({Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_1205, signal_1204, signal_471}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_457 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_959, signal_958, signal_349}), .a ({signal_961, signal_960, signal_350}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963]}), .c ({signal_1207, signal_1206, signal_472}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_458 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1029, signal_1028, signal_384}), .a ({signal_1035, signal_1034, signal_387}), .clk (clk), .r ({Fresh[968], Fresh[967], Fresh[966]}), .c ({signal_1209, signal_1208, signal_473}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_459 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1011, signal_1010, signal_375}), .a ({signal_943, signal_942, signal_341}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969]}), .c ({signal_1211, signal_1210, signal_474}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_460 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1037, signal_1036, signal_388}), .a ({signal_1081, signal_1080, signal_410}), .clk (clk), .r ({Fresh[974], Fresh[973], Fresh[972]}), .c ({signal_1213, signal_1212, signal_475}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_461 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_981, signal_980, signal_360}), .a ({signal_1031, signal_1030, signal_385}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975]}), .c ({signal_1215, signal_1214, signal_476}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_462 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1135, signal_1134, signal_437}), .a ({signal_939, signal_938, signal_339}), .clk (clk), .r ({Fresh[980], Fresh[979], Fresh[978]}), .c ({signal_1217, signal_1216, signal_477}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_463 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1067, signal_1066, signal_403}), .a ({signal_925, signal_924, signal_332}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981]}), .c ({signal_1219, signal_1218, signal_478}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_464 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_931, signal_930, signal_335}), .a ({signal_945, signal_944, signal_342}), .clk (clk), .r ({Fresh[986], Fresh[985], Fresh[984]}), .c ({signal_1221, signal_1220, signal_479}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_465 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_933, signal_932, signal_336}), .a ({signal_991, signal_990, signal_365}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987]}), .c ({signal_1223, signal_1222, signal_480}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_466 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_973, signal_972, signal_356}), .a ({signal_1117, signal_1116, signal_428}), .clk (clk), .r ({Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_1225, signal_1224, signal_481}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_467 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_999, signal_998, signal_369}), .a ({signal_1017, signal_1016, signal_378}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993]}), .c ({signal_1227, signal_1226, signal_482}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_468 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1043, signal_1042, signal_391}), .a ({signal_1055, signal_1054, signal_397}), .clk (clk), .r ({Fresh[998], Fresh[997], Fresh[996]}), .c ({signal_1229, signal_1228, signal_483}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_469 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1007, signal_1006, signal_373}), .a ({signal_917, signal_916, signal_328}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999]}), .c ({signal_1231, signal_1230, signal_484}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_470 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1103, signal_1102, signal_421}), .a ({signal_1013, signal_1012, signal_376}), .clk (clk), .r ({Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({signal_1233, signal_1232, signal_485}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_471 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_965, signal_964, signal_352}), .a ({signal_993, signal_992, signal_366}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005]}), .c ({signal_1235, signal_1234, signal_486}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_472 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1123, signal_1122, signal_431}), .a ({signal_1097, signal_1096, signal_418}), .clk (clk), .r ({Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({signal_1237, signal_1236, signal_487}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_473 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1057, signal_1056, signal_398}), .a ({signal_1111, signal_1110, signal_425}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011]}), .c ({signal_1239, signal_1238, signal_488}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_474 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_969, signal_968, signal_354}), .a ({signal_1083, signal_1082, signal_411}), .clk (clk), .r ({Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({signal_1241, signal_1240, signal_489}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_475 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_967, signal_966, signal_353}), .a ({signal_927, signal_926, signal_333}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017]}), .c ({signal_1243, signal_1242, signal_490}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_476 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_985, signal_984, signal_362}), .a ({signal_1023, signal_1022, signal_381}), .clk (clk), .r ({Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_1245, signal_1244, signal_491}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_477 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1021, signal_1020, signal_380}), .a ({signal_1069, signal_1068, signal_404}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023]}), .c ({signal_1247, signal_1246, signal_492}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_478 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_2910, signal_2908, signal_2906}), .a ({signal_987, signal_986, signal_363}), .clk (clk), .r ({Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({signal_1249, signal_1248, signal_493}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_479 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_977, signal_976, signal_358}), .a ({signal_1051, signal_1050, signal_395}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029]}), .c ({signal_1251, signal_1250, signal_494}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_480 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1139, signal_1138, signal_439}), .a ({signal_1119, signal_1118, signal_429}), .clk (clk), .r ({Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({signal_1253, signal_1252, signal_495}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_481 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1075, signal_1074, signal_407}), .a ({signal_905, signal_904, signal_322}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035]}), .c ({signal_1255, signal_1254, signal_496}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_482 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_971, signal_970, signal_355}), .a ({signal_1129, signal_1128, signal_434}), .clk (clk), .r ({Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({signal_1257, signal_1256, signal_497}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_483 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1041, signal_1040, signal_390}), .a ({signal_1079, signal_1078, signal_409}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041]}), .c ({signal_1259, signal_1258, signal_498}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_484 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_919, signal_918, signal_329}), .a ({signal_1015, signal_1014, signal_377}), .clk (clk), .r ({Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({signal_1261, signal_1260, signal_499}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_485 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_903, signal_902, signal_321}), .a ({signal_1107, signal_1106, signal_423}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047]}), .c ({signal_1263, signal_1262, signal_500}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_486 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1087, signal_1086, signal_413}), .a ({signal_1061, signal_1060, signal_400}), .clk (clk), .r ({Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_1265, signal_1264, signal_501}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_487 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1005, signal_1004, signal_372}), .a ({signal_1073, signal_1072, signal_406}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053]}), .c ({signal_1267, signal_1266, signal_502}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_488 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_2916, signal_2914, signal_2912}), .a ({signal_1115, signal_1114, signal_427}), .clk (clk), .r ({Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({signal_1269, signal_1268, signal_503}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_489 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1001, signal_1000, signal_370}), .a ({signal_955, signal_954, signal_347}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059]}), .c ({signal_1271, signal_1270, signal_504}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_490 ( .s ({signal_2880, signal_2872, signal_2864}), .b ({signal_1049, signal_1048, signal_394}), .a ({signal_937, signal_936, signal_338}), .clk (clk), .r ({Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({signal_1273, signal_1272, signal_505}) ) ;
    buf_clk cell_832 ( .C (clk), .D (signal_2925), .Q (signal_2926) ) ;
    buf_clk cell_842 ( .C (clk), .D (signal_2935), .Q (signal_2936) ) ;
    buf_clk cell_852 ( .C (clk), .D (signal_2945), .Q (signal_2946) ) ;
    buf_clk cell_862 ( .C (clk), .D (signal_2955), .Q (signal_2956) ) ;
    buf_clk cell_874 ( .C (clk), .D (signal_2967), .Q (signal_2968) ) ;
    buf_clk cell_886 ( .C (clk), .D (signal_2979), .Q (signal_2980) ) ;
    buf_clk cell_898 ( .C (clk), .D (signal_2991), .Q (signal_2992) ) ;
    buf_clk cell_912 ( .C (clk), .D (signal_3005), .Q (signal_3006) ) ;
    buf_clk cell_926 ( .C (clk), .D (signal_3019), .Q (signal_3020) ) ;

    /* cells in depth 11 */
    buf_clk cell_863 ( .C (clk), .D (signal_2956), .Q (signal_2957) ) ;
    buf_clk cell_875 ( .C (clk), .D (signal_2968), .Q (signal_2969) ) ;
    buf_clk cell_887 ( .C (clk), .D (signal_2980), .Q (signal_2981) ) ;
    buf_clk cell_899 ( .C (clk), .D (signal_2992), .Q (signal_2993) ) ;
    buf_clk cell_913 ( .C (clk), .D (signal_3006), .Q (signal_3007) ) ;
    buf_clk cell_927 ( .C (clk), .D (signal_3020), .Q (signal_3021) ) ;

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_491 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1213, signal_1212, signal_475}), .a ({signal_1151, signal_1150, signal_444}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065]}), .c ({signal_1277, signal_1276, signal_506}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_492 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1163, signal_1162, signal_450}), .a ({signal_1173, signal_1172, signal_455}), .clk (clk), .r ({Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({signal_1279, signal_1278, signal_507}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_493 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1241, signal_1240, signal_489}), .a ({signal_1203, signal_1202, signal_470}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071]}), .c ({signal_1281, signal_1280, signal_508}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_494 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1229, signal_1228, signal_483}), .a ({signal_1153, signal_1152, signal_445}), .clk (clk), .r ({Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({signal_1283, signal_1282, signal_509}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_495 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1261, signal_1260, signal_499}), .a ({signal_1177, signal_1176, signal_457}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077]}), .c ({signal_1285, signal_1284, signal_510}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_496 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1223, signal_1222, signal_480}), .a ({signal_1219, signal_1218, signal_478}), .clk (clk), .r ({Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_1287, signal_1286, signal_511}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_497 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1265, signal_1264, signal_501}), .a ({signal_1215, signal_1214, signal_476}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083]}), .c ({signal_1289, signal_1288, signal_512}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_498 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1243, signal_1242, signal_490}), .a ({signal_1199, signal_1198, signal_468}), .clk (clk), .r ({Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({signal_1291, signal_1290, signal_513}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_499 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1269, signal_1268, signal_503}), .a ({signal_1185, signal_1184, signal_461}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089]}), .c ({signal_1293, signal_1292, signal_514}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_500 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1179, signal_1178, signal_458}), .a ({signal_1187, signal_1186, signal_462}), .clk (clk), .r ({Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({signal_1295, signal_1294, signal_515}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_501 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1161, signal_1160, signal_449}), .a ({signal_1197, signal_1196, signal_467}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095]}), .c ({signal_1297, signal_1296, signal_516}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_502 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1259, signal_1258, signal_498}), .a ({signal_1245, signal_1244, signal_491}), .clk (clk), .r ({Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({signal_1299, signal_1298, signal_517}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_503 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1167, signal_1166, signal_452}), .a ({signal_1239, signal_1238, signal_488}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101]}), .c ({signal_1301, signal_1300, signal_518}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_504 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1247, signal_1246, signal_492}), .a ({signal_1201, signal_1200, signal_469}), .clk (clk), .r ({Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({signal_1303, signal_1302, signal_519}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_505 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1253, signal_1252, signal_495}), .a ({signal_1207, signal_1206, signal_472}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107]}), .c ({signal_1305, signal_1304, signal_520}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_506 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1255, signal_1254, signal_496}), .a ({signal_1191, signal_1190, signal_464}), .clk (clk), .r ({Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_1307, signal_1306, signal_521}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_507 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1251, signal_1250, signal_494}), .a ({signal_1183, signal_1182, signal_460}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113]}), .c ({signal_1309, signal_1308, signal_522}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_508 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1209, signal_1208, signal_473}), .a ({signal_1257, signal_1256, signal_497}), .clk (clk), .r ({Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({signal_1311, signal_1310, signal_523}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_509 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1249, signal_1248, signal_493}), .a ({signal_1181, signal_1180, signal_459}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119]}), .c ({signal_1313, signal_1312, signal_524}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_510 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1171, signal_1170, signal_454}), .a ({signal_1267, signal_1266, signal_502}), .clk (clk), .r ({Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({signal_1315, signal_1314, signal_525}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_511 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1271, signal_1270, signal_504}), .a ({signal_1221, signal_1220, signal_479}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125]}), .c ({signal_1317, signal_1316, signal_526}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_512 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1175, signal_1174, signal_456}), .a ({signal_1157, signal_1156, signal_447}), .clk (clk), .r ({Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({signal_1319, signal_1318, signal_527}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_513 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1155, signal_1154, signal_446}), .a ({signal_1195, signal_1194, signal_466}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131]}), .c ({signal_1321, signal_1320, signal_528}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_514 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1205, signal_1204, signal_471}), .a ({signal_1233, signal_1232, signal_485}), .clk (clk), .r ({Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({signal_1323, signal_1322, signal_529}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_515 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1227, signal_1226, signal_482}), .a ({signal_1165, signal_1164, signal_451}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137]}), .c ({signal_1325, signal_1324, signal_530}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_516 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1159, signal_1158, signal_448}), .a ({signal_1189, signal_1188, signal_463}), .clk (clk), .r ({Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_1327, signal_1326, signal_531}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_517 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1193, signal_1192, signal_465}), .a ({signal_1273, signal_1272, signal_505}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143]}), .c ({signal_1329, signal_1328, signal_532}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_518 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1169, signal_1168, signal_453}), .a ({signal_1263, signal_1262, signal_500}), .clk (clk), .r ({Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({signal_1331, signal_1330, signal_533}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_519 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1211, signal_1210, signal_474}), .a ({signal_1225, signal_1224, signal_481}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149]}), .c ({signal_1333, signal_1332, signal_534}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_520 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1217, signal_1216, signal_477}), .a ({signal_1231, signal_1230, signal_484}), .clk (clk), .r ({Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({signal_1335, signal_1334, signal_535}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_521 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1237, signal_1236, signal_487}), .a ({signal_1147, signal_1146, signal_442}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155]}), .c ({signal_1337, signal_1336, signal_536}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_522 ( .s ({signal_2946, signal_2936, signal_2926}), .b ({signal_1235, signal_1234, signal_486}), .a ({signal_1149, signal_1148, signal_443}), .clk (clk), .r ({Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({signal_1339, signal_1338, signal_537}) ) ;
    buf_clk cell_864 ( .C (clk), .D (signal_2957), .Q (signal_2958) ) ;
    buf_clk cell_876 ( .C (clk), .D (signal_2969), .Q (signal_2970) ) ;
    buf_clk cell_888 ( .C (clk), .D (signal_2981), .Q (signal_2982) ) ;
    buf_clk cell_900 ( .C (clk), .D (signal_2993), .Q (signal_2994) ) ;
    buf_clk cell_914 ( .C (clk), .D (signal_3007), .Q (signal_3008) ) ;
    buf_clk cell_928 ( .C (clk), .D (signal_3021), .Q (signal_3022) ) ;

    /* cells in depth 13 */
    buf_clk cell_901 ( .C (clk), .D (signal_2994), .Q (signal_2995) ) ;
    buf_clk cell_915 ( .C (clk), .D (signal_3008), .Q (signal_3009) ) ;
    buf_clk cell_929 ( .C (clk), .D (signal_3022), .Q (signal_3023) ) ;

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_523 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1327, signal_1326, signal_531}), .a ({signal_1301, signal_1300, signal_518}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161]}), .c ({signal_1343, signal_1342, signal_538}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_524 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1281, signal_1280, signal_508}), .a ({signal_1335, signal_1334, signal_535}), .clk (clk), .r ({Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({signal_1345, signal_1344, signal_539}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_525 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1313, signal_1312, signal_524}), .a ({signal_1311, signal_1310, signal_523}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167]}), .c ({signal_1347, signal_1346, signal_540}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_526 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1303, signal_1302, signal_519}), .a ({signal_1319, signal_1318, signal_527}), .clk (clk), .r ({Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_1349, signal_1348, signal_541}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_527 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1321, signal_1320, signal_528}), .a ({signal_1277, signal_1276, signal_506}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173]}), .c ({signal_1351, signal_1350, signal_542}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_528 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1317, signal_1316, signal_526}), .a ({signal_1339, signal_1338, signal_537}), .clk (clk), .r ({Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({signal_1353, signal_1352, signal_543}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_529 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1285, signal_1284, signal_510}), .a ({signal_1331, signal_1330, signal_533}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179]}), .c ({signal_1355, signal_1354, signal_544}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_530 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1279, signal_1278, signal_507}), .a ({signal_1287, signal_1286, signal_511}), .clk (clk), .r ({Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({signal_1357, signal_1356, signal_545}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_531 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1293, signal_1292, signal_514}), .a ({signal_1297, signal_1296, signal_516}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185]}), .c ({signal_1359, signal_1358, signal_546}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_532 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1305, signal_1304, signal_520}), .a ({signal_1315, signal_1314, signal_525}), .clk (clk), .r ({Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({signal_1361, signal_1360, signal_547}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_533 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1289, signal_1288, signal_512}), .a ({signal_1325, signal_1324, signal_530}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191]}), .c ({signal_1363, signal_1362, signal_548}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_534 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1295, signal_1294, signal_515}), .a ({signal_1333, signal_1332, signal_534}), .clk (clk), .r ({Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({signal_1365, signal_1364, signal_549}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_535 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1307, signal_1306, signal_521}), .a ({signal_1299, signal_1298, signal_517}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197]}), .c ({signal_1367, signal_1366, signal_550}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_536 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1323, signal_1322, signal_529}), .a ({signal_1337, signal_1336, signal_536}), .clk (clk), .r ({Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_1369, signal_1368, signal_551}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_537 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1291, signal_1290, signal_513}), .a ({signal_1329, signal_1328, signal_532}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203]}), .c ({signal_1371, signal_1370, signal_552}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_538 ( .s ({signal_2982, signal_2970, signal_2958}), .b ({signal_1283, signal_1282, signal_509}), .a ({signal_1309, signal_1308, signal_522}), .clk (clk), .r ({Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({signal_1373, signal_1372, signal_553}) ) ;
    buf_clk cell_902 ( .C (clk), .D (signal_2995), .Q (signal_2996) ) ;
    buf_clk cell_916 ( .C (clk), .D (signal_3009), .Q (signal_3010) ) ;
    buf_clk cell_930 ( .C (clk), .D (signal_3023), .Q (signal_3024) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_539 ( .s ({signal_3024, signal_3010, signal_2996}), .b ({signal_1345, signal_1344, signal_539}), .a ({signal_1357, signal_1356, signal_545}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209]}), .c ({signal_1377, signal_1376, signal_145}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_540 ( .s ({signal_3024, signal_3010, signal_2996}), .b ({signal_1363, signal_1362, signal_548}), .a ({signal_1359, signal_1358, signal_546}), .clk (clk), .r ({Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({signal_1379, signal_1378, signal_148}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_541 ( .s ({signal_3024, signal_3010, signal_2996}), .b ({signal_1353, signal_1352, signal_543}), .a ({signal_1361, signal_1360, signal_547}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215]}), .c ({signal_1381, signal_1380, signal_143}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_542 ( .s ({signal_3024, signal_3010, signal_2996}), .b ({signal_1373, signal_1372, signal_553}), .a ({signal_1369, signal_1368, signal_551}), .clk (clk), .r ({Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({signal_1383, signal_1382, signal_146}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_543 ( .s ({signal_3024, signal_3010, signal_2996}), .b ({signal_1347, signal_1346, signal_540}), .a ({signal_1371, signal_1370, signal_552}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221]}), .c ({signal_1385, signal_1384, signal_149}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_544 ( .s ({signal_3024, signal_3010, signal_2996}), .b ({signal_1367, signal_1366, signal_550}), .a ({signal_1351, signal_1350, signal_542}), .clk (clk), .r ({Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({signal_1387, signal_1386, signal_144}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_545 ( .s ({signal_3024, signal_3010, signal_2996}), .b ({signal_1343, signal_1342, signal_538}), .a ({signal_1365, signal_1364, signal_549}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227]}), .c ({signal_1389, signal_1388, signal_147}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_546 ( .s ({signal_3024, signal_3010, signal_2996}), .b ({signal_1355, signal_1354, signal_544}), .a ({signal_1349, signal_1348, signal_541}), .clk (clk), .r ({Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({signal_1391, signal_1390, signal_150}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_1381, signal_1380, signal_143}), .Q ({Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_1387, signal_1386, signal_144}), .Q ({Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_1377, signal_1376, signal_145}), .Q ({Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_1383, signal_1382, signal_146}), .Q ({Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_4 ( .clk (clk), .D ({signal_1389, signal_1388, signal_147}), .Q ({Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_5 ( .clk (clk), .D ({signal_1379, signal_1378, signal_148}), .Q ({Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_6 ( .clk (clk), .D ({signal_1385, signal_1384, signal_149}), .Q ({Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_7 ( .clk (clk), .D ({signal_1391, signal_1390, signal_150}), .Q ({Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
