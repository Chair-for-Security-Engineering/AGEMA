/* modified netlist. Source: module AES in file /AES_round-based/AGEMA/AES.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module AES_GHPC_ANF_ClockGating_d1 (plaintext_s0, key_s0, clk, reset, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [159:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_423 ;
    wire signal_425 ;
    wire signal_427 ;
    wire signal_429 ;
    wire signal_431 ;
    wire signal_433 ;
    wire signal_435 ;
    wire signal_437 ;
    wire signal_439 ;
    wire signal_441 ;
    wire signal_443 ;
    wire signal_445 ;
    wire signal_447 ;
    wire signal_449 ;
    wire signal_451 ;
    wire signal_453 ;
    wire signal_455 ;
    wire signal_457 ;
    wire signal_459 ;
    wire signal_461 ;
    wire signal_463 ;
    wire signal_465 ;
    wire signal_467 ;
    wire signal_469 ;
    wire signal_471 ;
    wire signal_473 ;
    wire signal_475 ;
    wire signal_477 ;
    wire signal_479 ;
    wire signal_481 ;
    wire signal_483 ;
    wire signal_485 ;
    wire signal_487 ;
    wire signal_489 ;
    wire signal_491 ;
    wire signal_493 ;
    wire signal_495 ;
    wire signal_497 ;
    wire signal_499 ;
    wire signal_501 ;
    wire signal_503 ;
    wire signal_505 ;
    wire signal_507 ;
    wire signal_509 ;
    wire signal_511 ;
    wire signal_513 ;
    wire signal_515 ;
    wire signal_517 ;
    wire signal_519 ;
    wire signal_521 ;
    wire signal_523 ;
    wire signal_525 ;
    wire signal_527 ;
    wire signal_529 ;
    wire signal_531 ;
    wire signal_533 ;
    wire signal_535 ;
    wire signal_537 ;
    wire signal_539 ;
    wire signal_541 ;
    wire signal_543 ;
    wire signal_545 ;
    wire signal_547 ;
    wire signal_549 ;
    wire signal_551 ;
    wire signal_553 ;
    wire signal_555 ;
    wire signal_557 ;
    wire signal_559 ;
    wire signal_561 ;
    wire signal_563 ;
    wire signal_565 ;
    wire signal_567 ;
    wire signal_569 ;
    wire signal_571 ;
    wire signal_573 ;
    wire signal_575 ;
    wire signal_577 ;
    wire signal_579 ;
    wire signal_581 ;
    wire signal_583 ;
    wire signal_585 ;
    wire signal_587 ;
    wire signal_589 ;
    wire signal_591 ;
    wire signal_593 ;
    wire signal_595 ;
    wire signal_597 ;
    wire signal_599 ;
    wire signal_601 ;
    wire signal_603 ;
    wire signal_605 ;
    wire signal_607 ;
    wire signal_609 ;
    wire signal_611 ;
    wire signal_613 ;
    wire signal_615 ;
    wire signal_617 ;
    wire signal_619 ;
    wire signal_621 ;
    wire signal_623 ;
    wire signal_625 ;
    wire signal_627 ;
    wire signal_629 ;
    wire signal_631 ;
    wire signal_633 ;
    wire signal_635 ;
    wire signal_637 ;
    wire signal_639 ;
    wire signal_641 ;
    wire signal_643 ;
    wire signal_645 ;
    wire signal_647 ;
    wire signal_649 ;
    wire signal_651 ;
    wire signal_653 ;
    wire signal_655 ;
    wire signal_657 ;
    wire signal_659 ;
    wire signal_661 ;
    wire signal_663 ;
    wire signal_665 ;
    wire signal_667 ;
    wire signal_669 ;
    wire signal_671 ;
    wire signal_673 ;
    wire signal_675 ;
    wire signal_792 ;
    wire signal_912 ;
    wire signal_1032 ;
    wire signal_1152 ;
    wire signal_1272 ;
    wire signal_1392 ;
    wire signal_1512 ;
    wire signal_1632 ;
    wire signal_1752 ;
    wire signal_1872 ;
    wire signal_1992 ;
    wire signal_2112 ;
    wire signal_2232 ;
    wire signal_2352 ;
    wire signal_2472 ;
    wire signal_2592 ;
    wire signal_2597 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2855 ;
    wire signal_2857 ;
    wire signal_2859 ;
    wire signal_2861 ;
    wire signal_2863 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2877 ;
    wire signal_2879 ;
    wire signal_2881 ;
    wire signal_2883 ;
    wire signal_2885 ;
    wire signal_2887 ;
    wire signal_2889 ;
    wire signal_2891 ;
    wire signal_2893 ;
    wire signal_2895 ;
    wire signal_2897 ;
    wire signal_2899 ;
    wire signal_2901 ;
    wire signal_2903 ;
    wire signal_2905 ;
    wire signal_2907 ;
    wire signal_2909 ;
    wire signal_2911 ;
    wire signal_2913 ;
    wire signal_2915 ;
    wire signal_2917 ;
    wire signal_2919 ;
    wire signal_2921 ;
    wire signal_2923 ;
    wire signal_2925 ;
    wire signal_2927 ;
    wire signal_2929 ;
    wire signal_2931 ;
    wire signal_2933 ;
    wire signal_2935 ;
    wire signal_2937 ;
    wire signal_2939 ;
    wire signal_2941 ;
    wire signal_2943 ;
    wire signal_2945 ;
    wire signal_2947 ;
    wire signal_2949 ;
    wire signal_2951 ;
    wire signal_2953 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2959 ;
    wire signal_2961 ;
    wire signal_2963 ;
    wire signal_2965 ;
    wire signal_2967 ;
    wire signal_2969 ;
    wire signal_2971 ;
    wire signal_2973 ;
    wire signal_2975 ;
    wire signal_2977 ;
    wire signal_2979 ;
    wire signal_2981 ;
    wire signal_2983 ;
    wire signal_2985 ;
    wire signal_2987 ;
    wire signal_2989 ;
    wire signal_2991 ;
    wire signal_2993 ;
    wire signal_2995 ;
    wire signal_2997 ;
    wire signal_2999 ;
    wire signal_3001 ;
    wire signal_3003 ;
    wire signal_3005 ;
    wire signal_3007 ;
    wire signal_3009 ;
    wire signal_3011 ;
    wire signal_3013 ;
    wire signal_3015 ;
    wire signal_3017 ;
    wire signal_3019 ;
    wire signal_3021 ;
    wire signal_3023 ;
    wire signal_3025 ;
    wire signal_3027 ;
    wire signal_3029 ;
    wire signal_3031 ;
    wire signal_3033 ;
    wire signal_3035 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3043 ;
    wire signal_3045 ;
    wire signal_3047 ;
    wire signal_3049 ;
    wire signal_3051 ;
    wire signal_3053 ;
    wire signal_3055 ;
    wire signal_3057 ;
    wire signal_3059 ;
    wire signal_3061 ;
    wire signal_3063 ;
    wire signal_3065 ;
    wire signal_3067 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3079 ;
    wire signal_3081 ;
    wire signal_3083 ;
    wire signal_3085 ;
    wire signal_3087 ;
    wire signal_3089 ;
    wire signal_3091 ;
    wire signal_3093 ;
    wire signal_3095 ;
    wire signal_3097 ;
    wire signal_3099 ;
    wire signal_3101 ;
    wire signal_3103 ;
    wire signal_3105 ;
    wire signal_3107 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3874 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3882 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3890 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3898 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3906 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3914 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3922 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3930 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3938 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3946 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3954 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3962 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3970 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3978 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3986 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4394 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4402 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4410 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4418 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4426 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4434 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4442 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4450 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4458 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4466 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4474 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4482 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4490 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4498 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4506 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4514 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5403 ;
    wire signal_5405 ;
    wire signal_5407 ;
    wire signal_5409 ;
    wire signal_5411 ;
    wire signal_5413 ;
    wire signal_5415 ;
    wire signal_5417 ;
    wire signal_5419 ;
    wire signal_5421 ;
    wire signal_5423 ;
    wire signal_5425 ;
    wire signal_5427 ;
    wire signal_5429 ;
    wire signal_5431 ;
    wire signal_5433 ;
    wire signal_5435 ;
    wire signal_5437 ;
    wire signal_5439 ;
    wire signal_5441 ;
    wire signal_5443 ;
    wire signal_5445 ;
    wire signal_5447 ;
    wire signal_5449 ;
    wire signal_5451 ;
    wire signal_5453 ;
    wire signal_5455 ;
    wire signal_5457 ;
    wire signal_5459 ;
    wire signal_5461 ;
    wire signal_5463 ;
    wire signal_5465 ;
    wire signal_5467 ;
    wire signal_5469 ;
    wire signal_5471 ;
    wire signal_5473 ;
    wire signal_5475 ;
    wire signal_5477 ;
    wire signal_5479 ;
    wire signal_5481 ;
    wire signal_5483 ;
    wire signal_5485 ;
    wire signal_5487 ;
    wire signal_5489 ;
    wire signal_5491 ;
    wire signal_5493 ;
    wire signal_5495 ;
    wire signal_5497 ;
    wire signal_5499 ;
    wire signal_5501 ;
    wire signal_5503 ;
    wire signal_5505 ;
    wire signal_5507 ;
    wire signal_5509 ;
    wire signal_5511 ;
    wire signal_5513 ;
    wire signal_5515 ;
    wire signal_5517 ;
    wire signal_5519 ;
    wire signal_5521 ;
    wire signal_5523 ;
    wire signal_5525 ;
    wire signal_5527 ;
    wire signal_5529 ;
    wire signal_5531 ;
    wire signal_5533 ;
    wire signal_5535 ;
    wire signal_5537 ;
    wire signal_5539 ;
    wire signal_5541 ;
    wire signal_5543 ;
    wire signal_5545 ;
    wire signal_5547 ;
    wire signal_5549 ;
    wire signal_5551 ;
    wire signal_5553 ;
    wire signal_5555 ;
    wire signal_5557 ;
    wire signal_5559 ;
    wire signal_5561 ;
    wire signal_5563 ;
    wire signal_5565 ;
    wire signal_5567 ;
    wire signal_5569 ;
    wire signal_5571 ;
    wire signal_5573 ;
    wire signal_5575 ;
    wire signal_5577 ;
    wire signal_5579 ;
    wire signal_5581 ;
    wire signal_5583 ;
    wire signal_5585 ;
    wire signal_5587 ;
    wire signal_5589 ;
    wire signal_5591 ;
    wire signal_5593 ;
    wire signal_5595 ;
    wire signal_5597 ;
    wire signal_5599 ;
    wire signal_5601 ;
    wire signal_5603 ;
    wire signal_5605 ;
    wire signal_5607 ;
    wire signal_5609 ;
    wire signal_5611 ;
    wire signal_5613 ;
    wire signal_5615 ;
    wire signal_5617 ;
    wire signal_5619 ;
    wire signal_5621 ;
    wire signal_5623 ;
    wire signal_5625 ;
    wire signal_5627 ;
    wire signal_5629 ;
    wire signal_5631 ;
    wire signal_5633 ;
    wire signal_5635 ;
    wire signal_5637 ;
    wire signal_5639 ;
    wire signal_5641 ;
    wire signal_5643 ;
    wire signal_5645 ;
    wire signal_5647 ;
    wire signal_5649 ;
    wire signal_5651 ;
    wire signal_5653 ;
    wire signal_5655 ;
    wire signal_5657 ;
    wire signal_5659 ;
    wire signal_5661 ;
    wire signal_5663 ;
    wire signal_5665 ;
    wire signal_5667 ;
    wire signal_5669 ;
    wire signal_5671 ;
    wire signal_5673 ;
    wire signal_5675 ;
    wire signal_5677 ;
    wire signal_5679 ;
    wire signal_5681 ;
    wire signal_5683 ;
    wire signal_5685 ;
    wire signal_5687 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5723 ;
    wire signal_5725 ;
    wire signal_5727 ;
    wire signal_5729 ;
    wire signal_5731 ;
    wire signal_5733 ;
    wire signal_5735 ;
    wire signal_5737 ;
    wire signal_5739 ;
    wire signal_5741 ;
    wire signal_5743 ;
    wire signal_5745 ;
    wire signal_5747 ;
    wire signal_5749 ;
    wire signal_5751 ;
    wire signal_5753 ;
    wire signal_5755 ;
    wire signal_5757 ;
    wire signal_5759 ;
    wire signal_5761 ;
    wire signal_5763 ;
    wire signal_5765 ;
    wire signal_5767 ;
    wire signal_5769 ;
    wire signal_5771 ;
    wire signal_5773 ;
    wire signal_5775 ;
    wire signal_5777 ;
    wire signal_5779 ;
    wire signal_5781 ;
    wire signal_5783 ;
    wire signal_5785 ;
    wire signal_5787 ;
    wire signal_5789 ;
    wire signal_5791 ;
    wire signal_5793 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5829 ;
    wire signal_5831 ;
    wire signal_5833 ;
    wire signal_5835 ;
    wire signal_5837 ;
    wire signal_5839 ;
    wire signal_5841 ;
    wire signal_5843 ;
    wire signal_5845 ;
    wire signal_5847 ;
    wire signal_5849 ;
    wire signal_5851 ;
    wire signal_5853 ;
    wire signal_5855 ;
    wire signal_5857 ;
    wire signal_5859 ;
    wire signal_5861 ;
    wire signal_5863 ;
    wire signal_5865 ;
    wire signal_5867 ;
    wire signal_5869 ;
    wire signal_5871 ;
    wire signal_5873 ;
    wire signal_5875 ;
    wire signal_5877 ;
    wire signal_5879 ;
    wire signal_5881 ;
    wire signal_5883 ;
    wire signal_5885 ;
    wire signal_5887 ;
    wire signal_5889 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5925 ;
    wire signal_5927 ;
    wire signal_5929 ;
    wire signal_5931 ;
    wire signal_5933 ;
    wire signal_5935 ;
    wire signal_5937 ;
    wire signal_5939 ;
    wire signal_5941 ;
    wire signal_5943 ;
    wire signal_5945 ;
    wire signal_5947 ;
    wire signal_5949 ;
    wire signal_5951 ;
    wire signal_5953 ;
    wire signal_5955 ;
    wire signal_5957 ;
    wire signal_5959 ;
    wire signal_5961 ;
    wire signal_5963 ;
    wire signal_5965 ;
    wire signal_5967 ;
    wire signal_5969 ;
    wire signal_5971 ;
    wire signal_5973 ;
    wire signal_5975 ;
    wire signal_5977 ;
    wire signal_5979 ;
    wire signal_5981 ;
    wire signal_5983 ;
    wire signal_5985 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5997 ;
    wire signal_5999 ;
    wire signal_6001 ;
    wire signal_6003 ;
    wire signal_6005 ;
    wire signal_6007 ;
    wire signal_6009 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6016 ;
    wire signal_6018 ;
    wire signal_6020 ;
    wire signal_6181 ;

    /* cells in depth 0 */
    INV_X1 cell_0 ( .A (signal_395), .ZN (signal_400) ) ;
    INV_X1 cell_1 ( .A (signal_395), .ZN (signal_401) ) ;
    INV_X1 cell_2 ( .A (signal_395), .ZN (signal_398) ) ;
    INV_X1 cell_3 ( .A (signal_395), .ZN (signal_396) ) ;
    INV_X1 cell_4 ( .A (signal_395), .ZN (signal_397) ) ;
    INV_X1 cell_5 ( .A (signal_395), .ZN (signal_399) ) ;
    NOR2_X1 cell_6 ( .A1 (signal_406), .A2 (signal_411), .ZN (signal_395) ) ;
    INV_X1 cell_7 ( .A (signal_4388), .ZN (signal_406) ) ;
    INV_X1 cell_8 ( .A (signal_395), .ZN (signal_402) ) ;
    NOR2_X1 cell_9 ( .A1 (signal_4386), .A2 (signal_4387), .ZN (signal_404) ) ;
    INV_X1 cell_10 ( .A (signal_404), .ZN (signal_403) ) ;
    NOR2_X1 cell_11 ( .A1 (signal_4388), .A2 (signal_403), .ZN (signal_4384) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_4388), .A2 (signal_4385), .ZN (signal_418) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_418), .A2 (signal_403), .ZN (signal_4383) ) ;
    NAND2_X1 cell_14 ( .A1 (signal_4385), .A2 (signal_404), .ZN (signal_411) ) ;
    INV_X1 cell_15 ( .A (signal_4386), .ZN (signal_409) ) ;
    AND2_X1 cell_16 ( .A1 (signal_409), .A2 (signal_4387), .ZN (signal_414) ) ;
    NAND2_X1 cell_17 ( .A1 (signal_418), .A2 (signal_414), .ZN (signal_405) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_402), .A2 (signal_405), .ZN (signal_4382) ) ;
    NOR2_X1 cell_19 ( .A1 (signal_4385), .A2 (signal_406), .ZN (signal_416) ) ;
    NAND2_X1 cell_20 ( .A1 (signal_414), .A2 (signal_416), .ZN (signal_408) ) ;
    NAND2_X1 cell_21 ( .A1 (signal_4385), .A2 (signal_4384), .ZN (signal_407) ) ;
    NAND2_X1 cell_22 ( .A1 (signal_408), .A2 (signal_407), .ZN (signal_4381) ) ;
    NOR2_X1 cell_23 ( .A1 (signal_4387), .A2 (signal_409), .ZN (signal_412) ) ;
    NAND2_X1 cell_24 ( .A1 (signal_418), .A2 (signal_412), .ZN (signal_410) ) ;
    NAND2_X1 cell_25 ( .A1 (signal_411), .A2 (signal_410), .ZN (signal_4380) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_416), .A2 (signal_412), .ZN (signal_413) ) ;
    NAND2_X1 cell_27 ( .A1 (signal_402), .A2 (signal_413), .ZN (signal_4379) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_156 ( .a ({signal_4549, signal_3870}), .b ({signal_4550, signal_4378}), .c ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_157 ( .a ({signal_4552, signal_3770}), .b ({signal_4553, signal_4278}), .c ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_158 ( .a ({signal_4555, signal_3769}), .b ({signal_4556, signal_4277}), .c ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_159 ( .a ({signal_4558, signal_3768}), .b ({signal_4559, signal_4276}), .c ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_160 ( .a ({signal_4561, signal_3767}), .b ({signal_4562, signal_4275}), .c ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_161 ( .a ({signal_4564, signal_3766}), .b ({signal_4565, signal_4274}), .c ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_162 ( .a ({signal_4567, signal_3765}), .b ({signal_4568, signal_4273}), .c ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_163 ( .a ({signal_4570, signal_3764}), .b ({signal_4571, signal_4272}), .c ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_164 ( .a ({signal_4573, signal_3763}), .b ({signal_4574, signal_4271}), .c ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_165 ( .a ({signal_4576, signal_3762}), .b ({signal_4577, signal_4270}), .c ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_166 ( .a ({signal_4579, signal_3761}), .b ({signal_4580, signal_4269}), .c ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_167 ( .a ({signal_4582, signal_3860}), .b ({signal_4583, signal_4368}), .c ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_168 ( .a ({signal_4585, signal_3760}), .b ({signal_4586, signal_4268}), .c ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_169 ( .a ({signal_4588, signal_3759}), .b ({signal_4589, signal_4267}), .c ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_170 ( .a ({signal_4591, signal_3758}), .b ({signal_4592, signal_4266}), .c ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_171 ( .a ({signal_4594, signal_3757}), .b ({signal_4595, signal_4265}), .c ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_172 ( .a ({signal_4597, signal_3756}), .b ({signal_4598, signal_4264}), .c ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_173 ( .a ({signal_4600, signal_3755}), .b ({signal_4601, signal_4263}), .c ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_174 ( .a ({signal_4603, signal_3754}), .b ({signal_4604, signal_4262}), .c ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_175 ( .a ({signal_4606, signal_3753}), .b ({signal_4607, signal_4261}), .c ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_176 ( .a ({signal_4609, signal_3752}), .b ({signal_4610, signal_4260}), .c ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_177 ( .a ({signal_4612, signal_3751}), .b ({signal_4613, signal_4259}), .c ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_178 ( .a ({signal_4615, signal_3859}), .b ({signal_4616, signal_4367}), .c ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_179 ( .a ({signal_4618, signal_3750}), .b ({signal_4619, signal_4258}), .c ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_180 ( .a ({signal_4621, signal_3749}), .b ({signal_4622, signal_4257}), .c ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_181 ( .a ({signal_4624, signal_3748}), .b ({signal_4625, signal_4256}), .c ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_182 ( .a ({signal_4627, signal_3747}), .b ({signal_4628, signal_4255}), .c ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_183 ( .a ({signal_4630, signal_3746}), .b ({signal_4631, signal_4254}), .c ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_184 ( .a ({signal_4633, signal_3745}), .b ({signal_4634, signal_4253}), .c ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_185 ( .a ({signal_4636, signal_3744}), .b ({signal_4637, signal_4252}), .c ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_186 ( .a ({signal_4639, signal_3743}), .b ({signal_4640, signal_4251}), .c ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_187 ( .a ({signal_4642, signal_3858}), .b ({signal_4643, signal_4366}), .c ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_188 ( .a ({signal_4645, signal_3857}), .b ({signal_4646, signal_4365}), .c ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_189 ( .a ({signal_4648, signal_3856}), .b ({signal_4649, signal_4364}), .c ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_190 ( .a ({signal_4651, signal_3855}), .b ({signal_4652, signal_4363}), .c ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_191 ( .a ({signal_4654, signal_3854}), .b ({signal_4655, signal_4362}), .c ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_192 ( .a ({signal_4657, signal_3853}), .b ({signal_4658, signal_4361}), .c ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_193 ( .a ({signal_4660, signal_3852}), .b ({signal_4661, signal_4360}), .c ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_194 ( .a ({signal_4663, signal_3851}), .b ({signal_4664, signal_4359}), .c ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_195 ( .a ({signal_4666, signal_3869}), .b ({signal_4667, signal_4377}), .c ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_196 ( .a ({signal_4669, signal_3850}), .b ({signal_4670, signal_4358}), .c ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_197 ( .a ({signal_4672, signal_3849}), .b ({signal_4673, signal_4357}), .c ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_198 ( .a ({signal_4675, signal_3848}), .b ({signal_4676, signal_4356}), .c ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_199 ( .a ({signal_4678, signal_3847}), .b ({signal_4679, signal_4355}), .c ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_200 ( .a ({signal_4681, signal_3846}), .b ({signal_4682, signal_4354}), .c ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_201 ( .a ({signal_4684, signal_3845}), .b ({signal_4685, signal_4353}), .c ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_202 ( .a ({signal_4687, signal_3844}), .b ({signal_4688, signal_4352}), .c ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_203 ( .a ({signal_4690, signal_3843}), .b ({signal_4691, signal_4351}), .c ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_204 ( .a ({signal_4693, signal_3842}), .b ({signal_4694, signal_4350}), .c ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_205 ( .a ({signal_4696, signal_3841}), .b ({signal_4697, signal_4349}), .c ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_206 ( .a ({signal_4699, signal_3868}), .b ({signal_4700, signal_4376}), .c ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_207 ( .a ({signal_4702, signal_3840}), .b ({signal_4703, signal_4348}), .c ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_208 ( .a ({signal_4705, signal_3839}), .b ({signal_4706, signal_4347}), .c ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_209 ( .a ({signal_4708, signal_3838}), .b ({signal_4709, signal_4346}), .c ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_210 ( .a ({signal_4711, signal_3837}), .b ({signal_4712, signal_4345}), .c ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_211 ( .a ({signal_4714, signal_3836}), .b ({signal_4715, signal_4344}), .c ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_212 ( .a ({signal_4717, signal_3835}), .b ({signal_4718, signal_4343}), .c ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_213 ( .a ({signal_4720, signal_3834}), .b ({signal_4721, signal_4342}), .c ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_214 ( .a ({signal_4723, signal_3833}), .b ({signal_4724, signal_4341}), .c ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_215 ( .a ({signal_4726, signal_3832}), .b ({signal_4727, signal_4340}), .c ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_216 ( .a ({signal_4729, signal_3831}), .b ({signal_4730, signal_4339}), .c ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_217 ( .a ({signal_4732, signal_3867}), .b ({signal_4733, signal_4375}), .c ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_218 ( .a ({signal_4735, signal_3830}), .b ({signal_4736, signal_4338}), .c ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_219 ( .a ({signal_4738, signal_3829}), .b ({signal_4739, signal_4337}), .c ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_220 ( .a ({signal_4741, signal_3828}), .b ({signal_4742, signal_4336}), .c ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_221 ( .a ({signal_4744, signal_3827}), .b ({signal_4745, signal_4335}), .c ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_222 ( .a ({signal_4747, signal_3826}), .b ({signal_4748, signal_4334}), .c ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_223 ( .a ({signal_4750, signal_3825}), .b ({signal_4751, signal_4333}), .c ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_224 ( .a ({signal_4753, signal_3824}), .b ({signal_4754, signal_4332}), .c ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_225 ( .a ({signal_4756, signal_3823}), .b ({signal_4757, signal_4331}), .c ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_226 ( .a ({signal_4759, signal_3822}), .b ({signal_4760, signal_4330}), .c ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_227 ( .a ({signal_4762, signal_3821}), .b ({signal_4763, signal_4329}), .c ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_228 ( .a ({signal_4765, signal_3866}), .b ({signal_4766, signal_4374}), .c ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_229 ( .a ({signal_4768, signal_3820}), .b ({signal_4769, signal_4328}), .c ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_230 ( .a ({signal_4771, signal_3819}), .b ({signal_4772, signal_4327}), .c ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_231 ( .a ({signal_4774, signal_3818}), .b ({signal_4775, signal_4326}), .c ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_232 ( .a ({signal_4777, signal_3817}), .b ({signal_4778, signal_4325}), .c ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_233 ( .a ({signal_4780, signal_3816}), .b ({signal_4781, signal_4324}), .c ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_234 ( .a ({signal_4783, signal_3815}), .b ({signal_4784, signal_4323}), .c ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_235 ( .a ({signal_4786, signal_3814}), .b ({signal_4787, signal_4322}), .c ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_236 ( .a ({signal_4789, signal_3813}), .b ({signal_4790, signal_4321}), .c ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_237 ( .a ({signal_4792, signal_3812}), .b ({signal_4793, signal_4320}), .c ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_238 ( .a ({signal_4795, signal_3811}), .b ({signal_4796, signal_4319}), .c ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_239 ( .a ({signal_4798, signal_3865}), .b ({signal_4799, signal_4373}), .c ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_240 ( .a ({signal_4801, signal_3810}), .b ({signal_4802, signal_4318}), .c ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_241 ( .a ({signal_4804, signal_3809}), .b ({signal_4805, signal_4317}), .c ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_242 ( .a ({signal_4807, signal_3808}), .b ({signal_4808, signal_4316}), .c ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_243 ( .a ({signal_4810, signal_3807}), .b ({signal_4811, signal_4315}), .c ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_244 ( .a ({signal_4813, signal_3806}), .b ({signal_4814, signal_4314}), .c ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_245 ( .a ({signal_4816, signal_3805}), .b ({signal_4817, signal_4313}), .c ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_246 ( .a ({signal_4819, signal_3804}), .b ({signal_4820, signal_4312}), .c ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_247 ( .a ({signal_4822, signal_3803}), .b ({signal_4823, signal_4311}), .c ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_248 ( .a ({signal_4825, signal_3802}), .b ({signal_4826, signal_4310}), .c ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_249 ( .a ({signal_4828, signal_3801}), .b ({signal_4829, signal_4309}), .c ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_250 ( .a ({signal_4831, signal_3864}), .b ({signal_4832, signal_4372}), .c ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_251 ( .a ({signal_4834, signal_3800}), .b ({signal_4835, signal_4308}), .c ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_252 ( .a ({signal_4837, signal_3799}), .b ({signal_4838, signal_4307}), .c ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_253 ( .a ({signal_4840, signal_3798}), .b ({signal_4841, signal_4306}), .c ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_254 ( .a ({signal_4843, signal_3797}), .b ({signal_4844, signal_4305}), .c ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_255 ( .a ({signal_4846, signal_3796}), .b ({signal_4847, signal_4304}), .c ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_256 ( .a ({signal_4849, signal_3795}), .b ({signal_4850, signal_4303}), .c ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_257 ( .a ({signal_4852, signal_3794}), .b ({signal_4853, signal_4302}), .c ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_258 ( .a ({signal_4855, signal_3793}), .b ({signal_4856, signal_4301}), .c ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_259 ( .a ({signal_4858, signal_3792}), .b ({signal_4859, signal_4300}), .c ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_260 ( .a ({signal_4861, signal_3791}), .b ({signal_4862, signal_4299}), .c ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_261 ( .a ({signal_4864, signal_3863}), .b ({signal_4865, signal_4371}), .c ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_262 ( .a ({signal_4867, signal_3790}), .b ({signal_4868, signal_4298}), .c ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_263 ( .a ({signal_4870, signal_3789}), .b ({signal_4871, signal_4297}), .c ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_264 ( .a ({signal_4873, signal_3788}), .b ({signal_4874, signal_4296}), .c ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_265 ( .a ({signal_4876, signal_3787}), .b ({signal_4877, signal_4295}), .c ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_266 ( .a ({signal_4879, signal_3786}), .b ({signal_4880, signal_4294}), .c ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_267 ( .a ({signal_4882, signal_3785}), .b ({signal_4883, signal_4293}), .c ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_268 ( .a ({signal_4885, signal_3784}), .b ({signal_4886, signal_4292}), .c ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_269 ( .a ({signal_4888, signal_3783}), .b ({signal_4889, signal_4291}), .c ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_270 ( .a ({signal_4891, signal_3782}), .b ({signal_4892, signal_4290}), .c ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_271 ( .a ({signal_4894, signal_3781}), .b ({signal_4895, signal_4289}), .c ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_272 ( .a ({signal_4897, signal_3862}), .b ({signal_4898, signal_4370}), .c ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_273 ( .a ({signal_4900, signal_3780}), .b ({signal_4901, signal_4288}), .c ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_274 ( .a ({signal_4903, signal_3779}), .b ({signal_4904, signal_4287}), .c ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_275 ( .a ({signal_4906, signal_3778}), .b ({signal_4907, signal_4286}), .c ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_276 ( .a ({signal_4909, signal_3777}), .b ({signal_4910, signal_4285}), .c ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_277 ( .a ({signal_4912, signal_3776}), .b ({signal_4913, signal_4284}), .c ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_278 ( .a ({signal_4915, signal_3775}), .b ({signal_4916, signal_4283}), .c ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_279 ( .a ({signal_4918, signal_3774}), .b ({signal_4919, signal_4282}), .c ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_280 ( .a ({signal_4921, signal_3773}), .b ({signal_4922, signal_4281}), .c ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_281 ( .a ({signal_4924, signal_3772}), .b ({signal_4925, signal_4280}), .c ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_282 ( .a ({signal_4927, signal_3771}), .b ({signal_4928, signal_4279}), .c ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_283 ( .a ({signal_4930, signal_3861}), .b ({signal_4931, signal_4369}), .c ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    NAND2_X1 cell_284 ( .A1 (signal_4385), .A2 (signal_414), .ZN (signal_415) ) ;
    NOR2_X1 cell_285 ( .A1 (signal_4388), .A2 (signal_415), .ZN (done) ) ;
    INV_X1 cell_286 ( .A (signal_416), .ZN (signal_417) ) ;
    NAND2_X1 cell_287 ( .A1 (signal_4386), .A2 (signal_4387), .ZN (signal_419) ) ;
    NOR2_X1 cell_288 ( .A1 (signal_417), .A2 (signal_419), .ZN (signal_393) ) ;
    INV_X1 cell_289 ( .A (signal_418), .ZN (signal_420) ) ;
    NOR2_X1 cell_290 ( .A1 (signal_420), .A2 (signal_419), .ZN (signal_394) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_679 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_4933, signal_792}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_807 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_4934, signal_912}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_935 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_4935, signal_1032}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1063 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_4936, signal_1152}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1191 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_4937, signal_1272}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1319 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_4938, signal_1392}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1447 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_4939, signal_1512}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1575 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_4940, signal_1632}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1703 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_4941, signal_1752}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1831 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_4942, signal_1872}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1959 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_4943, signal_1992}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_2087 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_4944, signal_2112}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_2215 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_4945, signal_2232}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_2343 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_4946, signal_2352}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_2471 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_4947, signal_2472}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_2599 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_4948, signal_2592}) ) ;
    INV_X1 cell_4187 ( .A (signal_3597), .ZN (signal_3607) ) ;
    MUX2_X1 cell_4188 ( .S (signal_3609), .A (signal_3598), .B (signal_3599), .Z (signal_3597) ) ;
    NOR2_X1 cell_4189 ( .A1 (reset), .A2 (signal_3600), .ZN (signal_3610) ) ;
    XNOR2_X1 cell_4190 ( .A (signal_4388), .B (signal_4387), .ZN (signal_3600) ) ;
    MUX2_X1 cell_4191 ( .S (signal_4385), .A (signal_3601), .B (signal_3602), .Z (signal_3608) ) ;
    NAND2_X1 cell_4192 ( .A1 (signal_3598), .A2 (signal_3603), .ZN (signal_3602) ) ;
    NAND2_X1 cell_4193 ( .A1 (signal_3609), .A2 (signal_3606), .ZN (signal_3603) ) ;
    NOR2_X1 cell_4194 ( .A1 (signal_3604), .A2 (signal_3612), .ZN (signal_3598) ) ;
    NOR2_X1 cell_4195 ( .A1 (signal_4387), .A2 (reset), .ZN (signal_3604) ) ;
    NOR2_X1 cell_4196 ( .A1 (signal_3609), .A2 (signal_3599), .ZN (signal_3601) ) ;
    NAND2_X1 cell_4197 ( .A1 (signal_4387), .A2 (signal_3605), .ZN (signal_3599) ) ;
    NOR2_X1 cell_4198 ( .A1 (reset), .A2 (signal_3611), .ZN (signal_3605) ) ;
    NOR2_X1 cell_4199 ( .A1 (reset), .A2 (signal_4388), .ZN (signal_3612) ) ;
    INV_X1 cell_4200 ( .A (reset), .ZN (signal_3606) ) ;
    INV_X1 cell_4201 ( .A (signal_4388), .ZN (signal_3611) ) ;
    INV_X1 cell_4205 ( .A (signal_4386), .ZN (signal_3609) ) ;
    ClockGatingController #(3) cell_4210 ( .clk (clk), .rst (reset), .GatedClk (signal_6181), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_28 ( .s (signal_402), .b ({signal_5012, signal_3994}), .a ({signal_5364, signal_4122}), .c ({signal_5394, signal_3742}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_29 ( .s (signal_402), .b ({signal_5150, signal_4415}), .a ({signal_5039, signal_4022}), .c ({signal_5237, signal_3642}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_30 ( .s (signal_402), .b ({signal_5149, signal_4414}), .a ({signal_5038, signal_4021}), .c ({signal_5238, signal_3641}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_31 ( .s (signal_402), .b ({signal_5148, signal_4413}), .a ({signal_5037, signal_4020}), .c ({signal_5239, signal_3640}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_32 ( .s (signal_402), .b ({signal_5152, signal_4420}), .a ({signal_5036, signal_4019}), .c ({signal_5240, signal_3639}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_33 ( .s (signal_402), .b ({signal_4973, signal_3890}), .a ({signal_5035, signal_4018}), .c ({signal_5241, signal_3638}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_34 ( .s (signal_402), .b ({signal_5146, signal_4410}), .a ({signal_5357, signal_4017}), .c ({signal_5395, signal_3637}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_35 ( .s (signal_402), .b ({signal_4972, signal_3888}), .a ({signal_5034, signal_4016}), .c ({signal_5242, signal_3636}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_36 ( .s (signal_396), .b ({signal_4971, signal_3887}), .a ({signal_5033, signal_4015}), .c ({signal_5243, signal_3635}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_37 ( .s (signal_397), .b ({signal_5145, signal_4407}), .a ({signal_5032, signal_4014}), .c ({signal_5244, signal_3634}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_38 ( .s (signal_398), .b ({signal_5144, signal_4406}), .a ({signal_5031, signal_4013}), .c ({signal_5245, signal_3633}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_39 ( .s (signal_399), .b ({signal_5008, signal_3984}), .a ({signal_5124, signal_4112}), .c ({signal_5246, signal_3732}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_40 ( .s (signal_400), .b ({signal_5143, signal_4405}), .a ({signal_5030, signal_4012}), .c ({signal_5247, signal_3632}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_41 ( .s (signal_401), .b ({signal_5147, signal_4412}), .a ({signal_5029, signal_4011}), .c ({signal_5248, signal_3631}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_42 ( .s (signal_400), .b ({signal_4970, signal_3882}), .a ({signal_5028, signal_4010}), .c ({signal_5249, signal_3630}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_43 ( .s (signal_399), .b ({signal_5141, signal_4402}), .a ({signal_5027, signal_4009}), .c ({signal_5250, signal_3629}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_44 ( .s (signal_399), .b ({signal_4969, signal_3880}), .a ({signal_5026, signal_4008}), .c ({signal_5251, signal_3628}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_45 ( .s (signal_396), .b ({signal_4968, signal_3879}), .a ({signal_5025, signal_4007}), .c ({signal_5252, signal_3627}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_46 ( .s (signal_397), .b ({signal_5140, signal_4399}), .a ({signal_5024, signal_4006}), .c ({signal_5253, signal_3626}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_47 ( .s (signal_398), .b ({signal_5139, signal_4398}), .a ({signal_5023, signal_4005}), .c ({signal_5254, signal_3625}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_48 ( .s (signal_400), .b ({signal_5138, signal_4397}), .a ({signal_5022, signal_4004}), .c ({signal_5255, signal_3624}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_49 ( .s (signal_401), .b ({signal_5142, signal_4404}), .a ({signal_5021, signal_4003}), .c ({signal_5256, signal_3623}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_50 ( .s (signal_401), .b ({signal_5007, signal_3983}), .a ({signal_5123, signal_4111}), .c ({signal_5257, signal_3731}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_51 ( .s (signal_400), .b ({signal_4967, signal_3874}), .a ({signal_5020, signal_4002}), .c ({signal_5258, signal_3622}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_52 ( .s (signal_399), .b ({signal_5136, signal_4394}), .a ({signal_5019, signal_4001}), .c ({signal_5259, signal_3621}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_53 ( .s (signal_400), .b ({signal_4966, signal_3872}), .a ({signal_5018, signal_4000}), .c ({signal_5260, signal_3620}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_54 ( .s (signal_401), .b ({signal_4965, signal_3871}), .a ({signal_5017, signal_3999}), .c ({signal_5261, signal_3619}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_55 ( .s (signal_397), .b ({signal_5135, signal_4391}), .a ({signal_5016, signal_3998}), .c ({signal_5262, signal_3618}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_56 ( .s (signal_401), .b ({signal_5134, signal_4390}), .a ({signal_5015, signal_3997}), .c ({signal_5263, signal_3617}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_57 ( .s (signal_397), .b ({signal_5133, signal_4389}), .a ({signal_5014, signal_3996}), .c ({signal_5264, signal_3616}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_58 ( .s (signal_398), .b ({signal_5137, signal_4396}), .a ({signal_5013, signal_3995}), .c ({signal_5265, signal_3615}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_59 ( .s (signal_396), .b ({signal_5205, signal_4503}), .a ({signal_5122, signal_4110}), .c ({signal_5266, signal_3730}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_60 ( .s (signal_398), .b ({signal_5204, signal_4502}), .a ({signal_5121, signal_4109}), .c ({signal_5267, signal_3729}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_61 ( .s (signal_397), .b ({signal_5203, signal_4501}), .a ({signal_5120, signal_4108}), .c ({signal_5268, signal_3728}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_62 ( .s (signal_398), .b ({signal_5207, signal_4508}), .a ({signal_5119, signal_4107}), .c ({signal_5269, signal_3727}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_63 ( .s (signal_396), .b ({signal_5006, signal_3978}), .a ({signal_5118, signal_4106}), .c ({signal_5270, signal_3726}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_64 ( .s (signal_399), .b ({signal_5201, signal_4498}), .a ({signal_5117, signal_4105}), .c ({signal_5271, signal_3725}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_65 ( .s (signal_400), .b ({signal_5005, signal_3976}), .a ({signal_5116, signal_4104}), .c ({signal_5272, signal_3724}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_66 ( .s (signal_401), .b ({signal_5004, signal_3975}), .a ({signal_5115, signal_4103}), .c ({signal_5273, signal_3723}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_67 ( .s (signal_399), .b ({signal_5211, signal_4514}), .a ({signal_5132, signal_4121}), .c ({signal_5274, signal_3741}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_68 ( .s (signal_400), .b ({signal_5200, signal_4495}), .a ({signal_5114, signal_4102}), .c ({signal_5275, signal_3722}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_69 ( .s (signal_397), .b ({signal_5199, signal_4494}), .a ({signal_5113, signal_4101}), .c ({signal_5276, signal_3721}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_70 ( .s (signal_398), .b ({signal_5198, signal_4493}), .a ({signal_5112, signal_4100}), .c ({signal_5277, signal_3720}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_71 ( .s (signal_396), .b ({signal_5202, signal_4500}), .a ({signal_5111, signal_4099}), .c ({signal_5278, signal_3719}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_72 ( .s (signal_401), .b ({signal_5003, signal_3970}), .a ({signal_5110, signal_4098}), .c ({signal_5279, signal_3718}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_73 ( .s (signal_399), .b ({signal_5196, signal_4490}), .a ({signal_5109, signal_4097}), .c ({signal_5280, signal_3717}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_74 ( .s (signal_397), .b ({signal_5002, signal_3968}), .a ({signal_5108, signal_4096}), .c ({signal_5281, signal_3716}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_75 ( .s (signal_398), .b ({signal_5001, signal_3967}), .a ({signal_5107, signal_4095}), .c ({signal_5282, signal_3715}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_76 ( .s (signal_396), .b ({signal_5195, signal_4487}), .a ({signal_5106, signal_4094}), .c ({signal_5283, signal_3714}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_77 ( .s (signal_400), .b ({signal_5194, signal_4486}), .a ({signal_5105, signal_4093}), .c ({signal_5284, signal_3713}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_78 ( .s (signal_396), .b ({signal_5011, signal_3992}), .a ({signal_5131, signal_4120}), .c ({signal_5285, signal_3740}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_79 ( .s (signal_401), .b ({signal_5193, signal_4485}), .a ({signal_5104, signal_4092}), .c ({signal_5286, signal_3712}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_80 ( .s (signal_399), .b ({signal_5197, signal_4492}), .a ({signal_5103, signal_4091}), .c ({signal_5287, signal_3711}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_81 ( .s (signal_397), .b ({signal_5000, signal_3962}), .a ({signal_5362, signal_4090}), .c ({signal_5396, signal_3710}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_82 ( .s (signal_398), .b ({signal_5191, signal_4482}), .a ({signal_5102, signal_4089}), .c ({signal_5288, signal_3709}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_83 ( .s (signal_396), .b ({signal_4999, signal_3960}), .a ({signal_5101, signal_4088}), .c ({signal_5289, signal_3708}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_84 ( .s (signal_401), .b ({signal_4998, signal_3959}), .a ({signal_5100, signal_4087}), .c ({signal_5290, signal_3707}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_85 ( .s (signal_401), .b ({signal_5190, signal_4479}), .a ({signal_5099, signal_4086}), .c ({signal_5291, signal_3706}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_86 ( .s (signal_401), .b ({signal_5189, signal_4478}), .a ({signal_5098, signal_4085}), .c ({signal_5292, signal_3705}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_87 ( .s (signal_401), .b ({signal_5188, signal_4477}), .a ({signal_5097, signal_4084}), .c ({signal_5293, signal_3704}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_88 ( .s (signal_401), .b ({signal_5192, signal_4484}), .a ({signal_5096, signal_4083}), .c ({signal_5294, signal_3703}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_89 ( .s (signal_401), .b ({signal_5010, signal_3991}), .a ({signal_5130, signal_4119}), .c ({signal_5295, signal_3739}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_90 ( .s (signal_401), .b ({signal_4997, signal_3954}), .a ({signal_5095, signal_4082}), .c ({signal_5296, signal_3702}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_91 ( .s (signal_401), .b ({signal_5186, signal_4474}), .a ({signal_5361, signal_4081}), .c ({signal_5397, signal_3701}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_92 ( .s (signal_401), .b ({signal_4996, signal_3952}), .a ({signal_5094, signal_4080}), .c ({signal_5297, signal_3700}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_93 ( .s (signal_401), .b ({signal_4995, signal_3951}), .a ({signal_5093, signal_4079}), .c ({signal_5298, signal_3699}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_94 ( .s (signal_401), .b ({signal_5185, signal_4471}), .a ({signal_5092, signal_4078}), .c ({signal_5299, signal_3698}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_95 ( .s (signal_401), .b ({signal_5184, signal_4470}), .a ({signal_5091, signal_4077}), .c ({signal_5300, signal_3697}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_96 ( .s (signal_400), .b ({signal_5183, signal_4469}), .a ({signal_5090, signal_4076}), .c ({signal_5301, signal_3696}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_97 ( .s (signal_400), .b ({signal_5187, signal_4476}), .a ({signal_5089, signal_4075}), .c ({signal_5302, signal_3695}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_98 ( .s (signal_400), .b ({signal_4994, signal_3946}), .a ({signal_5088, signal_4074}), .c ({signal_5303, signal_3694}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_99 ( .s (signal_400), .b ({signal_5181, signal_4466}), .a ({signal_5087, signal_4073}), .c ({signal_5304, signal_3693}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_100 ( .s (signal_400), .b ({signal_5210, signal_4511}), .a ({signal_5129, signal_4118}), .c ({signal_5305, signal_3738}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_101 ( .s (signal_400), .b ({signal_4993, signal_3944}), .a ({signal_5086, signal_4072}), .c ({signal_5306, signal_3692}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_102 ( .s (signal_400), .b ({signal_4992, signal_3943}), .a ({signal_5085, signal_4071}), .c ({signal_5307, signal_3691}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_103 ( .s (signal_400), .b ({signal_5180, signal_4463}), .a ({signal_5084, signal_4070}), .c ({signal_5308, signal_3690}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_104 ( .s (signal_400), .b ({signal_5179, signal_4462}), .a ({signal_5083, signal_4069}), .c ({signal_5309, signal_3689}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_105 ( .s (signal_400), .b ({signal_5178, signal_4461}), .a ({signal_5082, signal_4068}), .c ({signal_5310, signal_3688}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_106 ( .s (signal_400), .b ({signal_5182, signal_4468}), .a ({signal_5081, signal_4067}), .c ({signal_5311, signal_3687}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_107 ( .s (signal_400), .b ({signal_4991, signal_3938}), .a ({signal_5080, signal_4066}), .c ({signal_5312, signal_3686}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_108 ( .s (signal_399), .b ({signal_5176, signal_4458}), .a ({signal_5079, signal_4065}), .c ({signal_5313, signal_3685}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_109 ( .s (signal_399), .b ({signal_4990, signal_3936}), .a ({signal_5078, signal_4064}), .c ({signal_5314, signal_3684}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_110 ( .s (signal_399), .b ({signal_4989, signal_3935}), .a ({signal_5077, signal_4063}), .c ({signal_5315, signal_3683}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_111 ( .s (signal_399), .b ({signal_5209, signal_4510}), .a ({signal_5128, signal_4117}), .c ({signal_5316, signal_3737}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_112 ( .s (signal_399), .b ({signal_5175, signal_4455}), .a ({signal_5076, signal_4062}), .c ({signal_5317, signal_3682}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_113 ( .s (signal_399), .b ({signal_5174, signal_4454}), .a ({signal_5075, signal_4061}), .c ({signal_5318, signal_3681}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_114 ( .s (signal_399), .b ({signal_5173, signal_4453}), .a ({signal_5074, signal_4060}), .c ({signal_5319, signal_3680}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_115 ( .s (signal_399), .b ({signal_5177, signal_4460}), .a ({signal_5073, signal_4059}), .c ({signal_5320, signal_3679}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_116 ( .s (signal_399), .b ({signal_4988, signal_3930}), .a ({signal_5360, signal_4058}), .c ({signal_5398, signal_3678}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_117 ( .s (signal_399), .b ({signal_5171, signal_4450}), .a ({signal_5072, signal_4057}), .c ({signal_5321, signal_3677}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_118 ( .s (signal_399), .b ({signal_4987, signal_3928}), .a ({signal_5071, signal_4056}), .c ({signal_5322, signal_3676}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_119 ( .s (signal_399), .b ({signal_4986, signal_3927}), .a ({signal_5070, signal_4055}), .c ({signal_5323, signal_3675}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_120 ( .s (signal_398), .b ({signal_5170, signal_4447}), .a ({signal_5069, signal_4054}), .c ({signal_5324, signal_3674}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_121 ( .s (signal_398), .b ({signal_5169, signal_4446}), .a ({signal_5068, signal_4053}), .c ({signal_5325, signal_3673}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_122 ( .s (signal_398), .b ({signal_5208, signal_4509}), .a ({signal_5127, signal_4116}), .c ({signal_5326, signal_3736}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_123 ( .s (signal_398), .b ({signal_5168, signal_4445}), .a ({signal_5067, signal_4052}), .c ({signal_5327, signal_3672}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_124 ( .s (signal_398), .b ({signal_5172, signal_4452}), .a ({signal_5066, signal_4051}), .c ({signal_5328, signal_3671}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_125 ( .s (signal_398), .b ({signal_4985, signal_3922}), .a ({signal_5065, signal_4050}), .c ({signal_5329, signal_3670}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_126 ( .s (signal_398), .b ({signal_5166, signal_4442}), .a ({signal_5359, signal_4049}), .c ({signal_5399, signal_3669}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_127 ( .s (signal_398), .b ({signal_4984, signal_3920}), .a ({signal_5064, signal_4048}), .c ({signal_5330, signal_3668}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_128 ( .s (signal_398), .b ({signal_4983, signal_3919}), .a ({signal_5063, signal_4047}), .c ({signal_5331, signal_3667}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_129 ( .s (signal_398), .b ({signal_5165, signal_4439}), .a ({signal_5062, signal_4046}), .c ({signal_5332, signal_3666}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_130 ( .s (signal_398), .b ({signal_5164, signal_4438}), .a ({signal_5061, signal_4045}), .c ({signal_5333, signal_3665}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_131 ( .s (signal_398), .b ({signal_5163, signal_4437}), .a ({signal_5060, signal_4044}), .c ({signal_5334, signal_3664}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_132 ( .s (signal_397), .b ({signal_5167, signal_4444}), .a ({signal_5059, signal_4043}), .c ({signal_5335, signal_3663}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_133 ( .s (signal_397), .b ({signal_5212, signal_4516}), .a ({signal_5126, signal_4115}), .c ({signal_5336, signal_3735}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_134 ( .s (signal_397), .b ({signal_4982, signal_3914}), .a ({signal_5058, signal_4042}), .c ({signal_5337, signal_3662}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_135 ( .s (signal_397), .b ({signal_5161, signal_4434}), .a ({signal_5057, signal_4041}), .c ({signal_5338, signal_3661}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_136 ( .s (signal_397), .b ({signal_4981, signal_3912}), .a ({signal_5056, signal_4040}), .c ({signal_5339, signal_3660}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_137 ( .s (signal_397), .b ({signal_4980, signal_3911}), .a ({signal_5055, signal_4039}), .c ({signal_5340, signal_3659}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_138 ( .s (signal_397), .b ({signal_5160, signal_4431}), .a ({signal_5054, signal_4038}), .c ({signal_5341, signal_3658}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_139 ( .s (signal_397), .b ({signal_5159, signal_4430}), .a ({signal_5053, signal_4037}), .c ({signal_5342, signal_3657}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_140 ( .s (signal_397), .b ({signal_5158, signal_4429}), .a ({signal_5052, signal_4036}), .c ({signal_5343, signal_3656}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_141 ( .s (signal_397), .b ({signal_5162, signal_4436}), .a ({signal_5051, signal_4035}), .c ({signal_5344, signal_3655}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_142 ( .s (signal_397), .b ({signal_4979, signal_3906}), .a ({signal_5050, signal_4034}), .c ({signal_5345, signal_3654}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_143 ( .s (signal_397), .b ({signal_5156, signal_4426}), .a ({signal_5049, signal_4033}), .c ({signal_5346, signal_3653}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_144 ( .s (signal_396), .b ({signal_5009, signal_3986}), .a ({signal_5125, signal_4114}), .c ({signal_5347, signal_3734}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_145 ( .s (signal_396), .b ({signal_4978, signal_3904}), .a ({signal_5048, signal_4032}), .c ({signal_5348, signal_3652}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_146 ( .s (signal_396), .b ({signal_4977, signal_3903}), .a ({signal_5047, signal_4031}), .c ({signal_5349, signal_3651}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_147 ( .s (signal_396), .b ({signal_5155, signal_4423}), .a ({signal_5046, signal_4030}), .c ({signal_5350, signal_3650}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_148 ( .s (signal_396), .b ({signal_5154, signal_4422}), .a ({signal_5045, signal_4029}), .c ({signal_5351, signal_3649}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_149 ( .s (signal_396), .b ({signal_5153, signal_4421}), .a ({signal_5044, signal_4028}), .c ({signal_5352, signal_3648}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_150 ( .s (signal_396), .b ({signal_5157, signal_4428}), .a ({signal_5043, signal_4027}), .c ({signal_5353, signal_3647}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_151 ( .s (signal_396), .b ({signal_4976, signal_3898}), .a ({signal_5358, signal_4026}), .c ({signal_5400, signal_3646}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_152 ( .s (signal_396), .b ({signal_5151, signal_4418}), .a ({signal_5042, signal_4025}), .c ({signal_5354, signal_3645}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_153 ( .s (signal_396), .b ({signal_4975, signal_3896}), .a ({signal_5041, signal_4024}), .c ({signal_5355, signal_3644}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_154 ( .s (signal_396), .b ({signal_4974, signal_3895}), .a ({signal_5040, signal_4023}), .c ({signal_5356, signal_3643}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_155 ( .s (signal_396), .b ({signal_5206, signal_4506}), .a ({signal_5363, signal_4113}), .c ({signal_5401, signal_3733}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_291 ( .s (reset), .b ({signal_5394, signal_3742}), .a ({plaintext_s1[0], plaintext_s0[0]}), .c ({signal_5723, signal_421}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_294 ( .s (reset), .b ({signal_5274, signal_3741}), .a ({plaintext_s1[1], plaintext_s0[1]}), .c ({signal_5403, signal_423}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_297 ( .s (reset), .b ({signal_5285, signal_3740}), .a ({plaintext_s1[2], plaintext_s0[2]}), .c ({signal_5405, signal_425}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_300 ( .s (reset), .b ({signal_5295, signal_3739}), .a ({plaintext_s1[3], plaintext_s0[3]}), .c ({signal_5407, signal_427}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_303 ( .s (reset), .b ({signal_5305, signal_3738}), .a ({plaintext_s1[4], plaintext_s0[4]}), .c ({signal_5409, signal_429}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_306 ( .s (reset), .b ({signal_5316, signal_3737}), .a ({plaintext_s1[5], plaintext_s0[5]}), .c ({signal_5411, signal_431}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_309 ( .s (reset), .b ({signal_5326, signal_3736}), .a ({plaintext_s1[6], plaintext_s0[6]}), .c ({signal_5413, signal_433}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_312 ( .s (reset), .b ({signal_5336, signal_3735}), .a ({plaintext_s1[7], plaintext_s0[7]}), .c ({signal_5415, signal_435}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_315 ( .s (reset), .b ({signal_5347, signal_3734}), .a ({plaintext_s1[8], plaintext_s0[8]}), .c ({signal_5417, signal_437}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_318 ( .s (reset), .b ({signal_5401, signal_3733}), .a ({plaintext_s1[9], plaintext_s0[9]}), .c ({signal_5725, signal_439}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_321 ( .s (reset), .b ({signal_5246, signal_3732}), .a ({plaintext_s1[10], plaintext_s0[10]}), .c ({signal_5419, signal_441}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_324 ( .s (reset), .b ({signal_5257, signal_3731}), .a ({plaintext_s1[11], plaintext_s0[11]}), .c ({signal_5421, signal_443}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_327 ( .s (reset), .b ({signal_5266, signal_3730}), .a ({plaintext_s1[12], plaintext_s0[12]}), .c ({signal_5423, signal_445}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_330 ( .s (reset), .b ({signal_5267, signal_3729}), .a ({plaintext_s1[13], plaintext_s0[13]}), .c ({signal_5425, signal_447}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_333 ( .s (reset), .b ({signal_5268, signal_3728}), .a ({plaintext_s1[14], plaintext_s0[14]}), .c ({signal_5427, signal_449}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_336 ( .s (reset), .b ({signal_5269, signal_3727}), .a ({plaintext_s1[15], plaintext_s0[15]}), .c ({signal_5429, signal_451}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_339 ( .s (reset), .b ({signal_5270, signal_3726}), .a ({plaintext_s1[16], plaintext_s0[16]}), .c ({signal_5431, signal_453}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_342 ( .s (reset), .b ({signal_5271, signal_3725}), .a ({plaintext_s1[17], plaintext_s0[17]}), .c ({signal_5433, signal_455}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_345 ( .s (reset), .b ({signal_5272, signal_3724}), .a ({plaintext_s1[18], plaintext_s0[18]}), .c ({signal_5435, signal_457}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_348 ( .s (reset), .b ({signal_5273, signal_3723}), .a ({plaintext_s1[19], plaintext_s0[19]}), .c ({signal_5437, signal_459}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_351 ( .s (reset), .b ({signal_5275, signal_3722}), .a ({plaintext_s1[20], plaintext_s0[20]}), .c ({signal_5439, signal_461}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_354 ( .s (reset), .b ({signal_5276, signal_3721}), .a ({plaintext_s1[21], plaintext_s0[21]}), .c ({signal_5441, signal_463}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_357 ( .s (reset), .b ({signal_5277, signal_3720}), .a ({plaintext_s1[22], plaintext_s0[22]}), .c ({signal_5443, signal_465}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_360 ( .s (reset), .b ({signal_5278, signal_3719}), .a ({plaintext_s1[23], plaintext_s0[23]}), .c ({signal_5445, signal_467}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_363 ( .s (reset), .b ({signal_5279, signal_3718}), .a ({plaintext_s1[24], plaintext_s0[24]}), .c ({signal_5447, signal_469}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_366 ( .s (reset), .b ({signal_5280, signal_3717}), .a ({plaintext_s1[25], plaintext_s0[25]}), .c ({signal_5449, signal_471}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_369 ( .s (reset), .b ({signal_5281, signal_3716}), .a ({plaintext_s1[26], plaintext_s0[26]}), .c ({signal_5451, signal_473}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_372 ( .s (reset), .b ({signal_5282, signal_3715}), .a ({plaintext_s1[27], plaintext_s0[27]}), .c ({signal_5453, signal_475}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_375 ( .s (reset), .b ({signal_5283, signal_3714}), .a ({plaintext_s1[28], plaintext_s0[28]}), .c ({signal_5455, signal_477}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_378 ( .s (reset), .b ({signal_5284, signal_3713}), .a ({plaintext_s1[29], plaintext_s0[29]}), .c ({signal_5457, signal_479}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_381 ( .s (reset), .b ({signal_5286, signal_3712}), .a ({plaintext_s1[30], plaintext_s0[30]}), .c ({signal_5459, signal_481}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_384 ( .s (reset), .b ({signal_5287, signal_3711}), .a ({plaintext_s1[31], plaintext_s0[31]}), .c ({signal_5461, signal_483}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_387 ( .s (reset), .b ({signal_5396, signal_3710}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({signal_5727, signal_485}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_390 ( .s (reset), .b ({signal_5288, signal_3709}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({signal_5463, signal_487}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_393 ( .s (reset), .b ({signal_5289, signal_3708}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({signal_5465, signal_489}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_396 ( .s (reset), .b ({signal_5290, signal_3707}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({signal_5467, signal_491}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_399 ( .s (reset), .b ({signal_5291, signal_3706}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({signal_5469, signal_493}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_402 ( .s (reset), .b ({signal_5292, signal_3705}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({signal_5471, signal_495}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_405 ( .s (reset), .b ({signal_5293, signal_3704}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({signal_5473, signal_497}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_408 ( .s (reset), .b ({signal_5294, signal_3703}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({signal_5475, signal_499}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_411 ( .s (reset), .b ({signal_5296, signal_3702}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({signal_5477, signal_501}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_414 ( .s (reset), .b ({signal_5397, signal_3701}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({signal_5729, signal_503}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_417 ( .s (reset), .b ({signal_5297, signal_3700}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({signal_5479, signal_505}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_420 ( .s (reset), .b ({signal_5298, signal_3699}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({signal_5481, signal_507}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_423 ( .s (reset), .b ({signal_5299, signal_3698}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({signal_5483, signal_509}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_426 ( .s (reset), .b ({signal_5300, signal_3697}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({signal_5485, signal_511}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_429 ( .s (reset), .b ({signal_5301, signal_3696}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({signal_5487, signal_513}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_432 ( .s (reset), .b ({signal_5302, signal_3695}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({signal_5489, signal_515}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_435 ( .s (reset), .b ({signal_5303, signal_3694}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({signal_5491, signal_517}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_438 ( .s (reset), .b ({signal_5304, signal_3693}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({signal_5493, signal_519}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_441 ( .s (reset), .b ({signal_5306, signal_3692}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({signal_5495, signal_521}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_444 ( .s (reset), .b ({signal_5307, signal_3691}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({signal_5497, signal_523}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_447 ( .s (reset), .b ({signal_5308, signal_3690}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({signal_5499, signal_525}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_450 ( .s (reset), .b ({signal_5309, signal_3689}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({signal_5501, signal_527}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_453 ( .s (reset), .b ({signal_5310, signal_3688}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({signal_5503, signal_529}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_456 ( .s (reset), .b ({signal_5311, signal_3687}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({signal_5505, signal_531}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_459 ( .s (reset), .b ({signal_5312, signal_3686}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({signal_5507, signal_533}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_462 ( .s (reset), .b ({signal_5313, signal_3685}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({signal_5509, signal_535}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_465 ( .s (reset), .b ({signal_5314, signal_3684}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({signal_5511, signal_537}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_468 ( .s (reset), .b ({signal_5315, signal_3683}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({signal_5513, signal_539}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_471 ( .s (reset), .b ({signal_5317, signal_3682}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({signal_5515, signal_541}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_474 ( .s (reset), .b ({signal_5318, signal_3681}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({signal_5517, signal_543}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_477 ( .s (reset), .b ({signal_5319, signal_3680}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({signal_5519, signal_545}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_480 ( .s (reset), .b ({signal_5320, signal_3679}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({signal_5521, signal_547}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_483 ( .s (reset), .b ({signal_5398, signal_3678}), .a ({plaintext_s1[64], plaintext_s0[64]}), .c ({signal_5731, signal_549}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_486 ( .s (reset), .b ({signal_5321, signal_3677}), .a ({plaintext_s1[65], plaintext_s0[65]}), .c ({signal_5523, signal_551}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_489 ( .s (reset), .b ({signal_5322, signal_3676}), .a ({plaintext_s1[66], plaintext_s0[66]}), .c ({signal_5525, signal_553}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_492 ( .s (reset), .b ({signal_5323, signal_3675}), .a ({plaintext_s1[67], plaintext_s0[67]}), .c ({signal_5527, signal_555}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_495 ( .s (reset), .b ({signal_5324, signal_3674}), .a ({plaintext_s1[68], plaintext_s0[68]}), .c ({signal_5529, signal_557}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_498 ( .s (reset), .b ({signal_5325, signal_3673}), .a ({plaintext_s1[69], plaintext_s0[69]}), .c ({signal_5531, signal_559}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_501 ( .s (reset), .b ({signal_5327, signal_3672}), .a ({plaintext_s1[70], plaintext_s0[70]}), .c ({signal_5533, signal_561}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_504 ( .s (reset), .b ({signal_5328, signal_3671}), .a ({plaintext_s1[71], plaintext_s0[71]}), .c ({signal_5535, signal_563}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_507 ( .s (reset), .b ({signal_5329, signal_3670}), .a ({plaintext_s1[72], plaintext_s0[72]}), .c ({signal_5537, signal_565}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_510 ( .s (reset), .b ({signal_5399, signal_3669}), .a ({plaintext_s1[73], plaintext_s0[73]}), .c ({signal_5733, signal_567}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_513 ( .s (reset), .b ({signal_5330, signal_3668}), .a ({plaintext_s1[74], plaintext_s0[74]}), .c ({signal_5539, signal_569}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_516 ( .s (reset), .b ({signal_5331, signal_3667}), .a ({plaintext_s1[75], plaintext_s0[75]}), .c ({signal_5541, signal_571}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_519 ( .s (reset), .b ({signal_5332, signal_3666}), .a ({plaintext_s1[76], plaintext_s0[76]}), .c ({signal_5543, signal_573}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_522 ( .s (reset), .b ({signal_5333, signal_3665}), .a ({plaintext_s1[77], plaintext_s0[77]}), .c ({signal_5545, signal_575}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_525 ( .s (reset), .b ({signal_5334, signal_3664}), .a ({plaintext_s1[78], plaintext_s0[78]}), .c ({signal_5547, signal_577}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_528 ( .s (reset), .b ({signal_5335, signal_3663}), .a ({plaintext_s1[79], plaintext_s0[79]}), .c ({signal_5549, signal_579}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_531 ( .s (reset), .b ({signal_5337, signal_3662}), .a ({plaintext_s1[80], plaintext_s0[80]}), .c ({signal_5551, signal_581}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_534 ( .s (reset), .b ({signal_5338, signal_3661}), .a ({plaintext_s1[81], plaintext_s0[81]}), .c ({signal_5553, signal_583}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_537 ( .s (reset), .b ({signal_5339, signal_3660}), .a ({plaintext_s1[82], plaintext_s0[82]}), .c ({signal_5555, signal_585}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_540 ( .s (reset), .b ({signal_5340, signal_3659}), .a ({plaintext_s1[83], plaintext_s0[83]}), .c ({signal_5557, signal_587}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_543 ( .s (reset), .b ({signal_5341, signal_3658}), .a ({plaintext_s1[84], plaintext_s0[84]}), .c ({signal_5559, signal_589}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_546 ( .s (reset), .b ({signal_5342, signal_3657}), .a ({plaintext_s1[85], plaintext_s0[85]}), .c ({signal_5561, signal_591}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_549 ( .s (reset), .b ({signal_5343, signal_3656}), .a ({plaintext_s1[86], plaintext_s0[86]}), .c ({signal_5563, signal_593}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_552 ( .s (reset), .b ({signal_5344, signal_3655}), .a ({plaintext_s1[87], plaintext_s0[87]}), .c ({signal_5565, signal_595}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_555 ( .s (reset), .b ({signal_5345, signal_3654}), .a ({plaintext_s1[88], plaintext_s0[88]}), .c ({signal_5567, signal_597}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_558 ( .s (reset), .b ({signal_5346, signal_3653}), .a ({plaintext_s1[89], plaintext_s0[89]}), .c ({signal_5569, signal_599}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_561 ( .s (reset), .b ({signal_5348, signal_3652}), .a ({plaintext_s1[90], plaintext_s0[90]}), .c ({signal_5571, signal_601}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_564 ( .s (reset), .b ({signal_5349, signal_3651}), .a ({plaintext_s1[91], plaintext_s0[91]}), .c ({signal_5573, signal_603}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_567 ( .s (reset), .b ({signal_5350, signal_3650}), .a ({plaintext_s1[92], plaintext_s0[92]}), .c ({signal_5575, signal_605}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_570 ( .s (reset), .b ({signal_5351, signal_3649}), .a ({plaintext_s1[93], plaintext_s0[93]}), .c ({signal_5577, signal_607}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_573 ( .s (reset), .b ({signal_5352, signal_3648}), .a ({plaintext_s1[94], plaintext_s0[94]}), .c ({signal_5579, signal_609}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_576 ( .s (reset), .b ({signal_5353, signal_3647}), .a ({plaintext_s1[95], plaintext_s0[95]}), .c ({signal_5581, signal_611}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_579 ( .s (reset), .b ({signal_5400, signal_3646}), .a ({plaintext_s1[96], plaintext_s0[96]}), .c ({signal_5735, signal_613}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_582 ( .s (reset), .b ({signal_5354, signal_3645}), .a ({plaintext_s1[97], plaintext_s0[97]}), .c ({signal_5583, signal_615}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_585 ( .s (reset), .b ({signal_5355, signal_3644}), .a ({plaintext_s1[98], plaintext_s0[98]}), .c ({signal_5585, signal_617}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_588 ( .s (reset), .b ({signal_5356, signal_3643}), .a ({plaintext_s1[99], plaintext_s0[99]}), .c ({signal_5587, signal_619}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_591 ( .s (reset), .b ({signal_5237, signal_3642}), .a ({plaintext_s1[100], plaintext_s0[100]}), .c ({signal_5589, signal_621}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_594 ( .s (reset), .b ({signal_5238, signal_3641}), .a ({plaintext_s1[101], plaintext_s0[101]}), .c ({signal_5591, signal_623}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_597 ( .s (reset), .b ({signal_5239, signal_3640}), .a ({plaintext_s1[102], plaintext_s0[102]}), .c ({signal_5593, signal_625}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_600 ( .s (reset), .b ({signal_5240, signal_3639}), .a ({plaintext_s1[103], plaintext_s0[103]}), .c ({signal_5595, signal_627}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_603 ( .s (reset), .b ({signal_5241, signal_3638}), .a ({plaintext_s1[104], plaintext_s0[104]}), .c ({signal_5597, signal_629}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_606 ( .s (reset), .b ({signal_5395, signal_3637}), .a ({plaintext_s1[105], plaintext_s0[105]}), .c ({signal_5737, signal_631}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_609 ( .s (reset), .b ({signal_5242, signal_3636}), .a ({plaintext_s1[106], plaintext_s0[106]}), .c ({signal_5599, signal_633}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_612 ( .s (reset), .b ({signal_5243, signal_3635}), .a ({plaintext_s1[107], plaintext_s0[107]}), .c ({signal_5601, signal_635}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_615 ( .s (reset), .b ({signal_5244, signal_3634}), .a ({plaintext_s1[108], plaintext_s0[108]}), .c ({signal_5603, signal_637}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_618 ( .s (reset), .b ({signal_5245, signal_3633}), .a ({plaintext_s1[109], plaintext_s0[109]}), .c ({signal_5605, signal_639}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_621 ( .s (reset), .b ({signal_5247, signal_3632}), .a ({plaintext_s1[110], plaintext_s0[110]}), .c ({signal_5607, signal_641}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_624 ( .s (reset), .b ({signal_5248, signal_3631}), .a ({plaintext_s1[111], plaintext_s0[111]}), .c ({signal_5609, signal_643}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_627 ( .s (reset), .b ({signal_5249, signal_3630}), .a ({plaintext_s1[112], plaintext_s0[112]}), .c ({signal_5611, signal_645}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_630 ( .s (reset), .b ({signal_5250, signal_3629}), .a ({plaintext_s1[113], plaintext_s0[113]}), .c ({signal_5613, signal_647}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_633 ( .s (reset), .b ({signal_5251, signal_3628}), .a ({plaintext_s1[114], plaintext_s0[114]}), .c ({signal_5615, signal_649}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_636 ( .s (reset), .b ({signal_5252, signal_3627}), .a ({plaintext_s1[115], plaintext_s0[115]}), .c ({signal_5617, signal_651}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_639 ( .s (reset), .b ({signal_5253, signal_3626}), .a ({plaintext_s1[116], plaintext_s0[116]}), .c ({signal_5619, signal_653}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_642 ( .s (reset), .b ({signal_5254, signal_3625}), .a ({plaintext_s1[117], plaintext_s0[117]}), .c ({signal_5621, signal_655}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_645 ( .s (reset), .b ({signal_5255, signal_3624}), .a ({plaintext_s1[118], plaintext_s0[118]}), .c ({signal_5623, signal_657}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_648 ( .s (reset), .b ({signal_5256, signal_3623}), .a ({plaintext_s1[119], plaintext_s0[119]}), .c ({signal_5625, signal_659}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_651 ( .s (reset), .b ({signal_5258, signal_3622}), .a ({plaintext_s1[120], plaintext_s0[120]}), .c ({signal_5627, signal_661}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_654 ( .s (reset), .b ({signal_5259, signal_3621}), .a ({plaintext_s1[121], plaintext_s0[121]}), .c ({signal_5629, signal_663}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_657 ( .s (reset), .b ({signal_5260, signal_3620}), .a ({plaintext_s1[122], plaintext_s0[122]}), .c ({signal_5631, signal_665}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_660 ( .s (reset), .b ({signal_5261, signal_3619}), .a ({plaintext_s1[123], plaintext_s0[123]}), .c ({signal_5633, signal_667}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_663 ( .s (reset), .b ({signal_5262, signal_3618}), .a ({plaintext_s1[124], plaintext_s0[124]}), .c ({signal_5635, signal_669}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_666 ( .s (reset), .b ({signal_5263, signal_3617}), .a ({plaintext_s1[125], plaintext_s0[125]}), .c ({signal_5637, signal_671}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_669 ( .s (reset), .b ({signal_5264, signal_3616}), .a ({plaintext_s1[126], plaintext_s0[126]}), .c ({signal_5639, signal_673}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_672 ( .s (reset), .b ({signal_5265, signal_3615}), .a ({plaintext_s1[127], plaintext_s0[127]}), .c ({signal_5641, signal_675}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_2723 ( .a ({signal_4949, signal_2597}), .b ({signal_5141, signal_4402}), .c ({signal_5357, signal_4017}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_2815 ( .a ({signal_4950, signal_2660}), .b ({signal_4973, signal_3890}), .c ({signal_5358, signal_4026}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_2831 ( .a ({signal_4951, signal_2661}), .b ({signal_5161, signal_4434}), .c ({signal_5359, signal_4049}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_2923 ( .a ({signal_4952, signal_2724}), .b ({signal_4985, signal_3922}), .c ({signal_5360, signal_4058}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_2939 ( .a ({signal_4953, signal_2725}), .b ({signal_5181, signal_4466}), .c ({signal_5361, signal_4081}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_3031 ( .a ({signal_4954, signal_2788}), .b ({signal_4997, signal_3954}), .c ({signal_5362, signal_4090}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_3047 ( .a ({signal_4955, signal_2789}), .b ({signal_5201, signal_4498}), .c ({signal_5363, signal_4113}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_3139 ( .a ({signal_4956, signal_2852}), .b ({signal_5009, signal_3986}), .c ({signal_5364, signal_4122}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3155 ( .s (reset), .b ({signal_5923, signal_4250}), .a ({key_s1[0], key_s0[0]}), .c ({signal_5925, signal_2853}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3158 ( .s (reset), .b ({signal_5912, signal_4249}), .a ({key_s1[1], key_s0[1]}), .c ({signal_5927, signal_2855}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3161 ( .s (reset), .b ({signal_5901, signal_4248}), .a ({key_s1[2], key_s0[2]}), .c ({signal_5929, signal_2857}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3164 ( .s (reset), .b ({signal_5898, signal_4247}), .a ({key_s1[3], key_s0[3]}), .c ({signal_5931, signal_2859}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3167 ( .s (reset), .b ({signal_5897, signal_4246}), .a ({key_s1[4], key_s0[4]}), .c ({signal_5933, signal_2861}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3170 ( .s (reset), .b ({signal_5896, signal_4245}), .a ({key_s1[5], key_s0[5]}), .c ({signal_5935, signal_2863}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3173 ( .s (reset), .b ({signal_5895, signal_4244}), .a ({key_s1[6], key_s0[6]}), .c ({signal_5937, signal_2865}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3176 ( .s (reset), .b ({signal_5894, signal_4243}), .a ({key_s1[7], key_s0[7]}), .c ({signal_5939, signal_2867}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3179 ( .s (reset), .b ({signal_5893, signal_4242}), .a ({key_s1[8], key_s0[8]}), .c ({signal_5941, signal_2869}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3182 ( .s (reset), .b ({signal_5892, signal_4241}), .a ({key_s1[9], key_s0[9]}), .c ({signal_5943, signal_2871}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3185 ( .s (reset), .b ({signal_5922, signal_4240}), .a ({key_s1[10], key_s0[10]}), .c ({signal_5945, signal_2873}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3188 ( .s (reset), .b ({signal_5921, signal_4239}), .a ({key_s1[11], key_s0[11]}), .c ({signal_5947, signal_2875}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3191 ( .s (reset), .b ({signal_5920, signal_4238}), .a ({key_s1[12], key_s0[12]}), .c ({signal_5949, signal_2877}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3194 ( .s (reset), .b ({signal_5919, signal_4237}), .a ({key_s1[13], key_s0[13]}), .c ({signal_5951, signal_2879}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3197 ( .s (reset), .b ({signal_5918, signal_4236}), .a ({key_s1[14], key_s0[14]}), .c ({signal_5953, signal_2881}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3200 ( .s (reset), .b ({signal_5917, signal_4235}), .a ({key_s1[15], key_s0[15]}), .c ({signal_5955, signal_2883}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3203 ( .s (reset), .b ({signal_5916, signal_4234}), .a ({key_s1[16], key_s0[16]}), .c ({signal_5957, signal_2885}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3206 ( .s (reset), .b ({signal_5915, signal_4233}), .a ({key_s1[17], key_s0[17]}), .c ({signal_5959, signal_2887}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3209 ( .s (reset), .b ({signal_5914, signal_4232}), .a ({key_s1[18], key_s0[18]}), .c ({signal_5961, signal_2889}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3212 ( .s (reset), .b ({signal_5913, signal_4231}), .a ({key_s1[19], key_s0[19]}), .c ({signal_5963, signal_2891}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3215 ( .s (reset), .b ({signal_5911, signal_4230}), .a ({key_s1[20], key_s0[20]}), .c ({signal_5965, signal_2893}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3218 ( .s (reset), .b ({signal_5910, signal_4229}), .a ({key_s1[21], key_s0[21]}), .c ({signal_5967, signal_2895}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3221 ( .s (reset), .b ({signal_5909, signal_4228}), .a ({key_s1[22], key_s0[22]}), .c ({signal_5969, signal_2897}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3224 ( .s (reset), .b ({signal_5908, signal_4227}), .a ({key_s1[23], key_s0[23]}), .c ({signal_5971, signal_2899}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3227 ( .s (reset), .b ({signal_5995, signal_4226}), .a ({key_s1[24], key_s0[24]}), .c ({signal_5997, signal_2901}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3230 ( .s (reset), .b ({signal_5994, signal_4225}), .a ({key_s1[25], key_s0[25]}), .c ({signal_5999, signal_2903}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3233 ( .s (reset), .b ({signal_6014, signal_4224}), .a ({key_s1[26], key_s0[26]}), .c ({signal_6016, signal_2905}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3236 ( .s (reset), .b ({signal_6013, signal_4223}), .a ({key_s1[27], key_s0[27]}), .c ({signal_6018, signal_2907}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3239 ( .s (reset), .b ({signal_5991, signal_4222}), .a ({key_s1[28], key_s0[28]}), .c ({signal_6001, signal_2909}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3242 ( .s (reset), .b ({signal_6012, signal_4221}), .a ({key_s1[29], key_s0[29]}), .c ({signal_6020, signal_2911}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3245 ( .s (reset), .b ({signal_5989, signal_4220}), .a ({key_s1[30], key_s0[30]}), .c ({signal_6003, signal_2913}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3248 ( .s (reset), .b ({signal_5988, signal_4219}), .a ({key_s1[31], key_s0[31]}), .c ({signal_6005, signal_2915}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3251 ( .s (reset), .b ({signal_5827, signal_4218}), .a ({key_s1[32], key_s0[32]}), .c ({signal_5829, signal_2917}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3254 ( .s (reset), .b ({signal_5813, signal_4217}), .a ({key_s1[33], key_s0[33]}), .c ({signal_5831, signal_2919}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3257 ( .s (reset), .b ({signal_5805, signal_4216}), .a ({key_s1[34], key_s0[34]}), .c ({signal_5833, signal_2921}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3260 ( .s (reset), .b ({signal_5802, signal_4215}), .a ({key_s1[35], key_s0[35]}), .c ({signal_5835, signal_2923}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3263 ( .s (reset), .b ({signal_5801, signal_4214}), .a ({key_s1[36], key_s0[36]}), .c ({signal_5837, signal_2925}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3266 ( .s (reset), .b ({signal_5800, signal_4213}), .a ({key_s1[37], key_s0[37]}), .c ({signal_5839, signal_2927}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3269 ( .s (reset), .b ({signal_5799, signal_4212}), .a ({key_s1[38], key_s0[38]}), .c ({signal_5841, signal_2929}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3272 ( .s (reset), .b ({signal_5798, signal_4211}), .a ({key_s1[39], key_s0[39]}), .c ({signal_5843, signal_2931}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3275 ( .s (reset), .b ({signal_5797, signal_4210}), .a ({key_s1[40], key_s0[40]}), .c ({signal_5845, signal_2933}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3278 ( .s (reset), .b ({signal_5796, signal_4209}), .a ({key_s1[41], key_s0[41]}), .c ({signal_5847, signal_2935}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3281 ( .s (reset), .b ({signal_5826, signal_4208}), .a ({key_s1[42], key_s0[42]}), .c ({signal_5849, signal_2937}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3284 ( .s (reset), .b ({signal_5825, signal_4207}), .a ({key_s1[43], key_s0[43]}), .c ({signal_5851, signal_2939}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3287 ( .s (reset), .b ({signal_5821, signal_4206}), .a ({key_s1[44], key_s0[44]}), .c ({signal_5853, signal_2941}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3290 ( .s (reset), .b ({signal_5820, signal_4205}), .a ({key_s1[45], key_s0[45]}), .c ({signal_5855, signal_2943}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3293 ( .s (reset), .b ({signal_5819, signal_4204}), .a ({key_s1[46], key_s0[46]}), .c ({signal_5857, signal_2945}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3296 ( .s (reset), .b ({signal_5818, signal_4203}), .a ({key_s1[47], key_s0[47]}), .c ({signal_5859, signal_2947}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3299 ( .s (reset), .b ({signal_5817, signal_4202}), .a ({key_s1[48], key_s0[48]}), .c ({signal_5861, signal_2949}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3302 ( .s (reset), .b ({signal_5816, signal_4201}), .a ({key_s1[49], key_s0[49]}), .c ({signal_5863, signal_2951}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3305 ( .s (reset), .b ({signal_5815, signal_4200}), .a ({key_s1[50], key_s0[50]}), .c ({signal_5865, signal_2953}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3308 ( .s (reset), .b ({signal_5814, signal_4199}), .a ({key_s1[51], key_s0[51]}), .c ({signal_5867, signal_2955}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3311 ( .s (reset), .b ({signal_5812, signal_4198}), .a ({key_s1[52], key_s0[52]}), .c ({signal_5869, signal_2957}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3314 ( .s (reset), .b ({signal_5811, signal_4197}), .a ({key_s1[53], key_s0[53]}), .c ({signal_5871, signal_2959}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3317 ( .s (reset), .b ({signal_5810, signal_4196}), .a ({key_s1[54], key_s0[54]}), .c ({signal_5873, signal_2961}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3320 ( .s (reset), .b ({signal_5809, signal_4195}), .a ({key_s1[55], key_s0[55]}), .c ({signal_5875, signal_2963}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3323 ( .s (reset), .b ({signal_5907, signal_4194}), .a ({key_s1[56], key_s0[56]}), .c ({signal_5973, signal_2965}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3326 ( .s (reset), .b ({signal_5906, signal_4193}), .a ({key_s1[57], key_s0[57]}), .c ({signal_5975, signal_2967}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3329 ( .s (reset), .b ({signal_5993, signal_4192}), .a ({key_s1[58], key_s0[58]}), .c ({signal_6007, signal_2969}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3332 ( .s (reset), .b ({signal_5992, signal_4191}), .a ({key_s1[59], key_s0[59]}), .c ({signal_6009, signal_2971}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3335 ( .s (reset), .b ({signal_5903, signal_4190}), .a ({key_s1[60], key_s0[60]}), .c ({signal_5977, signal_2973}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3338 ( .s (reset), .b ({signal_5990, signal_4189}), .a ({key_s1[61], key_s0[61]}), .c ({signal_6011, signal_2975}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3341 ( .s (reset), .b ({signal_5900, signal_4188}), .a ({key_s1[62], key_s0[62]}), .c ({signal_5979, signal_2977}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3344 ( .s (reset), .b ({signal_5899, signal_4187}), .a ({key_s1[63], key_s0[63]}), .c ({signal_5981, signal_2979}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3347 ( .s (reset), .b ({signal_5718, signal_4186}), .a ({key_s1[64], key_s0[64]}), .c ({signal_5739, signal_2981}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3350 ( .s (reset), .b ({signal_5702, signal_4185}), .a ({key_s1[65], key_s0[65]}), .c ({signal_5741, signal_2983}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3353 ( .s (reset), .b ({signal_5697, signal_4184}), .a ({key_s1[66], key_s0[66]}), .c ({signal_5743, signal_2985}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3356 ( .s (reset), .b ({signal_5696, signal_4183}), .a ({key_s1[67], key_s0[67]}), .c ({signal_5745, signal_2987}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3359 ( .s (reset), .b ({signal_5695, signal_4182}), .a ({key_s1[68], key_s0[68]}), .c ({signal_5747, signal_2989}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3362 ( .s (reset), .b ({signal_5694, signal_4181}), .a ({key_s1[69], key_s0[69]}), .c ({signal_5749, signal_2991}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3365 ( .s (reset), .b ({signal_5693, signal_4180}), .a ({key_s1[70], key_s0[70]}), .c ({signal_5751, signal_2993}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3368 ( .s (reset), .b ({signal_5692, signal_4179}), .a ({key_s1[71], key_s0[71]}), .c ({signal_5753, signal_2995}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3371 ( .s (reset), .b ({signal_5691, signal_4178}), .a ({key_s1[72], key_s0[72]}), .c ({signal_5755, signal_2997}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3374 ( .s (reset), .b ({signal_5690, signal_4177}), .a ({key_s1[73], key_s0[73]}), .c ({signal_5757, signal_2999}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3377 ( .s (reset), .b ({signal_5717, signal_4176}), .a ({key_s1[74], key_s0[74]}), .c ({signal_5759, signal_3001}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3380 ( .s (reset), .b ({signal_5716, signal_4175}), .a ({key_s1[75], key_s0[75]}), .c ({signal_5761, signal_3003}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3383 ( .s (reset), .b ({signal_5710, signal_4174}), .a ({key_s1[76], key_s0[76]}), .c ({signal_5763, signal_3005}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3386 ( .s (reset), .b ({signal_5709, signal_4173}), .a ({key_s1[77], key_s0[77]}), .c ({signal_5765, signal_3007}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3389 ( .s (reset), .b ({signal_5708, signal_4172}), .a ({key_s1[78], key_s0[78]}), .c ({signal_5767, signal_3009}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3392 ( .s (reset), .b ({signal_5707, signal_4171}), .a ({key_s1[79], key_s0[79]}), .c ({signal_5769, signal_3011}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3395 ( .s (reset), .b ({signal_5706, signal_4170}), .a ({key_s1[80], key_s0[80]}), .c ({signal_5771, signal_3013}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3398 ( .s (reset), .b ({signal_5705, signal_4169}), .a ({key_s1[81], key_s0[81]}), .c ({signal_5773, signal_3015}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3401 ( .s (reset), .b ({signal_5704, signal_4168}), .a ({key_s1[82], key_s0[82]}), .c ({signal_5775, signal_3017}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3404 ( .s (reset), .b ({signal_5703, signal_4167}), .a ({key_s1[83], key_s0[83]}), .c ({signal_5777, signal_3019}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3407 ( .s (reset), .b ({signal_5701, signal_4166}), .a ({key_s1[84], key_s0[84]}), .c ({signal_5779, signal_3021}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3410 ( .s (reset), .b ({signal_5700, signal_4165}), .a ({key_s1[85], key_s0[85]}), .c ({signal_5781, signal_3023}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3413 ( .s (reset), .b ({signal_5699, signal_4164}), .a ({key_s1[86], key_s0[86]}), .c ({signal_5783, signal_3025}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3416 ( .s (reset), .b ({signal_5698, signal_4163}), .a ({key_s1[87], key_s0[87]}), .c ({signal_5785, signal_3027}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3419 ( .s (reset), .b ({signal_5808, signal_4162}), .a ({key_s1[88], key_s0[88]}), .c ({signal_5877, signal_3029}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3422 ( .s (reset), .b ({signal_5807, signal_4161}), .a ({key_s1[89], key_s0[89]}), .c ({signal_5879, signal_3031}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3425 ( .s (reset), .b ({signal_5905, signal_4160}), .a ({key_s1[90], key_s0[90]}), .c ({signal_5983, signal_3033}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3428 ( .s (reset), .b ({signal_5904, signal_4159}), .a ({key_s1[91], key_s0[91]}), .c ({signal_5985, signal_3035}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3431 ( .s (reset), .b ({signal_5806, signal_4158}), .a ({key_s1[92], key_s0[92]}), .c ({signal_5881, signal_3037}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3434 ( .s (reset), .b ({signal_5902, signal_4157}), .a ({key_s1[93], key_s0[93]}), .c ({signal_5987, signal_3039}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3437 ( .s (reset), .b ({signal_5804, signal_4156}), .a ({key_s1[94], key_s0[94]}), .c ({signal_5883, signal_3041}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3440 ( .s (reset), .b ({signal_5803, signal_4155}), .a ({key_s1[95], key_s0[95]}), .c ({signal_5885, signal_3043}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3443 ( .s (reset), .b ({signal_5388, signal_4154}), .a ({key_s1[96], key_s0[96]}), .c ({signal_5643, signal_3045}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3446 ( .s (reset), .b ({signal_5367, signal_4153}), .a ({key_s1[97], key_s0[97]}), .c ({signal_5645, signal_3047}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3449 ( .s (reset), .b ({signal_5366, signal_4152}), .a ({key_s1[98], key_s0[98]}), .c ({signal_5647, signal_3049}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3452 ( .s (reset), .b ({signal_5365, signal_4151}), .a ({key_s1[99], key_s0[99]}), .c ({signal_5649, signal_3051}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3455 ( .s (reset), .b ({signal_5387, signal_4150}), .a ({key_s1[100], key_s0[100]}), .c ({signal_5651, signal_3053}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3458 ( .s (reset), .b ({signal_5386, signal_4149}), .a ({key_s1[101], key_s0[101]}), .c ({signal_5653, signal_3055}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3461 ( .s (reset), .b ({signal_5385, signal_4148}), .a ({key_s1[102], key_s0[102]}), .c ({signal_5655, signal_3057}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3464 ( .s (reset), .b ({signal_5384, signal_4147}), .a ({key_s1[103], key_s0[103]}), .c ({signal_5657, signal_3059}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3467 ( .s (reset), .b ({signal_5383, signal_4146}), .a ({key_s1[104], key_s0[104]}), .c ({signal_5659, signal_3061}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3470 ( .s (reset), .b ({signal_5382, signal_4145}), .a ({key_s1[105], key_s0[105]}), .c ({signal_5661, signal_3063}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3473 ( .s (reset), .b ({signal_5381, signal_4144}), .a ({key_s1[106], key_s0[106]}), .c ({signal_5663, signal_3065}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3476 ( .s (reset), .b ({signal_5380, signal_4143}), .a ({key_s1[107], key_s0[107]}), .c ({signal_5665, signal_3067}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3479 ( .s (reset), .b ({signal_5379, signal_4142}), .a ({key_s1[108], key_s0[108]}), .c ({signal_5667, signal_3069}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3482 ( .s (reset), .b ({signal_5378, signal_4141}), .a ({key_s1[109], key_s0[109]}), .c ({signal_5669, signal_3071}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3485 ( .s (reset), .b ({signal_5377, signal_4140}), .a ({key_s1[110], key_s0[110]}), .c ({signal_5671, signal_3073}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3488 ( .s (reset), .b ({signal_5376, signal_4139}), .a ({key_s1[111], key_s0[111]}), .c ({signal_5673, signal_3075}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3491 ( .s (reset), .b ({signal_5375, signal_4138}), .a ({key_s1[112], key_s0[112]}), .c ({signal_5675, signal_3077}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3494 ( .s (reset), .b ({signal_5374, signal_4137}), .a ({key_s1[113], key_s0[113]}), .c ({signal_5677, signal_3079}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3497 ( .s (reset), .b ({signal_5373, signal_4136}), .a ({key_s1[114], key_s0[114]}), .c ({signal_5679, signal_3081}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3500 ( .s (reset), .b ({signal_5372, signal_4135}), .a ({key_s1[115], key_s0[115]}), .c ({signal_5681, signal_3083}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3503 ( .s (reset), .b ({signal_5371, signal_4134}), .a ({key_s1[116], key_s0[116]}), .c ({signal_5683, signal_3085}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3506 ( .s (reset), .b ({signal_5370, signal_4133}), .a ({key_s1[117], key_s0[117]}), .c ({signal_5685, signal_3087}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3509 ( .s (reset), .b ({signal_5369, signal_4132}), .a ({key_s1[118], key_s0[118]}), .c ({signal_5687, signal_3089}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3512 ( .s (reset), .b ({signal_5368, signal_4131}), .a ({key_s1[119], key_s0[119]}), .c ({signal_5689, signal_3091}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3515 ( .s (reset), .b ({signal_5715, signal_4130}), .a ({key_s1[120], key_s0[120]}), .c ({signal_5787, signal_3093}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3518 ( .s (reset), .b ({signal_5714, signal_4129}), .a ({key_s1[121], key_s0[121]}), .c ({signal_5789, signal_3095}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3521 ( .s (reset), .b ({signal_5824, signal_4128}), .a ({key_s1[122], key_s0[122]}), .c ({signal_5887, signal_3097}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3524 ( .s (reset), .b ({signal_5823, signal_4127}), .a ({key_s1[123], key_s0[123]}), .c ({signal_5889, signal_3099}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3527 ( .s (reset), .b ({signal_5713, signal_4126}), .a ({key_s1[124], key_s0[124]}), .c ({signal_5791, signal_3101}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3530 ( .s (reset), .b ({signal_5822, signal_4125}), .a ({key_s1[125], key_s0[125]}), .c ({signal_5891, signal_3103}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3533 ( .s (reset), .b ({signal_5712, signal_4124}), .a ({key_s1[126], key_s0[126]}), .c ({signal_5793, signal_3105}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3536 ( .s (reset), .b ({signal_5711, signal_4123}), .a ({key_s1[127], key_s0[127]}), .c ({signal_5795, signal_3107}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3539 ( .a ({signal_4931, signal_4369}), .b ({signal_5796, signal_4209}), .c ({signal_5892, signal_4241}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3540 ( .a ({signal_4898, signal_4370}), .b ({signal_5797, signal_4210}), .c ({signal_5893, signal_4242}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3541 ( .a ({signal_4865, signal_4371}), .b ({signal_5798, signal_4211}), .c ({signal_5894, signal_4243}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3542 ( .a ({signal_4832, signal_4372}), .b ({signal_5799, signal_4212}), .c ({signal_5895, signal_4244}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3543 ( .a ({signal_4799, signal_4373}), .b ({signal_5800, signal_4213}), .c ({signal_5896, signal_4245}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3544 ( .a ({signal_4766, signal_4374}), .b ({signal_5801, signal_4214}), .c ({signal_5897, signal_4246}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3545 ( .a ({signal_4739, signal_4337}), .b ({signal_5690, signal_4177}), .c ({signal_5796, signal_4209}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3546 ( .a ({signal_4844, signal_4305}), .b ({signal_5382, signal_4145}), .c ({signal_5690, signal_4177}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3547 ( .a ({signal_4736, signal_4338}), .b ({signal_5691, signal_4178}), .c ({signal_5797, signal_4210}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3548 ( .a ({signal_4841, signal_4306}), .b ({signal_5383, signal_4146}), .c ({signal_5691, signal_4178}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3549 ( .a ({signal_4733, signal_4375}), .b ({signal_5802, signal_4215}), .c ({signal_5898, signal_4247}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3550 ( .a ({signal_4730, signal_4339}), .b ({signal_5692, signal_4179}), .c ({signal_5798, signal_4211}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3551 ( .a ({signal_4838, signal_4307}), .b ({signal_5384, signal_4147}), .c ({signal_5692, signal_4179}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3552 ( .a ({signal_4727, signal_4340}), .b ({signal_5693, signal_4180}), .c ({signal_5799, signal_4212}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3553 ( .a ({signal_4835, signal_4308}), .b ({signal_5385, signal_4148}), .c ({signal_5693, signal_4180}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3554 ( .a ({signal_4724, signal_4341}), .b ({signal_5694, signal_4181}), .c ({signal_5800, signal_4213}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3555 ( .a ({signal_4829, signal_4309}), .b ({signal_5386, signal_4149}), .c ({signal_5694, signal_4181}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3556 ( .a ({signal_4721, signal_4342}), .b ({signal_5695, signal_4182}), .c ({signal_5801, signal_4214}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3557 ( .a ({signal_4826, signal_4310}), .b ({signal_5387, signal_4150}), .c ({signal_5695, signal_4182}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3558 ( .a ({signal_4718, signal_4343}), .b ({signal_5696, signal_4183}), .c ({signal_5802, signal_4215}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3559 ( .a ({signal_4823, signal_4311}), .b ({signal_5365, signal_4151}), .c ({signal_5696, signal_4183}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3560 ( .a ({signal_4928, signal_4279}), .b ({signal_5233, signal_4545}), .c ({signal_5365, signal_4151}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3561 ( .a ({signal_4706, signal_4347}), .b ({signal_5899, signal_4187}), .c ({signal_5988, signal_4219}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3562 ( .a ({signal_4811, signal_4315}), .b ({signal_5803, signal_4155}), .c ({signal_5899, signal_4187}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3563 ( .a ({signal_4916, signal_4283}), .b ({signal_5711, signal_4123}), .c ({signal_5803, signal_4155}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3564 ( .a ({signal_4703, signal_4348}), .b ({signal_5900, signal_4188}), .c ({signal_5989, signal_4220}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3565 ( .a ({signal_4808, signal_4316}), .b ({signal_5804, signal_4156}), .c ({signal_5900, signal_4188}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3566 ( .a ({signal_4913, signal_4284}), .b ({signal_5712, signal_4124}), .c ({signal_5804, signal_4156}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3567 ( .a ({signal_4700, signal_4376}), .b ({signal_5805, signal_4216}), .c ({signal_5901, signal_4248}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3568 ( .a ({signal_4715, signal_4344}), .b ({signal_5697, signal_4184}), .c ({signal_5805, signal_4216}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3569 ( .a ({signal_4820, signal_4312}), .b ({signal_5366, signal_4152}), .c ({signal_5697, signal_4184}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3570 ( .a ({signal_4925, signal_4280}), .b ({signal_5234, signal_4546}), .c ({signal_5366, signal_4152}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3571 ( .a ({signal_4697, signal_4349}), .b ({signal_5990, signal_4189}), .c ({signal_6012, signal_4221}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3572 ( .a ({signal_4805, signal_4317}), .b ({signal_5902, signal_4157}), .c ({signal_5990, signal_4189}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3573 ( .a ({signal_4910, signal_4285}), .b ({signal_5822, signal_4125}), .c ({signal_5902, signal_4157}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3574 ( .a ({signal_4694, signal_4350}), .b ({signal_5903, signal_4190}), .c ({signal_5991, signal_4222}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3575 ( .a ({signal_4802, signal_4318}), .b ({signal_5806, signal_4158}), .c ({signal_5903, signal_4190}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3576 ( .a ({signal_4907, signal_4286}), .b ({signal_5713, signal_4126}), .c ({signal_5806, signal_4158}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3577 ( .a ({signal_4691, signal_4351}), .b ({signal_5992, signal_4191}), .c ({signal_6013, signal_4223}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3578 ( .a ({signal_4796, signal_4319}), .b ({signal_5904, signal_4159}), .c ({signal_5992, signal_4191}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3579 ( .a ({signal_4904, signal_4287}), .b ({signal_5823, signal_4127}), .c ({signal_5904, signal_4159}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3580 ( .a ({signal_4688, signal_4352}), .b ({signal_5993, signal_4192}), .c ({signal_6014, signal_4224}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3581 ( .a ({signal_4793, signal_4320}), .b ({signal_5905, signal_4160}), .c ({signal_5993, signal_4192}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3582 ( .a ({signal_4901, signal_4288}), .b ({signal_5824, signal_4128}), .c ({signal_5905, signal_4160}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3583 ( .a ({signal_4685, signal_4353}), .b ({signal_5906, signal_4193}), .c ({signal_5994, signal_4225}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3584 ( .a ({signal_4790, signal_4321}), .b ({signal_5807, signal_4161}), .c ({signal_5906, signal_4193}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3585 ( .a ({signal_4895, signal_4289}), .b ({signal_5714, signal_4129}), .c ({signal_5807, signal_4161}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3586 ( .a ({signal_4682, signal_4354}), .b ({signal_5907, signal_4194}), .c ({signal_5995, signal_4226}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3587 ( .a ({signal_4787, signal_4322}), .b ({signal_5808, signal_4162}), .c ({signal_5907, signal_4194}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3588 ( .a ({signal_4892, signal_4290}), .b ({signal_5715, signal_4130}), .c ({signal_5808, signal_4162}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3589 ( .a ({signal_4679, signal_4355}), .b ({signal_5809, signal_4195}), .c ({signal_5908, signal_4227}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3590 ( .a ({signal_4784, signal_4323}), .b ({signal_5698, signal_4163}), .c ({signal_5809, signal_4195}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3591 ( .a ({signal_4889, signal_4291}), .b ({signal_5368, signal_4131}), .c ({signal_5698, signal_4163}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3592 ( .a ({signal_4676, signal_4356}), .b ({signal_5810, signal_4196}), .c ({signal_5909, signal_4228}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3593 ( .a ({signal_4781, signal_4324}), .b ({signal_5699, signal_4164}), .c ({signal_5810, signal_4196}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3594 ( .a ({signal_4886, signal_4292}), .b ({signal_5369, signal_4132}), .c ({signal_5699, signal_4164}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3595 ( .a ({signal_4673, signal_4357}), .b ({signal_5811, signal_4197}), .c ({signal_5910, signal_4229}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3596 ( .a ({signal_4778, signal_4325}), .b ({signal_5700, signal_4165}), .c ({signal_5811, signal_4197}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3597 ( .a ({signal_4883, signal_4293}), .b ({signal_5370, signal_4133}), .c ({signal_5700, signal_4165}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3598 ( .a ({signal_4670, signal_4358}), .b ({signal_5812, signal_4198}), .c ({signal_5911, signal_4230}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3599 ( .a ({signal_4775, signal_4326}), .b ({signal_5701, signal_4166}), .c ({signal_5812, signal_4198}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3600 ( .a ({signal_4880, signal_4294}), .b ({signal_5371, signal_4134}), .c ({signal_5701, signal_4166}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3601 ( .a ({signal_4667, signal_4377}), .b ({signal_5813, signal_4217}), .c ({signal_5912, signal_4249}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3602 ( .a ({signal_4712, signal_4345}), .b ({signal_5702, signal_4185}), .c ({signal_5813, signal_4217}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3603 ( .a ({signal_4817, signal_4313}), .b ({signal_5367, signal_4153}), .c ({signal_5702, signal_4185}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3604 ( .a ({signal_4922, signal_4281}), .b ({signal_5235, signal_4547}), .c ({signal_5367, signal_4153}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3605 ( .a ({signal_4664, signal_4359}), .b ({signal_5814, signal_4199}), .c ({signal_5913, signal_4231}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3606 ( .a ({signal_4772, signal_4327}), .b ({signal_5703, signal_4167}), .c ({signal_5814, signal_4199}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3607 ( .a ({signal_4877, signal_4295}), .b ({signal_5372, signal_4135}), .c ({signal_5703, signal_4167}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3608 ( .a ({signal_4661, signal_4360}), .b ({signal_5815, signal_4200}), .c ({signal_5914, signal_4232}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3609 ( .a ({signal_4769, signal_4328}), .b ({signal_5704, signal_4168}), .c ({signal_5815, signal_4200}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3610 ( .a ({signal_4874, signal_4296}), .b ({signal_5373, signal_4136}), .c ({signal_5704, signal_4168}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3611 ( .a ({signal_4658, signal_4361}), .b ({signal_5816, signal_4201}), .c ({signal_5915, signal_4233}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3612 ( .a ({signal_4763, signal_4329}), .b ({signal_5705, signal_4169}), .c ({signal_5816, signal_4201}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3613 ( .a ({signal_4871, signal_4297}), .b ({signal_5374, signal_4137}), .c ({signal_5705, signal_4169}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3614 ( .a ({signal_4655, signal_4362}), .b ({signal_5817, signal_4202}), .c ({signal_5916, signal_4234}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3615 ( .a ({signal_4760, signal_4330}), .b ({signal_5706, signal_4170}), .c ({signal_5817, signal_4202}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3616 ( .a ({signal_4868, signal_4298}), .b ({signal_5375, signal_4138}), .c ({signal_5706, signal_4170}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3617 ( .a ({signal_4652, signal_4363}), .b ({signal_5818, signal_4203}), .c ({signal_5917, signal_4235}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3618 ( .a ({signal_4757, signal_4331}), .b ({signal_5707, signal_4171}), .c ({signal_5818, signal_4203}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3619 ( .a ({signal_4862, signal_4299}), .b ({signal_5376, signal_4139}), .c ({signal_5707, signal_4171}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3620 ( .a ({signal_4649, signal_4364}), .b ({signal_5819, signal_4204}), .c ({signal_5918, signal_4236}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3621 ( .a ({signal_4754, signal_4332}), .b ({signal_5708, signal_4172}), .c ({signal_5819, signal_4204}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3622 ( .a ({signal_4859, signal_4300}), .b ({signal_5377, signal_4140}), .c ({signal_5708, signal_4172}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3623 ( .a ({signal_4646, signal_4365}), .b ({signal_5820, signal_4205}), .c ({signal_5919, signal_4237}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3624 ( .a ({signal_4751, signal_4333}), .b ({signal_5709, signal_4173}), .c ({signal_5820, signal_4205}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3625 ( .a ({signal_4856, signal_4301}), .b ({signal_5378, signal_4141}), .c ({signal_5709, signal_4173}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3626 ( .a ({signal_4643, signal_4366}), .b ({signal_5821, signal_4206}), .c ({signal_5920, signal_4238}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3627 ( .a ({signal_4748, signal_4334}), .b ({signal_5710, signal_4174}), .c ({signal_5821, signal_4206}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3628 ( .a ({signal_4853, signal_4302}), .b ({signal_5379, signal_4142}), .c ({signal_5710, signal_4174}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3629 ( .a ({signal_4640, signal_4251}), .b ({signal_5389, signal_4517}), .c ({signal_5711, signal_4123}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3630 ( .a ({signal_4637, signal_4252}), .b ({signal_5390, signal_4518}), .c ({signal_5712, signal_4124}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3631 ( .a ({signal_4634, signal_4253}), .b ({signal_5719, signal_4519}), .c ({signal_5822, signal_4125}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3632 ( .a ({signal_4631, signal_4254}), .b ({signal_5391, signal_4520}), .c ({signal_5713, signal_4126}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3633 ( .a ({signal_4628, signal_4255}), .b ({signal_5720, signal_4521}), .c ({signal_5823, signal_4127}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3634 ( .a ({signal_4625, signal_4256}), .b ({signal_5721, signal_4522}), .c ({signal_5824, signal_4128}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3635 ( .a ({signal_4622, signal_4257}), .b ({signal_5392, signal_4523}), .c ({signal_5714, signal_4129}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3636 ( .a ({signal_4619, signal_4258}), .b ({signal_5393, signal_4524}), .c ({signal_5715, signal_4130}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3637 ( .a ({signal_4616, signal_4367}), .b ({signal_5825, signal_4207}), .c ({signal_5921, signal_4239}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3638 ( .a ({signal_4745, signal_4335}), .b ({signal_5716, signal_4175}), .c ({signal_5825, signal_4207}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3639 ( .a ({signal_4850, signal_4303}), .b ({signal_5380, signal_4143}), .c ({signal_5716, signal_4175}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3640 ( .a ({signal_4613, signal_4259}), .b ({signal_5213, signal_4525}), .c ({signal_5368, signal_4131}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3641 ( .a ({signal_4610, signal_4260}), .b ({signal_5214, signal_4526}), .c ({signal_5369, signal_4132}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3642 ( .a ({signal_4607, signal_4261}), .b ({signal_5215, signal_4527}), .c ({signal_5370, signal_4133}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3643 ( .a ({signal_4604, signal_4262}), .b ({signal_5216, signal_4528}), .c ({signal_5371, signal_4134}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3644 ( .a ({signal_4601, signal_4263}), .b ({signal_5217, signal_4529}), .c ({signal_5372, signal_4135}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3645 ( .a ({signal_4598, signal_4264}), .b ({signal_5218, signal_4530}), .c ({signal_5373, signal_4136}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3646 ( .a ({signal_4595, signal_4265}), .b ({signal_5219, signal_4531}), .c ({signal_5374, signal_4137}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3647 ( .a ({signal_4592, signal_4266}), .b ({signal_5220, signal_4532}), .c ({signal_5375, signal_4138}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3648 ( .a ({signal_4589, signal_4267}), .b ({signal_5221, signal_4533}), .c ({signal_5376, signal_4139}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3649 ( .a ({signal_4586, signal_4268}), .b ({signal_5222, signal_4534}), .c ({signal_5377, signal_4140}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3650 ( .a ({signal_4583, signal_4368}), .b ({signal_5826, signal_4208}), .c ({signal_5922, signal_4240}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3651 ( .a ({signal_4742, signal_4336}), .b ({signal_5717, signal_4176}), .c ({signal_5826, signal_4208}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3652 ( .a ({signal_4847, signal_4304}), .b ({signal_5381, signal_4144}), .c ({signal_5717, signal_4176}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3653 ( .a ({signal_4580, signal_4269}), .b ({signal_5223, signal_4535}), .c ({signal_5378, signal_4141}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3654 ( .a ({signal_4577, signal_4270}), .b ({signal_5224, signal_4536}), .c ({signal_5379, signal_4142}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3655 ( .a ({signal_4574, signal_4271}), .b ({signal_5225, signal_4537}), .c ({signal_5380, signal_4143}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3656 ( .a ({signal_4571, signal_4272}), .b ({signal_5226, signal_4538}), .c ({signal_5381, signal_4144}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3657 ( .a ({signal_4568, signal_4273}), .b ({signal_5227, signal_4539}), .c ({signal_5382, signal_4145}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3658 ( .a ({signal_4565, signal_4274}), .b ({signal_5228, signal_4540}), .c ({signal_5383, signal_4146}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3659 ( .a ({signal_4562, signal_4275}), .b ({signal_5229, signal_4541}), .c ({signal_5384, signal_4147}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3660 ( .a ({signal_4559, signal_4276}), .b ({signal_5230, signal_4542}), .c ({signal_5385, signal_4148}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3661 ( .a ({signal_4556, signal_4277}), .b ({signal_5231, signal_4543}), .c ({signal_5386, signal_4149}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3662 ( .a ({signal_4553, signal_4278}), .b ({signal_5232, signal_4544}), .c ({signal_5387, signal_4150}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3663 ( .a ({signal_4550, signal_4378}), .b ({signal_5827, signal_4218}), .c ({signal_5923, signal_4250}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3664 ( .a ({signal_4709, signal_4346}), .b ({signal_5718, signal_4186}), .c ({signal_5827, signal_4218}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3665 ( .a ({signal_4814, signal_4314}), .b ({signal_5388, signal_4154}), .c ({signal_5718, signal_4186}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3666 ( .a ({signal_4919, signal_4282}), .b ({signal_5236, signal_4548}), .c ({signal_5388, signal_4154}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3667 ( .a ({signal_4964, signal_3116}), .b ({1'b0, signal_393}), .c ({signal_5389, signal_4517}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3668 ( .a ({signal_4963, signal_3115}), .b ({1'b0, signal_394}), .c ({signal_5390, signal_4518}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3669 ( .a ({signal_4962, signal_3114}), .b ({1'b0, signal_4379}), .c ({signal_5719, signal_4519}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3670 ( .a ({signal_4961, signal_3113}), .b ({1'b0, signal_4380}), .c ({signal_5391, signal_4520}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3671 ( .a ({signal_4960, signal_3112}), .b ({1'b0, signal_4381}), .c ({signal_5720, signal_4521}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3672 ( .a ({signal_4959, signal_3111}), .b ({1'b0, signal_4382}), .c ({signal_5721, signal_4522}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3673 ( .a ({signal_4958, signal_3110}), .b ({1'b0, signal_4383}), .c ({signal_5392, signal_4523}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3674 ( .a ({signal_4957, signal_3109}), .b ({1'b0, signal_4384}), .c ({signal_5393, signal_4524}) ) ;
    AES_step2_ANF #(.low_latency(0), .pipeline(0)) cell_4209 ( .in0 ({signal_912, signal_792, signal_4378, signal_4377, signal_4376, signal_4375, signal_4374, signal_4373, signal_4372, signal_4371, signal_4370, signal_4369, signal_4368, signal_4367, signal_4366, signal_4365, signal_4364, signal_4363, signal_4362, signal_4361, signal_4360, signal_4359, signal_4358, signal_4357, signal_4356, signal_4355, signal_4354, signal_4353, signal_4352, signal_4351, signal_4350, signal_4349, signal_4348, signal_4347, ciphertext_s0[0], ciphertext_s0[1], ciphertext_s0[2], ciphertext_s0[4], ciphertext_s0[5], ciphertext_s0[6], ciphertext_s0[7], ciphertext_s0[8], ciphertext_s0[9], ciphertext_s0[10], ciphertext_s0[12], ciphertext_s0[13], ciphertext_s0[14], ciphertext_s0[15], ciphertext_s0[16], ciphertext_s0[17], ciphertext_s0[18], ciphertext_s0[20], ciphertext_s0[21], ciphertext_s0[22], ciphertext_s0[23], ciphertext_s0[24], ciphertext_s0[25], ciphertext_s0[26], ciphertext_s0[28], ciphertext_s0[29], ciphertext_s0[30], ciphertext_s0[31], ciphertext_s0[32], ciphertext_s0[33], ciphertext_s0[34], ciphertext_s0[36], ciphertext_s0[37], ciphertext_s0[38], ciphertext_s0[39], ciphertext_s0[40], ciphertext_s0[41], ciphertext_s0[42], ciphertext_s0[44], ciphertext_s0[45], ciphertext_s0[46], ciphertext_s0[47], ciphertext_s0[48], ciphertext_s0[49], ciphertext_s0[50], ciphertext_s0[52], ciphertext_s0[53], ciphertext_s0[54], ciphertext_s0[55], ciphertext_s0[56], ciphertext_s0[57], ciphertext_s0[58], ciphertext_s0[60], ciphertext_s0[61], ciphertext_s0[62], ciphertext_s0[63], ciphertext_s0[64], ciphertext_s0[65], ciphertext_s0[66], ciphertext_s0[68], ciphertext_s0[69], ciphertext_s0[70], ciphertext_s0[71], ciphertext_s0[72], ciphertext_s0[73], ciphertext_s0[74], ciphertext_s0[76], ciphertext_s0[77], ciphertext_s0[78], ciphertext_s0[79], ciphertext_s0[80], ciphertext_s0[81], ciphertext_s0[82], ciphertext_s0[84], ciphertext_s0[85], ciphertext_s0[86], ciphertext_s0[87], ciphertext_s0[88], ciphertext_s0[89], ciphertext_s0[90], ciphertext_s0[92], ciphertext_s0[93], ciphertext_s0[94], ciphertext_s0[95], ciphertext_s0[96], ciphertext_s0[97], ciphertext_s0[98], ciphertext_s0[100], ciphertext_s0[101], ciphertext_s0[102], ciphertext_s0[103], ciphertext_s0[104], ciphertext_s0[105], ciphertext_s0[106], ciphertext_s0[108], ciphertext_s0[109], ciphertext_s0[110], ciphertext_s0[111], ciphertext_s0[112], ciphertext_s0[113], ciphertext_s0[114], ciphertext_s0[116], ciphertext_s0[117], ciphertext_s0[118], ciphertext_s0[119], ciphertext_s0[120], ciphertext_s0[121], ciphertext_s0[122], ciphertext_s0[124], ciphertext_s0[125], ciphertext_s0[126], ciphertext_s0[127], signal_2592, signal_2472, signal_2352, signal_2232, signal_2112, signal_1992, signal_1872, signal_1752, signal_1632, signal_1512, signal_1392, signal_1272, signal_1152, signal_1032}), .in1 ({signal_4934, signal_4933, signal_4550, signal_4667, signal_4700, signal_4733, signal_4766, signal_4799, signal_4832, signal_4865, signal_4898, signal_4931, signal_4583, signal_4616, signal_4643, signal_4646, signal_4649, signal_4652, signal_4655, signal_4658, signal_4661, signal_4664, signal_4670, signal_4673, signal_4676, signal_4679, signal_4682, signal_4685, signal_4688, signal_4691, signal_4694, signal_4697, signal_4703, signal_4706, ciphertext_s1[0], ciphertext_s1[1], ciphertext_s1[2], ciphertext_s1[4], ciphertext_s1[5], ciphertext_s1[6], ciphertext_s1[7], ciphertext_s1[8], ciphertext_s1[9], ciphertext_s1[10], ciphertext_s1[12], ciphertext_s1[13], ciphertext_s1[14], ciphertext_s1[15], ciphertext_s1[16], ciphertext_s1[17], ciphertext_s1[18], ciphertext_s1[20], ciphertext_s1[21], ciphertext_s1[22], ciphertext_s1[23], ciphertext_s1[24], ciphertext_s1[25], ciphertext_s1[26], ciphertext_s1[28], ciphertext_s1[29], ciphertext_s1[30], ciphertext_s1[31], ciphertext_s1[32], ciphertext_s1[33], ciphertext_s1[34], ciphertext_s1[36], ciphertext_s1[37], ciphertext_s1[38], ciphertext_s1[39], ciphertext_s1[40], ciphertext_s1[41], ciphertext_s1[42], ciphertext_s1[44], ciphertext_s1[45], ciphertext_s1[46], ciphertext_s1[47], ciphertext_s1[48], ciphertext_s1[49], ciphertext_s1[50], ciphertext_s1[52], ciphertext_s1[53], ciphertext_s1[54], ciphertext_s1[55], ciphertext_s1[56], ciphertext_s1[57], ciphertext_s1[58], ciphertext_s1[60], ciphertext_s1[61], ciphertext_s1[62], ciphertext_s1[63], ciphertext_s1[64], ciphertext_s1[65], ciphertext_s1[66], ciphertext_s1[68], ciphertext_s1[69], ciphertext_s1[70], ciphertext_s1[71], ciphertext_s1[72], ciphertext_s1[73], ciphertext_s1[74], ciphertext_s1[76], ciphertext_s1[77], ciphertext_s1[78], ciphertext_s1[79], ciphertext_s1[80], ciphertext_s1[81], ciphertext_s1[82], ciphertext_s1[84], ciphertext_s1[85], ciphertext_s1[86], ciphertext_s1[87], ciphertext_s1[88], ciphertext_s1[89], ciphertext_s1[90], ciphertext_s1[92], ciphertext_s1[93], ciphertext_s1[94], ciphertext_s1[95], ciphertext_s1[96], ciphertext_s1[97], ciphertext_s1[98], ciphertext_s1[100], ciphertext_s1[101], ciphertext_s1[102], ciphertext_s1[103], ciphertext_s1[104], ciphertext_s1[105], ciphertext_s1[106], ciphertext_s1[108], ciphertext_s1[109], ciphertext_s1[110], ciphertext_s1[111], ciphertext_s1[112], ciphertext_s1[113], ciphertext_s1[114], ciphertext_s1[116], ciphertext_s1[117], ciphertext_s1[118], ciphertext_s1[119], ciphertext_s1[120], ciphertext_s1[121], ciphertext_s1[122], ciphertext_s1[124], ciphertext_s1[125], ciphertext_s1[126], ciphertext_s1[127], signal_4948, signal_4947, signal_4946, signal_4945, signal_4944, signal_4943, signal_4942, signal_4941, signal_4940, signal_4939, signal_4938, signal_4937, signal_4936, signal_4935}), .clk (clk), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_4548, signal_4547, signal_4546, signal_4545, signal_4544, signal_4543, signal_4542, signal_4541, signal_4540, signal_4539, signal_4538, signal_4537, signal_4536, signal_4535, signal_4534, signal_4533, signal_4532, signal_4531, signal_4530, signal_4529, signal_4528, signal_4527, signal_4526, signal_4525, signal_4516, signal_4514, signal_4511, signal_4510, signal_4509, signal_4508, signal_4506, signal_4503, signal_4502, signal_4501, signal_4500, signal_4498, signal_4495, signal_4494, signal_4493, signal_4492, signal_4490, signal_4487, signal_4486, signal_4485, signal_4484, signal_4482, signal_4479, signal_4478, signal_4477, signal_4476, signal_4474, signal_4471, signal_4470, signal_4469, signal_4468, signal_4466, signal_4463, signal_4462, signal_4461, signal_4460, signal_4458, signal_4455, signal_4454, signal_4453, signal_4452, signal_4450, signal_4447, signal_4446, signal_4445, signal_4444, signal_4442, signal_4439, signal_4438, signal_4437, signal_4436, signal_4434, signal_4431, signal_4430, signal_4429, signal_4428, signal_4426, signal_4423, signal_4422, signal_4421, signal_4420, signal_4418, signal_4415, signal_4414, signal_4413, signal_4412, signal_4410, signal_4407, signal_4406, signal_4405, signal_4404, signal_4402, signal_4399, signal_4398, signal_4397, signal_4396, signal_4394, signal_4391, signal_4390, signal_4389, signal_4121, signal_4120, signal_4119, signal_4118, signal_4117, signal_4116, signal_4115, signal_4114, signal_4112, signal_4111, signal_4110, signal_4109, signal_4108, signal_4107, signal_4106, signal_4105, signal_4104, signal_4103, signal_4102, signal_4101, signal_4100, signal_4099, signal_4098, signal_4097, signal_4096, signal_4095, signal_4094, signal_4093, signal_4092, signal_4091, signal_4089, signal_4088, signal_4087, signal_4086, signal_4085, signal_4084, signal_4083, signal_4082, signal_4080, signal_4079, signal_4078, signal_4077, signal_4076, signal_4075, signal_4074, signal_4073, signal_4072, signal_4071, signal_4070, signal_4069, signal_4068, signal_4067, signal_4066, signal_4065, signal_4064, signal_4063, signal_4062, signal_4061, signal_4060, signal_4059, signal_4057, signal_4056, signal_4055, signal_4054, signal_4053, signal_4052, signal_4051, signal_4050, signal_4048, signal_4047, signal_4046, signal_4045, signal_4044, signal_4043, signal_4042, signal_4041, signal_4040, signal_4039, signal_4038, signal_4037, signal_4036, signal_4035, signal_4034, signal_4033, signal_4032, signal_4031, signal_4030, signal_4029, signal_4028, signal_4027, signal_4025, signal_4024, signal_4023, signal_4022, signal_4021, signal_4020, signal_4019, signal_4018, signal_4016, signal_4015, signal_4014, signal_4013, signal_4012, signal_4011, signal_4010, signal_4009, signal_4008, signal_4007, signal_4006, signal_4005, signal_4004, signal_4003, signal_4002, signal_4001, signal_4000, signal_3999, signal_3998, signal_3997, signal_3996, signal_3995, signal_3994, signal_3992, signal_3991, signal_3986, signal_3984, signal_3983, signal_3978, signal_3976, signal_3975, signal_3970, signal_3968, signal_3967, signal_3962, signal_3960, signal_3959, signal_3954, signal_3952, signal_3951, signal_3946, signal_3944, signal_3943, signal_3938, signal_3936, signal_3935, signal_3930, signal_3928, signal_3927, signal_3922, signal_3920, signal_3919, signal_3914, signal_3912, signal_3911, signal_3906, signal_3904, signal_3903, signal_3898, signal_3896, signal_3895, signal_3890, signal_3888, signal_3887, signal_3882, signal_3880, signal_3879, signal_3874, signal_3872, signal_3871, signal_3116, signal_3115, signal_3114, signal_3113, signal_3112, signal_3111, signal_3110, signal_3109, signal_2852, signal_2789, signal_2788, signal_2725, signal_2724, signal_2661, signal_2660, signal_2597}), .out1 ({signal_5236, signal_5235, signal_5234, signal_5233, signal_5232, signal_5231, signal_5230, signal_5229, signal_5228, signal_5227, signal_5226, signal_5225, signal_5224, signal_5223, signal_5222, signal_5221, signal_5220, signal_5219, signal_5218, signal_5217, signal_5216, signal_5215, signal_5214, signal_5213, signal_5212, signal_5211, signal_5210, signal_5209, signal_5208, signal_5207, signal_5206, signal_5205, signal_5204, signal_5203, signal_5202, signal_5201, signal_5200, signal_5199, signal_5198, signal_5197, signal_5196, signal_5195, signal_5194, signal_5193, signal_5192, signal_5191, signal_5190, signal_5189, signal_5188, signal_5187, signal_5186, signal_5185, signal_5184, signal_5183, signal_5182, signal_5181, signal_5180, signal_5179, signal_5178, signal_5177, signal_5176, signal_5175, signal_5174, signal_5173, signal_5172, signal_5171, signal_5170, signal_5169, signal_5168, signal_5167, signal_5166, signal_5165, signal_5164, signal_5163, signal_5162, signal_5161, signal_5160, signal_5159, signal_5158, signal_5157, signal_5156, signal_5155, signal_5154, signal_5153, signal_5152, signal_5151, signal_5150, signal_5149, signal_5148, signal_5147, signal_5146, signal_5145, signal_5144, signal_5143, signal_5142, signal_5141, signal_5140, signal_5139, signal_5138, signal_5137, signal_5136, signal_5135, signal_5134, signal_5133, signal_5132, signal_5131, signal_5130, signal_5129, signal_5128, signal_5127, signal_5126, signal_5125, signal_5124, signal_5123, signal_5122, signal_5121, signal_5120, signal_5119, signal_5118, signal_5117, signal_5116, signal_5115, signal_5114, signal_5113, signal_5112, signal_5111, signal_5110, signal_5109, signal_5108, signal_5107, signal_5106, signal_5105, signal_5104, signal_5103, signal_5102, signal_5101, signal_5100, signal_5099, signal_5098, signal_5097, signal_5096, signal_5095, signal_5094, signal_5093, signal_5092, signal_5091, signal_5090, signal_5089, signal_5088, signal_5087, signal_5086, signal_5085, signal_5084, signal_5083, signal_5082, signal_5081, signal_5080, signal_5079, signal_5078, signal_5077, signal_5076, signal_5075, signal_5074, signal_5073, signal_5072, signal_5071, signal_5070, signal_5069, signal_5068, signal_5067, signal_5066, signal_5065, signal_5064, signal_5063, signal_5062, signal_5061, signal_5060, signal_5059, signal_5058, signal_5057, signal_5056, signal_5055, signal_5054, signal_5053, signal_5052, signal_5051, signal_5050, signal_5049, signal_5048, signal_5047, signal_5046, signal_5045, signal_5044, signal_5043, signal_5042, signal_5041, signal_5040, signal_5039, signal_5038, signal_5037, signal_5036, signal_5035, signal_5034, signal_5033, signal_5032, signal_5031, signal_5030, signal_5029, signal_5028, signal_5027, signal_5026, signal_5025, signal_5024, signal_5023, signal_5022, signal_5021, signal_5020, signal_5019, signal_5018, signal_5017, signal_5016, signal_5015, signal_5014, signal_5013, signal_5012, signal_5011, signal_5010, signal_5009, signal_5008, signal_5007, signal_5006, signal_5005, signal_5004, signal_5003, signal_5002, signal_5001, signal_5000, signal_4999, signal_4998, signal_4997, signal_4996, signal_4995, signal_4994, signal_4993, signal_4992, signal_4991, signal_4990, signal_4989, signal_4988, signal_4987, signal_4986, signal_4985, signal_4984, signal_4983, signal_4982, signal_4981, signal_4980, signal_4979, signal_4978, signal_4977, signal_4976, signal_4975, signal_4974, signal_4973, signal_4972, signal_4971, signal_4970, signal_4969, signal_4968, signal_4967, signal_4966, signal_4965, signal_4964, signal_4963, signal_4962, signal_4961, signal_4960, signal_4959, signal_4958, signal_4957, signal_4956, signal_4955, signal_4954, signal_4953, signal_4952, signal_4951, signal_4950, signal_4949}) ) ;

    /* register cells */
    reg_masked #(.low_latency(0), .pipeline(0)) cell_293 ( .clk (signal_6181), .D ({signal_5723, signal_421}), .Q ({signal_4549, signal_3870}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_296 ( .clk (signal_6181), .D ({signal_5403, signal_423}), .Q ({signal_4666, signal_3869}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_299 ( .clk (signal_6181), .D ({signal_5405, signal_425}), .Q ({signal_4699, signal_3868}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_302 ( .clk (signal_6181), .D ({signal_5407, signal_427}), .Q ({signal_4732, signal_3867}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_305 ( .clk (signal_6181), .D ({signal_5409, signal_429}), .Q ({signal_4765, signal_3866}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_308 ( .clk (signal_6181), .D ({signal_5411, signal_431}), .Q ({signal_4798, signal_3865}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_311 ( .clk (signal_6181), .D ({signal_5413, signal_433}), .Q ({signal_4831, signal_3864}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_314 ( .clk (signal_6181), .D ({signal_5415, signal_435}), .Q ({signal_4864, signal_3863}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_317 ( .clk (signal_6181), .D ({signal_5417, signal_437}), .Q ({signal_4897, signal_3862}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_320 ( .clk (signal_6181), .D ({signal_5725, signal_439}), .Q ({signal_4930, signal_3861}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_323 ( .clk (signal_6181), .D ({signal_5419, signal_441}), .Q ({signal_4582, signal_3860}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_326 ( .clk (signal_6181), .D ({signal_5421, signal_443}), .Q ({signal_4615, signal_3859}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_329 ( .clk (signal_6181), .D ({signal_5423, signal_445}), .Q ({signal_4642, signal_3858}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_332 ( .clk (signal_6181), .D ({signal_5425, signal_447}), .Q ({signal_4645, signal_3857}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_335 ( .clk (signal_6181), .D ({signal_5427, signal_449}), .Q ({signal_4648, signal_3856}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_338 ( .clk (signal_6181), .D ({signal_5429, signal_451}), .Q ({signal_4651, signal_3855}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_341 ( .clk (signal_6181), .D ({signal_5431, signal_453}), .Q ({signal_4654, signal_3854}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_344 ( .clk (signal_6181), .D ({signal_5433, signal_455}), .Q ({signal_4657, signal_3853}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_347 ( .clk (signal_6181), .D ({signal_5435, signal_457}), .Q ({signal_4660, signal_3852}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_350 ( .clk (signal_6181), .D ({signal_5437, signal_459}), .Q ({signal_4663, signal_3851}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_353 ( .clk (signal_6181), .D ({signal_5439, signal_461}), .Q ({signal_4669, signal_3850}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_356 ( .clk (signal_6181), .D ({signal_5441, signal_463}), .Q ({signal_4672, signal_3849}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_359 ( .clk (signal_6181), .D ({signal_5443, signal_465}), .Q ({signal_4675, signal_3848}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_362 ( .clk (signal_6181), .D ({signal_5445, signal_467}), .Q ({signal_4678, signal_3847}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_365 ( .clk (signal_6181), .D ({signal_5447, signal_469}), .Q ({signal_4681, signal_3846}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_368 ( .clk (signal_6181), .D ({signal_5449, signal_471}), .Q ({signal_4684, signal_3845}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_371 ( .clk (signal_6181), .D ({signal_5451, signal_473}), .Q ({signal_4687, signal_3844}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_374 ( .clk (signal_6181), .D ({signal_5453, signal_475}), .Q ({signal_4690, signal_3843}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_377 ( .clk (signal_6181), .D ({signal_5455, signal_477}), .Q ({signal_4693, signal_3842}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_380 ( .clk (signal_6181), .D ({signal_5457, signal_479}), .Q ({signal_4696, signal_3841}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_383 ( .clk (signal_6181), .D ({signal_5459, signal_481}), .Q ({signal_4702, signal_3840}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_386 ( .clk (signal_6181), .D ({signal_5461, signal_483}), .Q ({signal_4705, signal_3839}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_389 ( .clk (signal_6181), .D ({signal_5727, signal_485}), .Q ({signal_4708, signal_3838}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_392 ( .clk (signal_6181), .D ({signal_5463, signal_487}), .Q ({signal_4711, signal_3837}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_395 ( .clk (signal_6181), .D ({signal_5465, signal_489}), .Q ({signal_4714, signal_3836}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_398 ( .clk (signal_6181), .D ({signal_5467, signal_491}), .Q ({signal_4717, signal_3835}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_401 ( .clk (signal_6181), .D ({signal_5469, signal_493}), .Q ({signal_4720, signal_3834}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_404 ( .clk (signal_6181), .D ({signal_5471, signal_495}), .Q ({signal_4723, signal_3833}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_407 ( .clk (signal_6181), .D ({signal_5473, signal_497}), .Q ({signal_4726, signal_3832}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_410 ( .clk (signal_6181), .D ({signal_5475, signal_499}), .Q ({signal_4729, signal_3831}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_413 ( .clk (signal_6181), .D ({signal_5477, signal_501}), .Q ({signal_4735, signal_3830}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_416 ( .clk (signal_6181), .D ({signal_5729, signal_503}), .Q ({signal_4738, signal_3829}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_419 ( .clk (signal_6181), .D ({signal_5479, signal_505}), .Q ({signal_4741, signal_3828}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_422 ( .clk (signal_6181), .D ({signal_5481, signal_507}), .Q ({signal_4744, signal_3827}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_425 ( .clk (signal_6181), .D ({signal_5483, signal_509}), .Q ({signal_4747, signal_3826}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_428 ( .clk (signal_6181), .D ({signal_5485, signal_511}), .Q ({signal_4750, signal_3825}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_431 ( .clk (signal_6181), .D ({signal_5487, signal_513}), .Q ({signal_4753, signal_3824}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_434 ( .clk (signal_6181), .D ({signal_5489, signal_515}), .Q ({signal_4756, signal_3823}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_437 ( .clk (signal_6181), .D ({signal_5491, signal_517}), .Q ({signal_4759, signal_3822}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_440 ( .clk (signal_6181), .D ({signal_5493, signal_519}), .Q ({signal_4762, signal_3821}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_443 ( .clk (signal_6181), .D ({signal_5495, signal_521}), .Q ({signal_4768, signal_3820}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_446 ( .clk (signal_6181), .D ({signal_5497, signal_523}), .Q ({signal_4771, signal_3819}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_449 ( .clk (signal_6181), .D ({signal_5499, signal_525}), .Q ({signal_4774, signal_3818}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_452 ( .clk (signal_6181), .D ({signal_5501, signal_527}), .Q ({signal_4777, signal_3817}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_455 ( .clk (signal_6181), .D ({signal_5503, signal_529}), .Q ({signal_4780, signal_3816}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_458 ( .clk (signal_6181), .D ({signal_5505, signal_531}), .Q ({signal_4783, signal_3815}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_461 ( .clk (signal_6181), .D ({signal_5507, signal_533}), .Q ({signal_4786, signal_3814}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_464 ( .clk (signal_6181), .D ({signal_5509, signal_535}), .Q ({signal_4789, signal_3813}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_467 ( .clk (signal_6181), .D ({signal_5511, signal_537}), .Q ({signal_4792, signal_3812}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_470 ( .clk (signal_6181), .D ({signal_5513, signal_539}), .Q ({signal_4795, signal_3811}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_473 ( .clk (signal_6181), .D ({signal_5515, signal_541}), .Q ({signal_4801, signal_3810}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_476 ( .clk (signal_6181), .D ({signal_5517, signal_543}), .Q ({signal_4804, signal_3809}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_479 ( .clk (signal_6181), .D ({signal_5519, signal_545}), .Q ({signal_4807, signal_3808}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_482 ( .clk (signal_6181), .D ({signal_5521, signal_547}), .Q ({signal_4810, signal_3807}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_485 ( .clk (signal_6181), .D ({signal_5731, signal_549}), .Q ({signal_4813, signal_3806}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_488 ( .clk (signal_6181), .D ({signal_5523, signal_551}), .Q ({signal_4816, signal_3805}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_491 ( .clk (signal_6181), .D ({signal_5525, signal_553}), .Q ({signal_4819, signal_3804}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_494 ( .clk (signal_6181), .D ({signal_5527, signal_555}), .Q ({signal_4822, signal_3803}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_497 ( .clk (signal_6181), .D ({signal_5529, signal_557}), .Q ({signal_4825, signal_3802}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_500 ( .clk (signal_6181), .D ({signal_5531, signal_559}), .Q ({signal_4828, signal_3801}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_503 ( .clk (signal_6181), .D ({signal_5533, signal_561}), .Q ({signal_4834, signal_3800}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_506 ( .clk (signal_6181), .D ({signal_5535, signal_563}), .Q ({signal_4837, signal_3799}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_509 ( .clk (signal_6181), .D ({signal_5537, signal_565}), .Q ({signal_4840, signal_3798}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_512 ( .clk (signal_6181), .D ({signal_5733, signal_567}), .Q ({signal_4843, signal_3797}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_515 ( .clk (signal_6181), .D ({signal_5539, signal_569}), .Q ({signal_4846, signal_3796}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_518 ( .clk (signal_6181), .D ({signal_5541, signal_571}), .Q ({signal_4849, signal_3795}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_521 ( .clk (signal_6181), .D ({signal_5543, signal_573}), .Q ({signal_4852, signal_3794}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_524 ( .clk (signal_6181), .D ({signal_5545, signal_575}), .Q ({signal_4855, signal_3793}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_527 ( .clk (signal_6181), .D ({signal_5547, signal_577}), .Q ({signal_4858, signal_3792}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_530 ( .clk (signal_6181), .D ({signal_5549, signal_579}), .Q ({signal_4861, signal_3791}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_533 ( .clk (signal_6181), .D ({signal_5551, signal_581}), .Q ({signal_4867, signal_3790}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_536 ( .clk (signal_6181), .D ({signal_5553, signal_583}), .Q ({signal_4870, signal_3789}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_539 ( .clk (signal_6181), .D ({signal_5555, signal_585}), .Q ({signal_4873, signal_3788}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_542 ( .clk (signal_6181), .D ({signal_5557, signal_587}), .Q ({signal_4876, signal_3787}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_545 ( .clk (signal_6181), .D ({signal_5559, signal_589}), .Q ({signal_4879, signal_3786}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_548 ( .clk (signal_6181), .D ({signal_5561, signal_591}), .Q ({signal_4882, signal_3785}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_551 ( .clk (signal_6181), .D ({signal_5563, signal_593}), .Q ({signal_4885, signal_3784}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_554 ( .clk (signal_6181), .D ({signal_5565, signal_595}), .Q ({signal_4888, signal_3783}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_557 ( .clk (signal_6181), .D ({signal_5567, signal_597}), .Q ({signal_4891, signal_3782}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_560 ( .clk (signal_6181), .D ({signal_5569, signal_599}), .Q ({signal_4894, signal_3781}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_563 ( .clk (signal_6181), .D ({signal_5571, signal_601}), .Q ({signal_4900, signal_3780}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_566 ( .clk (signal_6181), .D ({signal_5573, signal_603}), .Q ({signal_4903, signal_3779}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_569 ( .clk (signal_6181), .D ({signal_5575, signal_605}), .Q ({signal_4906, signal_3778}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_572 ( .clk (signal_6181), .D ({signal_5577, signal_607}), .Q ({signal_4909, signal_3777}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_575 ( .clk (signal_6181), .D ({signal_5579, signal_609}), .Q ({signal_4912, signal_3776}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_578 ( .clk (signal_6181), .D ({signal_5581, signal_611}), .Q ({signal_4915, signal_3775}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_581 ( .clk (signal_6181), .D ({signal_5735, signal_613}), .Q ({signal_4918, signal_3774}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_584 ( .clk (signal_6181), .D ({signal_5583, signal_615}), .Q ({signal_4921, signal_3773}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_587 ( .clk (signal_6181), .D ({signal_5585, signal_617}), .Q ({signal_4924, signal_3772}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_590 ( .clk (signal_6181), .D ({signal_5587, signal_619}), .Q ({signal_4927, signal_3771}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_593 ( .clk (signal_6181), .D ({signal_5589, signal_621}), .Q ({signal_4552, signal_3770}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_596 ( .clk (signal_6181), .D ({signal_5591, signal_623}), .Q ({signal_4555, signal_3769}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_599 ( .clk (signal_6181), .D ({signal_5593, signal_625}), .Q ({signal_4558, signal_3768}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_602 ( .clk (signal_6181), .D ({signal_5595, signal_627}), .Q ({signal_4561, signal_3767}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_605 ( .clk (signal_6181), .D ({signal_5597, signal_629}), .Q ({signal_4564, signal_3766}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_608 ( .clk (signal_6181), .D ({signal_5737, signal_631}), .Q ({signal_4567, signal_3765}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_611 ( .clk (signal_6181), .D ({signal_5599, signal_633}), .Q ({signal_4570, signal_3764}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_614 ( .clk (signal_6181), .D ({signal_5601, signal_635}), .Q ({signal_4573, signal_3763}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_617 ( .clk (signal_6181), .D ({signal_5603, signal_637}), .Q ({signal_4576, signal_3762}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_620 ( .clk (signal_6181), .D ({signal_5605, signal_639}), .Q ({signal_4579, signal_3761}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_623 ( .clk (signal_6181), .D ({signal_5607, signal_641}), .Q ({signal_4585, signal_3760}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_626 ( .clk (signal_6181), .D ({signal_5609, signal_643}), .Q ({signal_4588, signal_3759}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_629 ( .clk (signal_6181), .D ({signal_5611, signal_645}), .Q ({signal_4591, signal_3758}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_632 ( .clk (signal_6181), .D ({signal_5613, signal_647}), .Q ({signal_4594, signal_3757}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_635 ( .clk (signal_6181), .D ({signal_5615, signal_649}), .Q ({signal_4597, signal_3756}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_638 ( .clk (signal_6181), .D ({signal_5617, signal_651}), .Q ({signal_4600, signal_3755}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_641 ( .clk (signal_6181), .D ({signal_5619, signal_653}), .Q ({signal_4603, signal_3754}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_644 ( .clk (signal_6181), .D ({signal_5621, signal_655}), .Q ({signal_4606, signal_3753}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_647 ( .clk (signal_6181), .D ({signal_5623, signal_657}), .Q ({signal_4609, signal_3752}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_650 ( .clk (signal_6181), .D ({signal_5625, signal_659}), .Q ({signal_4612, signal_3751}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_653 ( .clk (signal_6181), .D ({signal_5627, signal_661}), .Q ({signal_4618, signal_3750}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_656 ( .clk (signal_6181), .D ({signal_5629, signal_663}), .Q ({signal_4621, signal_3749}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_659 ( .clk (signal_6181), .D ({signal_5631, signal_665}), .Q ({signal_4624, signal_3748}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_662 ( .clk (signal_6181), .D ({signal_5633, signal_667}), .Q ({signal_4627, signal_3747}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_665 ( .clk (signal_6181), .D ({signal_5635, signal_669}), .Q ({signal_4630, signal_3746}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_668 ( .clk (signal_6181), .D ({signal_5637, signal_671}), .Q ({signal_4633, signal_3745}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_671 ( .clk (signal_6181), .D ({signal_5639, signal_673}), .Q ({signal_4636, signal_3744}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_674 ( .clk (signal_6181), .D ({signal_5641, signal_675}), .Q ({signal_4639, signal_3743}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3157 ( .clk (signal_6181), .D ({signal_5925, signal_2853}), .Q ({signal_4550, signal_4378}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3160 ( .clk (signal_6181), .D ({signal_5927, signal_2855}), .Q ({signal_4667, signal_4377}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3163 ( .clk (signal_6181), .D ({signal_5929, signal_2857}), .Q ({signal_4700, signal_4376}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3166 ( .clk (signal_6181), .D ({signal_5931, signal_2859}), .Q ({signal_4733, signal_4375}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3169 ( .clk (signal_6181), .D ({signal_5933, signal_2861}), .Q ({signal_4766, signal_4374}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3172 ( .clk (signal_6181), .D ({signal_5935, signal_2863}), .Q ({signal_4799, signal_4373}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3175 ( .clk (signal_6181), .D ({signal_5937, signal_2865}), .Q ({signal_4832, signal_4372}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3178 ( .clk (signal_6181), .D ({signal_5939, signal_2867}), .Q ({signal_4865, signal_4371}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3181 ( .clk (signal_6181), .D ({signal_5941, signal_2869}), .Q ({signal_4898, signal_4370}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3184 ( .clk (signal_6181), .D ({signal_5943, signal_2871}), .Q ({signal_4931, signal_4369}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3187 ( .clk (signal_6181), .D ({signal_5945, signal_2873}), .Q ({signal_4583, signal_4368}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3190 ( .clk (signal_6181), .D ({signal_5947, signal_2875}), .Q ({signal_4616, signal_4367}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3193 ( .clk (signal_6181), .D ({signal_5949, signal_2877}), .Q ({signal_4643, signal_4366}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3196 ( .clk (signal_6181), .D ({signal_5951, signal_2879}), .Q ({signal_4646, signal_4365}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3199 ( .clk (signal_6181), .D ({signal_5953, signal_2881}), .Q ({signal_4649, signal_4364}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3202 ( .clk (signal_6181), .D ({signal_5955, signal_2883}), .Q ({signal_4652, signal_4363}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3205 ( .clk (signal_6181), .D ({signal_5957, signal_2885}), .Q ({signal_4655, signal_4362}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3208 ( .clk (signal_6181), .D ({signal_5959, signal_2887}), .Q ({signal_4658, signal_4361}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3211 ( .clk (signal_6181), .D ({signal_5961, signal_2889}), .Q ({signal_4661, signal_4360}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3214 ( .clk (signal_6181), .D ({signal_5963, signal_2891}), .Q ({signal_4664, signal_4359}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3217 ( .clk (signal_6181), .D ({signal_5965, signal_2893}), .Q ({signal_4670, signal_4358}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3220 ( .clk (signal_6181), .D ({signal_5967, signal_2895}), .Q ({signal_4673, signal_4357}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3223 ( .clk (signal_6181), .D ({signal_5969, signal_2897}), .Q ({signal_4676, signal_4356}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3226 ( .clk (signal_6181), .D ({signal_5971, signal_2899}), .Q ({signal_4679, signal_4355}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3229 ( .clk (signal_6181), .D ({signal_5997, signal_2901}), .Q ({signal_4682, signal_4354}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3232 ( .clk (signal_6181), .D ({signal_5999, signal_2903}), .Q ({signal_4685, signal_4353}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3235 ( .clk (signal_6181), .D ({signal_6016, signal_2905}), .Q ({signal_4688, signal_4352}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3238 ( .clk (signal_6181), .D ({signal_6018, signal_2907}), .Q ({signal_4691, signal_4351}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3241 ( .clk (signal_6181), .D ({signal_6001, signal_2909}), .Q ({signal_4694, signal_4350}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3244 ( .clk (signal_6181), .D ({signal_6020, signal_2911}), .Q ({signal_4697, signal_4349}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3247 ( .clk (signal_6181), .D ({signal_6003, signal_2913}), .Q ({signal_4703, signal_4348}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3250 ( .clk (signal_6181), .D ({signal_6005, signal_2915}), .Q ({signal_4706, signal_4347}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3253 ( .clk (signal_6181), .D ({signal_5829, signal_2917}), .Q ({signal_4709, signal_4346}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3256 ( .clk (signal_6181), .D ({signal_5831, signal_2919}), .Q ({signal_4712, signal_4345}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3259 ( .clk (signal_6181), .D ({signal_5833, signal_2921}), .Q ({signal_4715, signal_4344}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3262 ( .clk (signal_6181), .D ({signal_5835, signal_2923}), .Q ({signal_4718, signal_4343}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3265 ( .clk (signal_6181), .D ({signal_5837, signal_2925}), .Q ({signal_4721, signal_4342}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3268 ( .clk (signal_6181), .D ({signal_5839, signal_2927}), .Q ({signal_4724, signal_4341}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3271 ( .clk (signal_6181), .D ({signal_5841, signal_2929}), .Q ({signal_4727, signal_4340}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3274 ( .clk (signal_6181), .D ({signal_5843, signal_2931}), .Q ({signal_4730, signal_4339}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3277 ( .clk (signal_6181), .D ({signal_5845, signal_2933}), .Q ({signal_4736, signal_4338}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3280 ( .clk (signal_6181), .D ({signal_5847, signal_2935}), .Q ({signal_4739, signal_4337}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3283 ( .clk (signal_6181), .D ({signal_5849, signal_2937}), .Q ({signal_4742, signal_4336}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3286 ( .clk (signal_6181), .D ({signal_5851, signal_2939}), .Q ({signal_4745, signal_4335}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3289 ( .clk (signal_6181), .D ({signal_5853, signal_2941}), .Q ({signal_4748, signal_4334}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3292 ( .clk (signal_6181), .D ({signal_5855, signal_2943}), .Q ({signal_4751, signal_4333}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3295 ( .clk (signal_6181), .D ({signal_5857, signal_2945}), .Q ({signal_4754, signal_4332}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3298 ( .clk (signal_6181), .D ({signal_5859, signal_2947}), .Q ({signal_4757, signal_4331}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3301 ( .clk (signal_6181), .D ({signal_5861, signal_2949}), .Q ({signal_4760, signal_4330}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3304 ( .clk (signal_6181), .D ({signal_5863, signal_2951}), .Q ({signal_4763, signal_4329}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3307 ( .clk (signal_6181), .D ({signal_5865, signal_2953}), .Q ({signal_4769, signal_4328}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3310 ( .clk (signal_6181), .D ({signal_5867, signal_2955}), .Q ({signal_4772, signal_4327}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3313 ( .clk (signal_6181), .D ({signal_5869, signal_2957}), .Q ({signal_4775, signal_4326}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3316 ( .clk (signal_6181), .D ({signal_5871, signal_2959}), .Q ({signal_4778, signal_4325}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3319 ( .clk (signal_6181), .D ({signal_5873, signal_2961}), .Q ({signal_4781, signal_4324}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3322 ( .clk (signal_6181), .D ({signal_5875, signal_2963}), .Q ({signal_4784, signal_4323}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3325 ( .clk (signal_6181), .D ({signal_5973, signal_2965}), .Q ({signal_4787, signal_4322}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3328 ( .clk (signal_6181), .D ({signal_5975, signal_2967}), .Q ({signal_4790, signal_4321}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3331 ( .clk (signal_6181), .D ({signal_6007, signal_2969}), .Q ({signal_4793, signal_4320}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3334 ( .clk (signal_6181), .D ({signal_6009, signal_2971}), .Q ({signal_4796, signal_4319}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3337 ( .clk (signal_6181), .D ({signal_5977, signal_2973}), .Q ({signal_4802, signal_4318}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3340 ( .clk (signal_6181), .D ({signal_6011, signal_2975}), .Q ({signal_4805, signal_4317}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3343 ( .clk (signal_6181), .D ({signal_5979, signal_2977}), .Q ({signal_4808, signal_4316}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3346 ( .clk (signal_6181), .D ({signal_5981, signal_2979}), .Q ({signal_4811, signal_4315}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3349 ( .clk (signal_6181), .D ({signal_5739, signal_2981}), .Q ({signal_4814, signal_4314}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3352 ( .clk (signal_6181), .D ({signal_5741, signal_2983}), .Q ({signal_4817, signal_4313}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3355 ( .clk (signal_6181), .D ({signal_5743, signal_2985}), .Q ({signal_4820, signal_4312}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3358 ( .clk (signal_6181), .D ({signal_5745, signal_2987}), .Q ({signal_4823, signal_4311}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3361 ( .clk (signal_6181), .D ({signal_5747, signal_2989}), .Q ({signal_4826, signal_4310}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3364 ( .clk (signal_6181), .D ({signal_5749, signal_2991}), .Q ({signal_4829, signal_4309}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3367 ( .clk (signal_6181), .D ({signal_5751, signal_2993}), .Q ({signal_4835, signal_4308}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3370 ( .clk (signal_6181), .D ({signal_5753, signal_2995}), .Q ({signal_4838, signal_4307}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3373 ( .clk (signal_6181), .D ({signal_5755, signal_2997}), .Q ({signal_4841, signal_4306}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3376 ( .clk (signal_6181), .D ({signal_5757, signal_2999}), .Q ({signal_4844, signal_4305}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3379 ( .clk (signal_6181), .D ({signal_5759, signal_3001}), .Q ({signal_4847, signal_4304}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3382 ( .clk (signal_6181), .D ({signal_5761, signal_3003}), .Q ({signal_4850, signal_4303}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3385 ( .clk (signal_6181), .D ({signal_5763, signal_3005}), .Q ({signal_4853, signal_4302}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3388 ( .clk (signal_6181), .D ({signal_5765, signal_3007}), .Q ({signal_4856, signal_4301}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3391 ( .clk (signal_6181), .D ({signal_5767, signal_3009}), .Q ({signal_4859, signal_4300}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3394 ( .clk (signal_6181), .D ({signal_5769, signal_3011}), .Q ({signal_4862, signal_4299}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3397 ( .clk (signal_6181), .D ({signal_5771, signal_3013}), .Q ({signal_4868, signal_4298}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3400 ( .clk (signal_6181), .D ({signal_5773, signal_3015}), .Q ({signal_4871, signal_4297}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3403 ( .clk (signal_6181), .D ({signal_5775, signal_3017}), .Q ({signal_4874, signal_4296}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3406 ( .clk (signal_6181), .D ({signal_5777, signal_3019}), .Q ({signal_4877, signal_4295}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3409 ( .clk (signal_6181), .D ({signal_5779, signal_3021}), .Q ({signal_4880, signal_4294}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3412 ( .clk (signal_6181), .D ({signal_5781, signal_3023}), .Q ({signal_4883, signal_4293}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3415 ( .clk (signal_6181), .D ({signal_5783, signal_3025}), .Q ({signal_4886, signal_4292}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3418 ( .clk (signal_6181), .D ({signal_5785, signal_3027}), .Q ({signal_4889, signal_4291}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3421 ( .clk (signal_6181), .D ({signal_5877, signal_3029}), .Q ({signal_4892, signal_4290}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3424 ( .clk (signal_6181), .D ({signal_5879, signal_3031}), .Q ({signal_4895, signal_4289}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3427 ( .clk (signal_6181), .D ({signal_5983, signal_3033}), .Q ({signal_4901, signal_4288}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3430 ( .clk (signal_6181), .D ({signal_5985, signal_3035}), .Q ({signal_4904, signal_4287}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3433 ( .clk (signal_6181), .D ({signal_5881, signal_3037}), .Q ({signal_4907, signal_4286}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3436 ( .clk (signal_6181), .D ({signal_5987, signal_3039}), .Q ({signal_4910, signal_4285}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3439 ( .clk (signal_6181), .D ({signal_5883, signal_3041}), .Q ({signal_4913, signal_4284}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3442 ( .clk (signal_6181), .D ({signal_5885, signal_3043}), .Q ({signal_4916, signal_4283}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3445 ( .clk (signal_6181), .D ({signal_5643, signal_3045}), .Q ({signal_4919, signal_4282}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3448 ( .clk (signal_6181), .D ({signal_5645, signal_3047}), .Q ({signal_4922, signal_4281}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3451 ( .clk (signal_6181), .D ({signal_5647, signal_3049}), .Q ({signal_4925, signal_4280}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3454 ( .clk (signal_6181), .D ({signal_5649, signal_3051}), .Q ({signal_4928, signal_4279}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3457 ( .clk (signal_6181), .D ({signal_5651, signal_3053}), .Q ({signal_4553, signal_4278}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3460 ( .clk (signal_6181), .D ({signal_5653, signal_3055}), .Q ({signal_4556, signal_4277}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3463 ( .clk (signal_6181), .D ({signal_5655, signal_3057}), .Q ({signal_4559, signal_4276}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3466 ( .clk (signal_6181), .D ({signal_5657, signal_3059}), .Q ({signal_4562, signal_4275}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3469 ( .clk (signal_6181), .D ({signal_5659, signal_3061}), .Q ({signal_4565, signal_4274}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3472 ( .clk (signal_6181), .D ({signal_5661, signal_3063}), .Q ({signal_4568, signal_4273}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3475 ( .clk (signal_6181), .D ({signal_5663, signal_3065}), .Q ({signal_4571, signal_4272}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3478 ( .clk (signal_6181), .D ({signal_5665, signal_3067}), .Q ({signal_4574, signal_4271}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3481 ( .clk (signal_6181), .D ({signal_5667, signal_3069}), .Q ({signal_4577, signal_4270}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3484 ( .clk (signal_6181), .D ({signal_5669, signal_3071}), .Q ({signal_4580, signal_4269}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3487 ( .clk (signal_6181), .D ({signal_5671, signal_3073}), .Q ({signal_4586, signal_4268}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3490 ( .clk (signal_6181), .D ({signal_5673, signal_3075}), .Q ({signal_4589, signal_4267}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3493 ( .clk (signal_6181), .D ({signal_5675, signal_3077}), .Q ({signal_4592, signal_4266}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3496 ( .clk (signal_6181), .D ({signal_5677, signal_3079}), .Q ({signal_4595, signal_4265}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3499 ( .clk (signal_6181), .D ({signal_5679, signal_3081}), .Q ({signal_4598, signal_4264}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3502 ( .clk (signal_6181), .D ({signal_5681, signal_3083}), .Q ({signal_4601, signal_4263}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3505 ( .clk (signal_6181), .D ({signal_5683, signal_3085}), .Q ({signal_4604, signal_4262}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3508 ( .clk (signal_6181), .D ({signal_5685, signal_3087}), .Q ({signal_4607, signal_4261}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3511 ( .clk (signal_6181), .D ({signal_5687, signal_3089}), .Q ({signal_4610, signal_4260}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3514 ( .clk (signal_6181), .D ({signal_5689, signal_3091}), .Q ({signal_4613, signal_4259}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3517 ( .clk (signal_6181), .D ({signal_5787, signal_3093}), .Q ({signal_4619, signal_4258}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3520 ( .clk (signal_6181), .D ({signal_5789, signal_3095}), .Q ({signal_4622, signal_4257}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3523 ( .clk (signal_6181), .D ({signal_5887, signal_3097}), .Q ({signal_4625, signal_4256}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3526 ( .clk (signal_6181), .D ({signal_5889, signal_3099}), .Q ({signal_4628, signal_4255}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3529 ( .clk (signal_6181), .D ({signal_5791, signal_3101}), .Q ({signal_4631, signal_4254}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3532 ( .clk (signal_6181), .D ({signal_5891, signal_3103}), .Q ({signal_4634, signal_4253}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3535 ( .clk (signal_6181), .D ({signal_5793, signal_3105}), .Q ({signal_4637, signal_4252}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_3538 ( .clk (signal_6181), .D ({signal_5795, signal_3107}), .Q ({signal_4640, signal_4251}) ) ;
    DFF_X1 cell_4202 ( .CK (signal_6181), .D (signal_3612), .Q (signal_4388), .QN () ) ;
    DFF_X1 cell_4204 ( .CK (signal_6181), .D (signal_3610), .Q (signal_4387), .QN () ) ;
    DFF_X1 cell_4206 ( .CK (signal_6181), .D (signal_3607), .Q (signal_4386), .QN () ) ;
    DFF_X1 cell_4208 ( .CK (signal_6181), .D (signal_3608), .Q (signal_4385), .QN () ) ;
endmodule
