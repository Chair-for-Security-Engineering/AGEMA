/* modified netlist. Source: module sbox in file ../sbox_lookup/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC2_BDDcudd_Pipeline_d3 (SI_s0, clk, SI_s1, SI_s2, SI_s3, Fresh, SO_s0, SO_s1, SO_s2, SO_s3);
    input [3:0] SI_s0 ;
    input clk ;
    input [3:0] SI_s1 ;
    input [3:0] SI_s2 ;
    input [3:0] SI_s3 ;
    input [101:0] Fresh ;
    output [3:0] SO_s0 ;
    output [3:0] SO_s1 ;
    output [3:0] SO_s2 ;
    output [3:0] SO_s3 ;
    wire signal_15 ;
    wire signal_16 ;
    wire signal_17 ;
    wire signal_18 ;
    wire signal_34 ;
    wire signal_35 ;
    wire signal_36 ;
    wire signal_37 ;
    wire signal_38 ;
    wire signal_39 ;
    wire signal_40 ;
    wire signal_41 ;
    wire signal_42 ;
    wire signal_43 ;
    wire signal_44 ;
    wire signal_45 ;
    wire signal_46 ;
    wire signal_50 ;
    wire signal_51 ;
    wire signal_52 ;
    wire signal_53 ;
    wire signal_54 ;
    wire signal_55 ;
    wire signal_59 ;
    wire signal_60 ;
    wire signal_61 ;
    wire signal_62 ;
    wire signal_63 ;
    wire signal_64 ;
    wire signal_65 ;
    wire signal_66 ;
    wire signal_67 ;
    wire signal_68 ;
    wire signal_69 ;
    wire signal_70 ;
    wire signal_71 ;
    wire signal_72 ;
    wire signal_73 ;
    wire signal_74 ;
    wire signal_75 ;
    wire signal_76 ;
    wire signal_77 ;
    wire signal_78 ;
    wire signal_79 ;
    wire signal_80 ;
    wire signal_81 ;
    wire signal_82 ;
    wire signal_86 ;
    wire signal_87 ;
    wire signal_88 ;
    wire signal_89 ;
    wire signal_90 ;
    wire signal_91 ;
    wire signal_92 ;
    wire signal_93 ;
    wire signal_94 ;
    wire signal_98 ;
    wire signal_99 ;
    wire signal_100 ;
    wire signal_101 ;
    wire signal_102 ;
    wire signal_103 ;
    wire signal_104 ;
    wire signal_105 ;
    wire signal_106 ;
    wire signal_107 ;
    wire signal_108 ;
    wire signal_109 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;

    /* cells in depth 0 */

    /* cells in depth 1 */
    buf_clk cell_40 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( signal_224 ) ) ;
    buf_clk cell_42 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( signal_226 ) ) ;
    buf_clk cell_44 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( signal_228 ) ) ;
    buf_clk cell_46 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( signal_230 ) ) ;
    buf_clk cell_48 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( signal_232 ) ) ;
    buf_clk cell_52 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( signal_236 ) ) ;
    buf_clk cell_56 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( signal_240 ) ) ;
    buf_clk cell_60 ( .C ( clk ), .D ( SI_s3[0] ), .Q ( signal_244 ) ) ;
    buf_clk cell_64 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( signal_248 ) ) ;
    buf_clk cell_68 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( signal_252 ) ) ;
    buf_clk cell_72 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( signal_256 ) ) ;
    buf_clk cell_76 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( signal_260 ) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_23 ( .s ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_52, signal_51, signal_50, signal_34}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_24 ( .s ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_55, signal_54, signal_53, signal_35}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_25 ( .s ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_61, signal_60, signal_59, signal_36}) ) ;
    buf_clk cell_41 ( .C ( clk ), .D ( signal_224 ), .Q ( signal_225 ) ) ;
    buf_clk cell_43 ( .C ( clk ), .D ( signal_226 ), .Q ( signal_227 ) ) ;
    buf_clk cell_45 ( .C ( clk ), .D ( signal_228 ), .Q ( signal_229 ) ) ;
    buf_clk cell_47 ( .C ( clk ), .D ( signal_230 ), .Q ( signal_231 ) ) ;
    buf_clk cell_49 ( .C ( clk ), .D ( signal_232 ), .Q ( signal_233 ) ) ;
    buf_clk cell_53 ( .C ( clk ), .D ( signal_236 ), .Q ( signal_237 ) ) ;
    buf_clk cell_57 ( .C ( clk ), .D ( signal_240 ), .Q ( signal_241 ) ) ;
    buf_clk cell_61 ( .C ( clk ), .D ( signal_244 ), .Q ( signal_245 ) ) ;
    buf_clk cell_65 ( .C ( clk ), .D ( signal_248 ), .Q ( signal_249 ) ) ;
    buf_clk cell_69 ( .C ( clk ), .D ( signal_252 ), .Q ( signal_253 ) ) ;
    buf_clk cell_73 ( .C ( clk ), .D ( signal_256 ), .Q ( signal_257 ) ) ;
    buf_clk cell_77 ( .C ( clk ), .D ( signal_260 ), .Q ( signal_261 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_50 ( .C ( clk ), .D ( signal_233 ), .Q ( signal_234 ) ) ;
    buf_clk cell_54 ( .C ( clk ), .D ( signal_237 ), .Q ( signal_238 ) ) ;
    buf_clk cell_58 ( .C ( clk ), .D ( signal_241 ), .Q ( signal_242 ) ) ;
    buf_clk cell_62 ( .C ( clk ), .D ( signal_245 ), .Q ( signal_246 ) ) ;
    buf_clk cell_66 ( .C ( clk ), .D ( signal_249 ), .Q ( signal_250 ) ) ;
    buf_clk cell_70 ( .C ( clk ), .D ( signal_253 ), .Q ( signal_254 ) ) ;
    buf_clk cell_74 ( .C ( clk ), .D ( signal_257 ), .Q ( signal_258 ) ) ;
    buf_clk cell_78 ( .C ( clk ), .D ( signal_261 ), .Q ( signal_262 ) ) ;
    buf_clk cell_80 ( .C ( clk ), .D ( signal_35 ), .Q ( signal_264 ) ) ;
    buf_clk cell_82 ( .C ( clk ), .D ( signal_53 ), .Q ( signal_266 ) ) ;
    buf_clk cell_84 ( .C ( clk ), .D ( signal_54 ), .Q ( signal_268 ) ) ;
    buf_clk cell_86 ( .C ( clk ), .D ( signal_55 ), .Q ( signal_270 ) ) ;
    buf_clk cell_96 ( .C ( clk ), .D ( signal_36 ), .Q ( signal_280 ) ) ;
    buf_clk cell_100 ( .C ( clk ), .D ( signal_59 ), .Q ( signal_284 ) ) ;
    buf_clk cell_104 ( .C ( clk ), .D ( signal_60 ), .Q ( signal_288 ) ) ;
    buf_clk cell_108 ( .C ( clk ), .D ( signal_61 ), .Q ( signal_292 ) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_26 ( .s ({signal_231, signal_229, signal_227, signal_225}), .b ({signal_52, signal_51, signal_50, signal_34}), .a ({signal_55, signal_54, signal_53, signal_35}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_64, signal_63, signal_62, signal_37}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_27 ( .s ({signal_231, signal_229, signal_227, signal_225}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_55, signal_54, signal_53, signal_35}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_67, signal_66, signal_65, signal_38}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_28 ( .s ({signal_231, signal_229, signal_227, signal_225}), .b ({signal_52, signal_51, signal_50, signal_34}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_70, signal_69, signal_68, signal_39}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_29 ( .s ({signal_231, signal_229, signal_227, signal_225}), .b ({signal_55, signal_54, signal_53, signal_35}), .a ({signal_52, signal_51, signal_50, signal_34}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_73, signal_72, signal_71, signal_40}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_30 ( .s ({signal_231, signal_229, signal_227, signal_225}), .b ({signal_55, signal_54, signal_53, signal_35}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_76, signal_75, signal_74, signal_41}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_31 ( .s ({signal_231, signal_229, signal_227, signal_225}), .b ({signal_55, signal_54, signal_53, signal_35}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_79, signal_78, signal_77, signal_42}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_32 ( .s ({signal_231, signal_229, signal_227, signal_225}), .b ({signal_52, signal_51, signal_50, signal_34}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_82, signal_81, signal_80, signal_43}) ) ;
    buf_clk cell_51 ( .C ( clk ), .D ( signal_234 ), .Q ( signal_235 ) ) ;
    buf_clk cell_55 ( .C ( clk ), .D ( signal_238 ), .Q ( signal_239 ) ) ;
    buf_clk cell_59 ( .C ( clk ), .D ( signal_242 ), .Q ( signal_243 ) ) ;
    buf_clk cell_63 ( .C ( clk ), .D ( signal_246 ), .Q ( signal_247 ) ) ;
    buf_clk cell_67 ( .C ( clk ), .D ( signal_250 ), .Q ( signal_251 ) ) ;
    buf_clk cell_71 ( .C ( clk ), .D ( signal_254 ), .Q ( signal_255 ) ) ;
    buf_clk cell_75 ( .C ( clk ), .D ( signal_258 ), .Q ( signal_259 ) ) ;
    buf_clk cell_79 ( .C ( clk ), .D ( signal_262 ), .Q ( signal_263 ) ) ;
    buf_clk cell_81 ( .C ( clk ), .D ( signal_264 ), .Q ( signal_265 ) ) ;
    buf_clk cell_83 ( .C ( clk ), .D ( signal_266 ), .Q ( signal_267 ) ) ;
    buf_clk cell_85 ( .C ( clk ), .D ( signal_268 ), .Q ( signal_269 ) ) ;
    buf_clk cell_87 ( .C ( clk ), .D ( signal_270 ), .Q ( signal_271 ) ) ;
    buf_clk cell_97 ( .C ( clk ), .D ( signal_280 ), .Q ( signal_281 ) ) ;
    buf_clk cell_101 ( .C ( clk ), .D ( signal_284 ), .Q ( signal_285 ) ) ;
    buf_clk cell_105 ( .C ( clk ), .D ( signal_288 ), .Q ( signal_289 ) ) ;
    buf_clk cell_109 ( .C ( clk ), .D ( signal_292 ), .Q ( signal_293 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_88 ( .C ( clk ), .D ( signal_251 ), .Q ( signal_272 ) ) ;
    buf_clk cell_90 ( .C ( clk ), .D ( signal_255 ), .Q ( signal_274 ) ) ;
    buf_clk cell_92 ( .C ( clk ), .D ( signal_259 ), .Q ( signal_276 ) ) ;
    buf_clk cell_94 ( .C ( clk ), .D ( signal_263 ), .Q ( signal_278 ) ) ;
    buf_clk cell_98 ( .C ( clk ), .D ( signal_281 ), .Q ( signal_282 ) ) ;
    buf_clk cell_102 ( .C ( clk ), .D ( signal_285 ), .Q ( signal_286 ) ) ;
    buf_clk cell_106 ( .C ( clk ), .D ( signal_289 ), .Q ( signal_290 ) ) ;
    buf_clk cell_110 ( .C ( clk ), .D ( signal_293 ), .Q ( signal_294 ) ) ;

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_33 ( .s ({signal_247, signal_243, signal_239, signal_235}), .b ({signal_73, signal_72, signal_71, signal_40}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_88, signal_87, signal_86, signal_44}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_34 ( .s ({signal_247, signal_243, signal_239, signal_235}), .b ({signal_67, signal_66, signal_65, signal_38}), .a ({signal_76, signal_75, signal_74, signal_41}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_91, signal_90, signal_89, signal_45}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_35 ( .s ({signal_247, signal_243, signal_239, signal_235}), .b ({signal_79, signal_78, signal_77, signal_42}), .a ({signal_70, signal_69, signal_68, signal_39}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_94, signal_93, signal_92, signal_46}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_36 ( .s ({signal_263, signal_259, signal_255, signal_251}), .b ({signal_64, signal_63, signal_62, signal_37}), .a ({signal_271, signal_269, signal_267, signal_265}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_100, signal_99, signal_98, signal_16}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_37 ( .s ({signal_247, signal_243, signal_239, signal_235}), .b ({signal_82, signal_81, signal_80, signal_43}), .a ({signal_76, signal_75, signal_74, signal_41}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_103, signal_102, signal_101, signal_15}) ) ;
    buf_clk cell_89 ( .C ( clk ), .D ( signal_272 ), .Q ( signal_273 ) ) ;
    buf_clk cell_91 ( .C ( clk ), .D ( signal_274 ), .Q ( signal_275 ) ) ;
    buf_clk cell_93 ( .C ( clk ), .D ( signal_276 ), .Q ( signal_277 ) ) ;
    buf_clk cell_95 ( .C ( clk ), .D ( signal_278 ), .Q ( signal_279 ) ) ;
    buf_clk cell_99 ( .C ( clk ), .D ( signal_282 ), .Q ( signal_283 ) ) ;
    buf_clk cell_103 ( .C ( clk ), .D ( signal_286 ), .Q ( signal_287 ) ) ;
    buf_clk cell_107 ( .C ( clk ), .D ( signal_290 ), .Q ( signal_291 ) ) ;
    buf_clk cell_111 ( .C ( clk ), .D ( signal_294 ), .Q ( signal_295 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_112 ( .C ( clk ), .D ( signal_15 ), .Q ( signal_296 ) ) ;
    buf_clk cell_114 ( .C ( clk ), .D ( signal_101 ), .Q ( signal_298 ) ) ;
    buf_clk cell_116 ( .C ( clk ), .D ( signal_102 ), .Q ( signal_300 ) ) ;
    buf_clk cell_118 ( .C ( clk ), .D ( signal_103 ), .Q ( signal_302 ) ) ;
    buf_clk cell_120 ( .C ( clk ), .D ( signal_16 ), .Q ( signal_304 ) ) ;
    buf_clk cell_122 ( .C ( clk ), .D ( signal_98 ), .Q ( signal_306 ) ) ;
    buf_clk cell_124 ( .C ( clk ), .D ( signal_99 ), .Q ( signal_308 ) ) ;
    buf_clk cell_126 ( .C ( clk ), .D ( signal_100 ), .Q ( signal_310 ) ) ;

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_38 ( .s ({signal_279, signal_277, signal_275, signal_273}), .b ({signal_88, signal_87, signal_86, signal_44}), .a ({signal_91, signal_90, signal_89, signal_45}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_106, signal_105, signal_104, signal_18}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_39 ( .s ({signal_279, signal_277, signal_275, signal_273}), .b ({signal_94, signal_93, signal_92, signal_46}), .a ({signal_295, signal_291, signal_287, signal_283}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_109, signal_108, signal_107, signal_17}) ) ;
    buf_clk cell_113 ( .C ( clk ), .D ( signal_296 ), .Q ( signal_297 ) ) ;
    buf_clk cell_115 ( .C ( clk ), .D ( signal_298 ), .Q ( signal_299 ) ) ;
    buf_clk cell_117 ( .C ( clk ), .D ( signal_300 ), .Q ( signal_301 ) ) ;
    buf_clk cell_119 ( .C ( clk ), .D ( signal_302 ), .Q ( signal_303 ) ) ;
    buf_clk cell_121 ( .C ( clk ), .D ( signal_304 ), .Q ( signal_305 ) ) ;
    buf_clk cell_123 ( .C ( clk ), .D ( signal_306 ), .Q ( signal_307 ) ) ;
    buf_clk cell_125 ( .C ( clk ), .D ( signal_308 ), .Q ( signal_309 ) ) ;
    buf_clk cell_127 ( .C ( clk ), .D ( signal_310 ), .Q ( signal_311 ) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_303, signal_301, signal_299, signal_297}), .Q ({SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_311, signal_309, signal_307, signal_305}), .Q ({SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_109, signal_108, signal_107, signal_17}), .Q ({SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_106, signal_105, signal_104, signal_18}), .Q ({SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
