
module SkinnyTop_HPC2_Pipeline_d1 ( Plaintext_s0, Key_s0, clk, rst, Key_s1, 
        Plaintext_s1, Fresh, Ciphertext_s0, done, Ciphertext_s1 );
  input [63:0] Plaintext_s0;
  input [63:0] Key_s0;
  input [63:0] Key_s1;
  input [63:0] Plaintext_s1;
  input [63:0] Fresh;
  output [63:0] Ciphertext_s0;
  output [63:0] Ciphertext_s1;
  input clk, rst;
  output done;
  wire   SubCellInst_SboxInst_0_n3, new_AGEMA_signal_1167,
         SubCellInst_SboxInst_0_XX_1_, new_AGEMA_signal_1169,
         SubCellInst_SboxInst_0_XX_2_, new_AGEMA_signal_1453,
         SubCellInst_SboxInst_0_Q0, new_AGEMA_signal_1454,
         SubCellInst_SboxInst_0_Q1, new_AGEMA_signal_1455,
         SubCellInst_SboxInst_0_Q4, new_AGEMA_signal_1456,
         SubCellInst_SboxInst_0_Q6, new_AGEMA_signal_1550,
         SubCellInst_SboxInst_0_L1, new_AGEMA_signal_1457,
         SubCellInst_SboxInst_0_L2, SubCellInst_SboxInst_1_n3,
         new_AGEMA_signal_1173, SubCellInst_SboxInst_1_XX_1_,
         new_AGEMA_signal_1175, SubCellInst_SboxInst_1_XX_2_,
         new_AGEMA_signal_1459, SubCellInst_SboxInst_1_Q0,
         new_AGEMA_signal_1460, SubCellInst_SboxInst_1_Q1,
         new_AGEMA_signal_1461, SubCellInst_SboxInst_1_Q4,
         new_AGEMA_signal_1462, SubCellInst_SboxInst_1_Q6,
         new_AGEMA_signal_1553, SubCellInst_SboxInst_1_L1,
         new_AGEMA_signal_1463, SubCellInst_SboxInst_1_L2,
         SubCellInst_SboxInst_2_n3, new_AGEMA_signal_1179,
         SubCellInst_SboxInst_2_XX_1_, new_AGEMA_signal_1181,
         SubCellInst_SboxInst_2_XX_2_, new_AGEMA_signal_1465,
         SubCellInst_SboxInst_2_Q0, new_AGEMA_signal_1466,
         SubCellInst_SboxInst_2_Q1, new_AGEMA_signal_1467,
         SubCellInst_SboxInst_2_Q4, new_AGEMA_signal_1468,
         SubCellInst_SboxInst_2_Q6, new_AGEMA_signal_1556,
         SubCellInst_SboxInst_2_L1, new_AGEMA_signal_1469,
         SubCellInst_SboxInst_2_L2, SubCellInst_SboxInst_3_n3,
         new_AGEMA_signal_1185, SubCellInst_SboxInst_3_XX_1_,
         new_AGEMA_signal_1187, SubCellInst_SboxInst_3_XX_2_,
         new_AGEMA_signal_1471, SubCellInst_SboxInst_3_Q0,
         new_AGEMA_signal_1472, SubCellInst_SboxInst_3_Q1,
         new_AGEMA_signal_1473, SubCellInst_SboxInst_3_Q4,
         new_AGEMA_signal_1474, SubCellInst_SboxInst_3_Q6,
         new_AGEMA_signal_1559, SubCellInst_SboxInst_3_L1,
         new_AGEMA_signal_1475, SubCellInst_SboxInst_3_L2,
         SubCellInst_SboxInst_4_n3, new_AGEMA_signal_1191,
         SubCellInst_SboxInst_4_XX_1_, new_AGEMA_signal_1193,
         SubCellInst_SboxInst_4_XX_2_, new_AGEMA_signal_1477,
         SubCellInst_SboxInst_4_Q0, new_AGEMA_signal_1478,
         SubCellInst_SboxInst_4_Q1, new_AGEMA_signal_1479,
         SubCellInst_SboxInst_4_Q4, new_AGEMA_signal_1480,
         SubCellInst_SboxInst_4_Q6, new_AGEMA_signal_1562,
         SubCellInst_SboxInst_4_L1, new_AGEMA_signal_1481,
         SubCellInst_SboxInst_4_L2, SubCellInst_SboxInst_5_n3,
         new_AGEMA_signal_1197, SubCellInst_SboxInst_5_XX_1_,
         new_AGEMA_signal_1199, SubCellInst_SboxInst_5_XX_2_,
         new_AGEMA_signal_1483, SubCellInst_SboxInst_5_Q0,
         new_AGEMA_signal_1484, SubCellInst_SboxInst_5_Q1,
         new_AGEMA_signal_1485, SubCellInst_SboxInst_5_Q4,
         new_AGEMA_signal_1486, SubCellInst_SboxInst_5_Q6,
         new_AGEMA_signal_1565, SubCellInst_SboxInst_5_L1,
         new_AGEMA_signal_1487, SubCellInst_SboxInst_5_L2,
         SubCellInst_SboxInst_6_n3, new_AGEMA_signal_1203,
         SubCellInst_SboxInst_6_XX_1_, new_AGEMA_signal_1205,
         SubCellInst_SboxInst_6_XX_2_, new_AGEMA_signal_1489,
         SubCellInst_SboxInst_6_Q0, new_AGEMA_signal_1490,
         SubCellInst_SboxInst_6_Q1, new_AGEMA_signal_1491,
         SubCellInst_SboxInst_6_Q4, new_AGEMA_signal_1492,
         SubCellInst_SboxInst_6_Q6, new_AGEMA_signal_1568,
         SubCellInst_SboxInst_6_L1, new_AGEMA_signal_1493,
         SubCellInst_SboxInst_6_L2, SubCellInst_SboxInst_7_n3,
         new_AGEMA_signal_1209, SubCellInst_SboxInst_7_XX_1_,
         new_AGEMA_signal_1211, SubCellInst_SboxInst_7_XX_2_,
         new_AGEMA_signal_1495, SubCellInst_SboxInst_7_Q0,
         new_AGEMA_signal_1496, SubCellInst_SboxInst_7_Q1,
         new_AGEMA_signal_1497, SubCellInst_SboxInst_7_Q4,
         new_AGEMA_signal_1498, SubCellInst_SboxInst_7_Q6,
         new_AGEMA_signal_1571, SubCellInst_SboxInst_7_L1,
         new_AGEMA_signal_1499, SubCellInst_SboxInst_7_L2,
         SubCellInst_SboxInst_8_n3, new_AGEMA_signal_1215,
         SubCellInst_SboxInst_8_XX_1_, new_AGEMA_signal_1217,
         SubCellInst_SboxInst_8_XX_2_, new_AGEMA_signal_1501,
         SubCellInst_SboxInst_8_Q0, new_AGEMA_signal_1502,
         SubCellInst_SboxInst_8_Q1, new_AGEMA_signal_1503,
         SubCellInst_SboxInst_8_Q4, new_AGEMA_signal_1504,
         SubCellInst_SboxInst_8_Q6, new_AGEMA_signal_1574,
         SubCellInst_SboxInst_8_L1, new_AGEMA_signal_1505,
         SubCellInst_SboxInst_8_L2, SubCellInst_SboxInst_9_n3,
         new_AGEMA_signal_1221, SubCellInst_SboxInst_9_XX_1_,
         new_AGEMA_signal_1223, SubCellInst_SboxInst_9_XX_2_,
         new_AGEMA_signal_1507, SubCellInst_SboxInst_9_Q0,
         new_AGEMA_signal_1508, SubCellInst_SboxInst_9_Q1,
         new_AGEMA_signal_1509, SubCellInst_SboxInst_9_Q4,
         new_AGEMA_signal_1510, SubCellInst_SboxInst_9_Q6,
         new_AGEMA_signal_1577, SubCellInst_SboxInst_9_L1,
         new_AGEMA_signal_1511, SubCellInst_SboxInst_9_L2,
         SubCellInst_SboxInst_10_n3, new_AGEMA_signal_1227,
         SubCellInst_SboxInst_10_XX_1_, new_AGEMA_signal_1229,
         SubCellInst_SboxInst_10_XX_2_, new_AGEMA_signal_1513,
         SubCellInst_SboxInst_10_Q0, new_AGEMA_signal_1514,
         SubCellInst_SboxInst_10_Q1, new_AGEMA_signal_1515,
         SubCellInst_SboxInst_10_Q4, new_AGEMA_signal_1516,
         SubCellInst_SboxInst_10_Q6, new_AGEMA_signal_1580,
         SubCellInst_SboxInst_10_L1, new_AGEMA_signal_1517,
         SubCellInst_SboxInst_10_L2, SubCellInst_SboxInst_11_n3,
         new_AGEMA_signal_1233, SubCellInst_SboxInst_11_XX_1_,
         new_AGEMA_signal_1235, SubCellInst_SboxInst_11_XX_2_,
         new_AGEMA_signal_1519, SubCellInst_SboxInst_11_Q0,
         new_AGEMA_signal_1520, SubCellInst_SboxInst_11_Q1,
         new_AGEMA_signal_1521, SubCellInst_SboxInst_11_Q4,
         new_AGEMA_signal_1522, SubCellInst_SboxInst_11_Q6,
         new_AGEMA_signal_1583, SubCellInst_SboxInst_11_L1,
         new_AGEMA_signal_1523, SubCellInst_SboxInst_11_L2,
         SubCellInst_SboxInst_12_n3, new_AGEMA_signal_1239,
         SubCellInst_SboxInst_12_XX_1_, new_AGEMA_signal_1241,
         SubCellInst_SboxInst_12_XX_2_, new_AGEMA_signal_1525,
         SubCellInst_SboxInst_12_Q0, new_AGEMA_signal_1526,
         SubCellInst_SboxInst_12_Q1, new_AGEMA_signal_1527,
         SubCellInst_SboxInst_12_Q4, new_AGEMA_signal_1528,
         SubCellInst_SboxInst_12_Q6, new_AGEMA_signal_1586,
         SubCellInst_SboxInst_12_L1, new_AGEMA_signal_1529,
         SubCellInst_SboxInst_12_L2, SubCellInst_SboxInst_13_n3,
         new_AGEMA_signal_1245, SubCellInst_SboxInst_13_XX_1_,
         new_AGEMA_signal_1247, SubCellInst_SboxInst_13_XX_2_,
         new_AGEMA_signal_1531, SubCellInst_SboxInst_13_Q0,
         new_AGEMA_signal_1532, SubCellInst_SboxInst_13_Q1,
         new_AGEMA_signal_1533, SubCellInst_SboxInst_13_Q4,
         new_AGEMA_signal_1534, SubCellInst_SboxInst_13_Q6,
         new_AGEMA_signal_1589, SubCellInst_SboxInst_13_L1,
         new_AGEMA_signal_1535, SubCellInst_SboxInst_13_L2,
         SubCellInst_SboxInst_14_n3, new_AGEMA_signal_1251,
         SubCellInst_SboxInst_14_XX_1_, new_AGEMA_signal_1253,
         SubCellInst_SboxInst_14_XX_2_, new_AGEMA_signal_1537,
         SubCellInst_SboxInst_14_Q0, new_AGEMA_signal_1538,
         SubCellInst_SboxInst_14_Q1, new_AGEMA_signal_1539,
         SubCellInst_SboxInst_14_Q4, new_AGEMA_signal_1540,
         SubCellInst_SboxInst_14_Q6, new_AGEMA_signal_1592,
         SubCellInst_SboxInst_14_L1, new_AGEMA_signal_1541,
         SubCellInst_SboxInst_14_L2, SubCellInst_SboxInst_15_n3,
         new_AGEMA_signal_1257, SubCellInst_SboxInst_15_XX_1_,
         new_AGEMA_signal_1259, SubCellInst_SboxInst_15_XX_2_,
         new_AGEMA_signal_1543, SubCellInst_SboxInst_15_Q0,
         new_AGEMA_signal_1544, SubCellInst_SboxInst_15_Q1,
         new_AGEMA_signal_1545, SubCellInst_SboxInst_15_Q4,
         new_AGEMA_signal_1546, SubCellInst_SboxInst_15_Q6,
         new_AGEMA_signal_1595, SubCellInst_SboxInst_15_L1,
         new_AGEMA_signal_1547, SubCellInst_SboxInst_15_L2,
         new_AGEMA_signal_1262, new_AGEMA_signal_1260, new_AGEMA_signal_1265,
         new_AGEMA_signal_1263, new_AGEMA_signal_1268, new_AGEMA_signal_1266,
         new_AGEMA_signal_1271, new_AGEMA_signal_1269, new_AGEMA_signal_1274,
         new_AGEMA_signal_1272, new_AGEMA_signal_1277, new_AGEMA_signal_1275,
         new_AGEMA_signal_1280, new_AGEMA_signal_1278, new_AGEMA_signal_1283,
         new_AGEMA_signal_1281, new_AGEMA_signal_1286, new_AGEMA_signal_1284,
         new_AGEMA_signal_1289, new_AGEMA_signal_1287, new_AGEMA_signal_1292,
         new_AGEMA_signal_1290, new_AGEMA_signal_1295, new_AGEMA_signal_1293,
         new_AGEMA_signal_1298, new_AGEMA_signal_1296, new_AGEMA_signal_1301,
         new_AGEMA_signal_1299, new_AGEMA_signal_1304, new_AGEMA_signal_1302,
         new_AGEMA_signal_1307, new_AGEMA_signal_1305, new_AGEMA_signal_1310,
         new_AGEMA_signal_1308, new_AGEMA_signal_1313, new_AGEMA_signal_1311,
         new_AGEMA_signal_1316, new_AGEMA_signal_1314, new_AGEMA_signal_1319,
         new_AGEMA_signal_1317, new_AGEMA_signal_1322, new_AGEMA_signal_1320,
         new_AGEMA_signal_1325, new_AGEMA_signal_1323, new_AGEMA_signal_1328,
         new_AGEMA_signal_1326, new_AGEMA_signal_1331, new_AGEMA_signal_1329,
         new_AGEMA_signal_1334, new_AGEMA_signal_1332, new_AGEMA_signal_1337,
         new_AGEMA_signal_1335, new_AGEMA_signal_1340, new_AGEMA_signal_1338,
         new_AGEMA_signal_1343, new_AGEMA_signal_1341, new_AGEMA_signal_1346,
         new_AGEMA_signal_1344, new_AGEMA_signal_1349, new_AGEMA_signal_1347,
         new_AGEMA_signal_1352, new_AGEMA_signal_1350, new_AGEMA_signal_1355,
         new_AGEMA_signal_1353, new_AGEMA_signal_1358, new_AGEMA_signal_1356,
         new_AGEMA_signal_1361, new_AGEMA_signal_1359, new_AGEMA_signal_1364,
         new_AGEMA_signal_1362, new_AGEMA_signal_1367, new_AGEMA_signal_1365,
         new_AGEMA_signal_1370, new_AGEMA_signal_1368, new_AGEMA_signal_1373,
         new_AGEMA_signal_1371, new_AGEMA_signal_1376, new_AGEMA_signal_1374,
         new_AGEMA_signal_1379, new_AGEMA_signal_1377, new_AGEMA_signal_1382,
         new_AGEMA_signal_1380, new_AGEMA_signal_1385, new_AGEMA_signal_1383,
         new_AGEMA_signal_1388, new_AGEMA_signal_1386, new_AGEMA_signal_1391,
         new_AGEMA_signal_1389, new_AGEMA_signal_1394, new_AGEMA_signal_1392,
         new_AGEMA_signal_1397, new_AGEMA_signal_1395, new_AGEMA_signal_1400,
         new_AGEMA_signal_1398, new_AGEMA_signal_1403, new_AGEMA_signal_1401,
         new_AGEMA_signal_1406, new_AGEMA_signal_1404, new_AGEMA_signal_1409,
         new_AGEMA_signal_1407, new_AGEMA_signal_1412, new_AGEMA_signal_1410,
         new_AGEMA_signal_1415, new_AGEMA_signal_1413, new_AGEMA_signal_1418,
         new_AGEMA_signal_1416, new_AGEMA_signal_1421, new_AGEMA_signal_1419,
         new_AGEMA_signal_1424, new_AGEMA_signal_1422, new_AGEMA_signal_1427,
         new_AGEMA_signal_1425, new_AGEMA_signal_1430, new_AGEMA_signal_1428,
         new_AGEMA_signal_1433, new_AGEMA_signal_1431, new_AGEMA_signal_1436,
         new_AGEMA_signal_1434, new_AGEMA_signal_1439, new_AGEMA_signal_1437,
         new_AGEMA_signal_1442, new_AGEMA_signal_1440, new_AGEMA_signal_1445,
         new_AGEMA_signal_1443, new_AGEMA_signal_1448, new_AGEMA_signal_1446,
         new_AGEMA_signal_1451, new_AGEMA_signal_1449, FSM_1,
         new_AGEMA_signal_2189, new_AGEMA_signal_2191, new_AGEMA_signal_2193,
         new_AGEMA_signal_2195, new_AGEMA_signal_2197, new_AGEMA_signal_2199,
         new_AGEMA_signal_2201, new_AGEMA_signal_2203, new_AGEMA_signal_2205,
         new_AGEMA_signal_2207, new_AGEMA_signal_2209, new_AGEMA_signal_2211,
         new_AGEMA_signal_2213, new_AGEMA_signal_2215, new_AGEMA_signal_2217,
         new_AGEMA_signal_2219, new_AGEMA_signal_2221, new_AGEMA_signal_2223,
         new_AGEMA_signal_2225, new_AGEMA_signal_2227, new_AGEMA_signal_2229,
         new_AGEMA_signal_2231, new_AGEMA_signal_2233, new_AGEMA_signal_2235,
         new_AGEMA_signal_2237, new_AGEMA_signal_2239, new_AGEMA_signal_2241,
         new_AGEMA_signal_2243, new_AGEMA_signal_2245, new_AGEMA_signal_2247,
         new_AGEMA_signal_2249, new_AGEMA_signal_2251, new_AGEMA_signal_2253,
         new_AGEMA_signal_2255, new_AGEMA_signal_2257, new_AGEMA_signal_2259,
         new_AGEMA_signal_2261, new_AGEMA_signal_2263, new_AGEMA_signal_2265,
         new_AGEMA_signal_2267, new_AGEMA_signal_2269, new_AGEMA_signal_2271,
         new_AGEMA_signal_2273, new_AGEMA_signal_2275, new_AGEMA_signal_2277,
         new_AGEMA_signal_2279, new_AGEMA_signal_2281, new_AGEMA_signal_2283,
         new_AGEMA_signal_2285, new_AGEMA_signal_2287, new_AGEMA_signal_2289,
         new_AGEMA_signal_2291, new_AGEMA_signal_2293, new_AGEMA_signal_2295,
         new_AGEMA_signal_2297, new_AGEMA_signal_2299, new_AGEMA_signal_2301,
         new_AGEMA_signal_2303, new_AGEMA_signal_2305, new_AGEMA_signal_2307,
         new_AGEMA_signal_2309, new_AGEMA_signal_2311, new_AGEMA_signal_2313,
         new_AGEMA_signal_2315, new_AGEMA_signal_2317, new_AGEMA_signal_2319,
         new_AGEMA_signal_2321, new_AGEMA_signal_2323, new_AGEMA_signal_2325,
         new_AGEMA_signal_2327, new_AGEMA_signal_2329, new_AGEMA_signal_2331,
         new_AGEMA_signal_2333, new_AGEMA_signal_2335, new_AGEMA_signal_2337,
         new_AGEMA_signal_2339, new_AGEMA_signal_2341, new_AGEMA_signal_2343,
         new_AGEMA_signal_2345, new_AGEMA_signal_2347, new_AGEMA_signal_2349,
         new_AGEMA_signal_2351, new_AGEMA_signal_2353, new_AGEMA_signal_2355,
         new_AGEMA_signal_2357, new_AGEMA_signal_2359, new_AGEMA_signal_2361,
         new_AGEMA_signal_2363, new_AGEMA_signal_2365, new_AGEMA_signal_2367,
         new_AGEMA_signal_2369, new_AGEMA_signal_2371, new_AGEMA_signal_2373,
         new_AGEMA_signal_2375, new_AGEMA_signal_2377, new_AGEMA_signal_2379,
         new_AGEMA_signal_2381, new_AGEMA_signal_2383, new_AGEMA_signal_2385,
         new_AGEMA_signal_2387, new_AGEMA_signal_2389, new_AGEMA_signal_2391,
         new_AGEMA_signal_2393, new_AGEMA_signal_2395, new_AGEMA_signal_2397,
         new_AGEMA_signal_2399, new_AGEMA_signal_2401, new_AGEMA_signal_2403,
         new_AGEMA_signal_2405, new_AGEMA_signal_2407, new_AGEMA_signal_2409,
         new_AGEMA_signal_2411, new_AGEMA_signal_2413, new_AGEMA_signal_2415,
         new_AGEMA_signal_2417, new_AGEMA_signal_2419, new_AGEMA_signal_2421,
         new_AGEMA_signal_2423, new_AGEMA_signal_2425, new_AGEMA_signal_2427,
         new_AGEMA_signal_2429, new_AGEMA_signal_2431, new_AGEMA_signal_2433,
         new_AGEMA_signal_2435, new_AGEMA_signal_2437, new_AGEMA_signal_2439,
         new_AGEMA_signal_2441, new_AGEMA_signal_2443, new_AGEMA_signal_2445,
         new_AGEMA_signal_2447, new_AGEMA_signal_2449, new_AGEMA_signal_2451,
         new_AGEMA_signal_2453, new_AGEMA_signal_2455, new_AGEMA_signal_2457,
         new_AGEMA_signal_2459, new_AGEMA_signal_2461, new_AGEMA_signal_2463,
         new_AGEMA_signal_2465, new_AGEMA_signal_2467, new_AGEMA_signal_2469,
         new_AGEMA_signal_2471, new_AGEMA_signal_2473, new_AGEMA_signal_2475,
         new_AGEMA_signal_2477, new_AGEMA_signal_2479, new_AGEMA_signal_2481,
         new_AGEMA_signal_2483, new_AGEMA_signal_2485, new_AGEMA_signal_2487,
         new_AGEMA_signal_2489, new_AGEMA_signal_2491, new_AGEMA_signal_2493,
         new_AGEMA_signal_2495, new_AGEMA_signal_2497, new_AGEMA_signal_2499,
         new_AGEMA_signal_2501, new_AGEMA_signal_2503, new_AGEMA_signal_2505,
         new_AGEMA_signal_2507, new_AGEMA_signal_2509, new_AGEMA_signal_2511,
         new_AGEMA_signal_2513, new_AGEMA_signal_2515, new_AGEMA_signal_2517,
         new_AGEMA_signal_2519, new_AGEMA_signal_2521, new_AGEMA_signal_2523,
         new_AGEMA_signal_2525, new_AGEMA_signal_2527, new_AGEMA_signal_2529,
         new_AGEMA_signal_2531, new_AGEMA_signal_2533, new_AGEMA_signal_2535,
         new_AGEMA_signal_2537, new_AGEMA_signal_2539, new_AGEMA_signal_2541,
         new_AGEMA_signal_2543, new_AGEMA_signal_2545, new_AGEMA_signal_2547,
         new_AGEMA_signal_2549, new_AGEMA_signal_2551, new_AGEMA_signal_2553,
         new_AGEMA_signal_2555, new_AGEMA_signal_2557, new_AGEMA_signal_2559,
         new_AGEMA_signal_2561, new_AGEMA_signal_2563, new_AGEMA_signal_2565,
         new_AGEMA_signal_2567, new_AGEMA_signal_2569, new_AGEMA_signal_2571,
         new_AGEMA_signal_2573, new_AGEMA_signal_2575, new_AGEMA_signal_2577,
         new_AGEMA_signal_2579, new_AGEMA_signal_2581, new_AGEMA_signal_2583,
         new_AGEMA_signal_2585, new_AGEMA_signal_2587, new_AGEMA_signal_2589,
         new_AGEMA_signal_2591, new_AGEMA_signal_2593, new_AGEMA_signal_2595,
         new_AGEMA_signal_2597, new_AGEMA_signal_2599, new_AGEMA_signal_2601,
         new_AGEMA_signal_2603, new_AGEMA_signal_2605, new_AGEMA_signal_2607,
         new_AGEMA_signal_2609, new_AGEMA_signal_2611, new_AGEMA_signal_2613,
         new_AGEMA_signal_2615, new_AGEMA_signal_2617, new_AGEMA_signal_2619,
         new_AGEMA_signal_2621, new_AGEMA_signal_2623, new_AGEMA_signal_2625,
         new_AGEMA_signal_2627, new_AGEMA_signal_2629, new_AGEMA_signal_2631,
         new_AGEMA_signal_2633, new_AGEMA_signal_2635, new_AGEMA_signal_2637,
         new_AGEMA_signal_2639, new_AGEMA_signal_2641, new_AGEMA_signal_2645,
         new_AGEMA_signal_2649, new_AGEMA_signal_2653, new_AGEMA_signal_2657,
         new_AGEMA_signal_2661, new_AGEMA_signal_2665, new_AGEMA_signal_2669,
         new_AGEMA_signal_2673, new_AGEMA_signal_2677, new_AGEMA_signal_2681,
         new_AGEMA_signal_2685, new_AGEMA_signal_2689, new_AGEMA_signal_2693,
         new_AGEMA_signal_2697, new_AGEMA_signal_2701, new_AGEMA_signal_2705,
         new_AGEMA_signal_2709, new_AGEMA_signal_2713, new_AGEMA_signal_2717,
         new_AGEMA_signal_2721, new_AGEMA_signal_2725, new_AGEMA_signal_2729,
         new_AGEMA_signal_2733, new_AGEMA_signal_2737, new_AGEMA_signal_2741,
         new_AGEMA_signal_2745, new_AGEMA_signal_2749, new_AGEMA_signal_2753,
         new_AGEMA_signal_2757, new_AGEMA_signal_2761, new_AGEMA_signal_2765,
         new_AGEMA_signal_2769, new_AGEMA_signal_2773, new_AGEMA_signal_2777,
         new_AGEMA_signal_2781, new_AGEMA_signal_2785, new_AGEMA_signal_2789,
         new_AGEMA_signal_2793, new_AGEMA_signal_2797, new_AGEMA_signal_2801,
         new_AGEMA_signal_2805, new_AGEMA_signal_2809, new_AGEMA_signal_2813,
         new_AGEMA_signal_2817, new_AGEMA_signal_2821, new_AGEMA_signal_2825,
         new_AGEMA_signal_2829, new_AGEMA_signal_2833, new_AGEMA_signal_2837,
         new_AGEMA_signal_2841, new_AGEMA_signal_2845, new_AGEMA_signal_2849,
         new_AGEMA_signal_2853, new_AGEMA_signal_2857, new_AGEMA_signal_2861,
         new_AGEMA_signal_2865, new_AGEMA_signal_2869, new_AGEMA_signal_2873,
         new_AGEMA_signal_2877, new_AGEMA_signal_2881, new_AGEMA_signal_2885,
         new_AGEMA_signal_2889, new_AGEMA_signal_2893, new_AGEMA_signal_2897,
         new_AGEMA_signal_2901, new_AGEMA_signal_2903, new_AGEMA_signal_2909,
         new_AGEMA_signal_2911, new_AGEMA_signal_2913, new_AGEMA_signal_2917,
         new_AGEMA_signal_2925, new_AGEMA_signal_2927, new_AGEMA_signal_2933,
         new_AGEMA_signal_2935, new_AGEMA_signal_2937, new_AGEMA_signal_2941,
         new_AGEMA_signal_2949, new_AGEMA_signal_2951, new_AGEMA_signal_2957,
         new_AGEMA_signal_2959, new_AGEMA_signal_2961, new_AGEMA_signal_2965,
         new_AGEMA_signal_2973, new_AGEMA_signal_2975, new_AGEMA_signal_2981,
         new_AGEMA_signal_2983, new_AGEMA_signal_2985, new_AGEMA_signal_2989,
         new_AGEMA_signal_2997, new_AGEMA_signal_2999, new_AGEMA_signal_3005,
         new_AGEMA_signal_3007, new_AGEMA_signal_3009, new_AGEMA_signal_3013,
         new_AGEMA_signal_3021, new_AGEMA_signal_3023, new_AGEMA_signal_3029,
         new_AGEMA_signal_3031, new_AGEMA_signal_3033, new_AGEMA_signal_3037,
         new_AGEMA_signal_3045, new_AGEMA_signal_3047, new_AGEMA_signal_3053,
         new_AGEMA_signal_3055, new_AGEMA_signal_3057, new_AGEMA_signal_3061,
         new_AGEMA_signal_3069, new_AGEMA_signal_3071, new_AGEMA_signal_3077,
         new_AGEMA_signal_3079, new_AGEMA_signal_3081, new_AGEMA_signal_3085,
         new_AGEMA_signal_3093, new_AGEMA_signal_3095, new_AGEMA_signal_3101,
         new_AGEMA_signal_3103, new_AGEMA_signal_3105, new_AGEMA_signal_3109,
         new_AGEMA_signal_3117, new_AGEMA_signal_3119, new_AGEMA_signal_3125,
         new_AGEMA_signal_3127, new_AGEMA_signal_3129, new_AGEMA_signal_3133,
         new_AGEMA_signal_3141, new_AGEMA_signal_3143, new_AGEMA_signal_3149,
         new_AGEMA_signal_3151, new_AGEMA_signal_3153, new_AGEMA_signal_3157,
         new_AGEMA_signal_3165, new_AGEMA_signal_3167, new_AGEMA_signal_3173,
         new_AGEMA_signal_3175, new_AGEMA_signal_3177, new_AGEMA_signal_3181,
         new_AGEMA_signal_3189, new_AGEMA_signal_3191, new_AGEMA_signal_3197,
         new_AGEMA_signal_3199, new_AGEMA_signal_3201, new_AGEMA_signal_3205,
         new_AGEMA_signal_3213, new_AGEMA_signal_3215, new_AGEMA_signal_3221,
         new_AGEMA_signal_3223, new_AGEMA_signal_3225, new_AGEMA_signal_3229,
         new_AGEMA_signal_3237, new_AGEMA_signal_3239, new_AGEMA_signal_3245,
         new_AGEMA_signal_3247, new_AGEMA_signal_3249, new_AGEMA_signal_3253,
         new_AGEMA_signal_3261, new_AGEMA_signal_3263, new_AGEMA_signal_3269,
         new_AGEMA_signal_3271, new_AGEMA_signal_3273, new_AGEMA_signal_3277,
         new_AGEMA_signal_3285, new_AGEMA_signal_3289, new_AGEMA_signal_3293,
         new_AGEMA_signal_3297, new_AGEMA_signal_3301, new_AGEMA_signal_3305,
         new_AGEMA_signal_3309, new_AGEMA_signal_3313, new_AGEMA_signal_3317,
         new_AGEMA_signal_3321, new_AGEMA_signal_3325, new_AGEMA_signal_3329,
         new_AGEMA_signal_3333, new_AGEMA_signal_3337, new_AGEMA_signal_3341,
         new_AGEMA_signal_3345, new_AGEMA_signal_3349, new_AGEMA_signal_3353,
         new_AGEMA_signal_3357, new_AGEMA_signal_3361, new_AGEMA_signal_3365,
         new_AGEMA_signal_3369, new_AGEMA_signal_3373, new_AGEMA_signal_3377,
         new_AGEMA_signal_3381, new_AGEMA_signal_3385, new_AGEMA_signal_3389,
         new_AGEMA_signal_3393, new_AGEMA_signal_3397, new_AGEMA_signal_3401,
         new_AGEMA_signal_3405, new_AGEMA_signal_3409, new_AGEMA_signal_3413,
         new_AGEMA_signal_3417, new_AGEMA_signal_3421, new_AGEMA_signal_3425,
         new_AGEMA_signal_3557, new_AGEMA_signal_3561, new_AGEMA_signal_3565,
         new_AGEMA_signal_3569, new_AGEMA_signal_3573, new_AGEMA_signal_3577,
         new_AGEMA_signal_3581, new_AGEMA_signal_3585, new_AGEMA_signal_3589,
         new_AGEMA_signal_3593, new_AGEMA_signal_3597, new_AGEMA_signal_3601,
         new_AGEMA_signal_3605, new_AGEMA_signal_3609, new_AGEMA_signal_3613,
         new_AGEMA_signal_3617, new_AGEMA_signal_3621, new_AGEMA_signal_3625,
         new_AGEMA_signal_3629, new_AGEMA_signal_3633, new_AGEMA_signal_3637,
         new_AGEMA_signal_3641, new_AGEMA_signal_3645, new_AGEMA_signal_3649,
         new_AGEMA_signal_3653, new_AGEMA_signal_3657, new_AGEMA_signal_3661,
         new_AGEMA_signal_3665, new_AGEMA_signal_3669, new_AGEMA_signal_3673,
         new_AGEMA_signal_3677, new_AGEMA_signal_3681, new_AGEMA_signal_3685,
         new_AGEMA_signal_3689, new_AGEMA_signal_3693, new_AGEMA_signal_3697,
         new_AGEMA_signal_3701, new_AGEMA_signal_3705, new_AGEMA_signal_3709,
         new_AGEMA_signal_3713, new_AGEMA_signal_3717, new_AGEMA_signal_3721,
         new_AGEMA_signal_3725, new_AGEMA_signal_3729, new_AGEMA_signal_3733,
         new_AGEMA_signal_3737, new_AGEMA_signal_3741, new_AGEMA_signal_3745,
         new_AGEMA_signal_3749, new_AGEMA_signal_3753, new_AGEMA_signal_3757,
         new_AGEMA_signal_3761, new_AGEMA_signal_3765, new_AGEMA_signal_3769,
         new_AGEMA_signal_3773, new_AGEMA_signal_3777, new_AGEMA_signal_3781,
         new_AGEMA_signal_3785, new_AGEMA_signal_3789, new_AGEMA_signal_3793,
         new_AGEMA_signal_3797, new_AGEMA_signal_3801, new_AGEMA_signal_3805,
         new_AGEMA_signal_3809, new_AGEMA_signal_3813, new_AGEMA_signal_3817,
         new_AGEMA_signal_3821, new_AGEMA_signal_3825, new_AGEMA_signal_3829,
         new_AGEMA_signal_3833, new_AGEMA_signal_3837, new_AGEMA_signal_3841,
         new_AGEMA_signal_3845, new_AGEMA_signal_3849, new_AGEMA_signal_3853,
         new_AGEMA_signal_3857, new_AGEMA_signal_3861, new_AGEMA_signal_3865,
         new_AGEMA_signal_3869, new_AGEMA_signal_3873, new_AGEMA_signal_3877,
         new_AGEMA_signal_3881, new_AGEMA_signal_3885, new_AGEMA_signal_3889,
         new_AGEMA_signal_3893, new_AGEMA_signal_3897, new_AGEMA_signal_3901,
         new_AGEMA_signal_3905, new_AGEMA_signal_3909, new_AGEMA_signal_3913,
         new_AGEMA_signal_3917, new_AGEMA_signal_3921, new_AGEMA_signal_3925,
         new_AGEMA_signal_3929, new_AGEMA_signal_3933, new_AGEMA_signal_3937,
         new_AGEMA_signal_3941, new_AGEMA_signal_3945, new_AGEMA_signal_3949,
         new_AGEMA_signal_3953, new_AGEMA_signal_3957, new_AGEMA_signal_3961,
         new_AGEMA_signal_3965, new_AGEMA_signal_3969, new_AGEMA_signal_3973,
         new_AGEMA_signal_3977, new_AGEMA_signal_3981, new_AGEMA_signal_3985,
         new_AGEMA_signal_3989, new_AGEMA_signal_3993, new_AGEMA_signal_3997,
         new_AGEMA_signal_4001, new_AGEMA_signal_4005, new_AGEMA_signal_4009,
         new_AGEMA_signal_4013, new_AGEMA_signal_4017, new_AGEMA_signal_4021,
         new_AGEMA_signal_4025, new_AGEMA_signal_4029, new_AGEMA_signal_4033,
         new_AGEMA_signal_4037, new_AGEMA_signal_4041, new_AGEMA_signal_4045,
         new_AGEMA_signal_4049, new_AGEMA_signal_4053, new_AGEMA_signal_4057,
         new_AGEMA_signal_4061, new_AGEMA_signal_4065, new_AGEMA_signal_4069,
         new_AGEMA_signal_4073, new_AGEMA_signal_4077, new_AGEMA_signal_4081,
         new_AGEMA_signal_4085, new_AGEMA_signal_4089, new_AGEMA_signal_2190,
         new_AGEMA_signal_1922, new_AGEMA_signal_2194, new_AGEMA_signal_2192,
         new_AGEMA_signal_1915, new_AGEMA_signal_1982, new_AGEMA_signal_2198,
         new_AGEMA_signal_2196, new_AGEMA_signal_1975, new_AGEMA_signal_1924,
         new_AGEMA_signal_2202, new_AGEMA_signal_2200, new_AGEMA_signal_1917,
         new_AGEMA_signal_1984, new_AGEMA_signal_2206, new_AGEMA_signal_2204,
         new_AGEMA_signal_1977, new_AGEMA_signal_1926, new_AGEMA_signal_2210,
         new_AGEMA_signal_2208, new_AGEMA_signal_1919, new_AGEMA_signal_1986,
         new_AGEMA_signal_2214, new_AGEMA_signal_2212, new_AGEMA_signal_1979,
         new_AGEMA_signal_2042, new_AGEMA_signal_2218, new_AGEMA_signal_2216,
         new_AGEMA_signal_2033, new_AGEMA_signal_2085, new_AGEMA_signal_2222,
         new_AGEMA_signal_2220, new_AGEMA_signal_2077, new_AGEMA_signal_1928,
         new_AGEMA_signal_2226, new_AGEMA_signal_2224, new_AGEMA_signal_1909,
         new_AGEMA_signal_1988, new_AGEMA_signal_2230, new_AGEMA_signal_2228,
         new_AGEMA_signal_1968, new_AGEMA_signal_1930, new_AGEMA_signal_2234,
         new_AGEMA_signal_2232, new_AGEMA_signal_1911, new_AGEMA_signal_1990,
         new_AGEMA_signal_2238, new_AGEMA_signal_2236, new_AGEMA_signal_1970,
         new_AGEMA_signal_2048, new_AGEMA_signal_2242, new_AGEMA_signal_2240,
         new_AGEMA_signal_2023, new_AGEMA_signal_2091, new_AGEMA_signal_2246,
         new_AGEMA_signal_2244, new_AGEMA_signal_2071, new_AGEMA_signal_1932,
         new_AGEMA_signal_2250, new_AGEMA_signal_2248, new_AGEMA_signal_1913,
         new_AGEMA_signal_1992, new_AGEMA_signal_2254, new_AGEMA_signal_2252,
         new_AGEMA_signal_1973, new_AGEMA_signal_1821, new_AGEMA_signal_2258,
         new_AGEMA_signal_2256, new_AGEMA_signal_1810, new_AGEMA_signal_1874,
         new_AGEMA_signal_2262, new_AGEMA_signal_2260, new_AGEMA_signal_1854,
         new_AGEMA_signal_1823, new_AGEMA_signal_2266, new_AGEMA_signal_2264,
         new_AGEMA_signal_1812, new_AGEMA_signal_1876, new_AGEMA_signal_2270,
         new_AGEMA_signal_2268, new_AGEMA_signal_1856, new_AGEMA_signal_1825,
         new_AGEMA_signal_2274, new_AGEMA_signal_2272, new_AGEMA_signal_1814,
         new_AGEMA_signal_1878, new_AGEMA_signal_2278, new_AGEMA_signal_2276,
         new_AGEMA_signal_1858, new_AGEMA_signal_1940, new_AGEMA_signal_2282,
         new_AGEMA_signal_2280, new_AGEMA_signal_1898, new_AGEMA_signal_2000,
         new_AGEMA_signal_2286, new_AGEMA_signal_2284, new_AGEMA_signal_1958,
         new_AGEMA_signal_1942, new_AGEMA_signal_2290, new_AGEMA_signal_2288,
         new_AGEMA_signal_1901, new_AGEMA_signal_2002, new_AGEMA_signal_2294,
         new_AGEMA_signal_2292, new_AGEMA_signal_1960, new_AGEMA_signal_1944,
         new_AGEMA_signal_2298, new_AGEMA_signal_2296, new_AGEMA_signal_1903,
         new_AGEMA_signal_2004, new_AGEMA_signal_2302, new_AGEMA_signal_2300,
         new_AGEMA_signal_1963, new_AGEMA_signal_1946, new_AGEMA_signal_2306,
         new_AGEMA_signal_2304, new_AGEMA_signal_1906, new_AGEMA_signal_2006,
         new_AGEMA_signal_2310, new_AGEMA_signal_2308, new_AGEMA_signal_1965,
         new_AGEMA_signal_2060, new_AGEMA_signal_2314, new_AGEMA_signal_2312,
         new_AGEMA_signal_2017, new_AGEMA_signal_2103, new_AGEMA_signal_2318,
         new_AGEMA_signal_2316, new_AGEMA_signal_2067, new_AGEMA_signal_1724,
         SubCellInst_SboxInst_0_YY_1_, new_AGEMA_signal_1660,
         SubCellInst_SboxInst_0_YY_0_, new_AGEMA_signal_1548,
         SubCellInst_SboxInst_0_T0, new_AGEMA_signal_1596,
         SubCellInst_SboxInst_0_Q2, new_AGEMA_signal_2322,
         new_AGEMA_signal_2320, new_AGEMA_signal_1549,
         SubCellInst_SboxInst_0_T2, new_AGEMA_signal_1597,
         SubCellInst_SboxInst_0_Q7, new_AGEMA_signal_2326,
         new_AGEMA_signal_2324, new_AGEMA_signal_1598,
         SubCellInst_SboxInst_0_L3, new_AGEMA_signal_2330,
         new_AGEMA_signal_2328, new_AGEMA_signal_2334, new_AGEMA_signal_2332,
         new_AGEMA_signal_1726, SubCellInst_SboxInst_1_YY_1_,
         new_AGEMA_signal_1664, SubCellInst_SboxInst_1_YY_0_,
         new_AGEMA_signal_1551, SubCellInst_SboxInst_1_T0,
         new_AGEMA_signal_1600, SubCellInst_SboxInst_1_Q2,
         new_AGEMA_signal_2338, new_AGEMA_signal_2336, new_AGEMA_signal_1552,
         SubCellInst_SboxInst_1_T2, new_AGEMA_signal_1601,
         SubCellInst_SboxInst_1_Q7, new_AGEMA_signal_2342,
         new_AGEMA_signal_2340, new_AGEMA_signal_1602,
         SubCellInst_SboxInst_1_L3, new_AGEMA_signal_2346,
         new_AGEMA_signal_2344, new_AGEMA_signal_2350, new_AGEMA_signal_2348,
         new_AGEMA_signal_1728, SubCellInst_SboxInst_2_YY_1_,
         new_AGEMA_signal_1668, SubCellInst_SboxInst_2_YY_0_,
         new_AGEMA_signal_1554, SubCellInst_SboxInst_2_T0,
         new_AGEMA_signal_1604, SubCellInst_SboxInst_2_Q2,
         new_AGEMA_signal_2354, new_AGEMA_signal_2352, new_AGEMA_signal_1555,
         SubCellInst_SboxInst_2_T2, new_AGEMA_signal_1605,
         SubCellInst_SboxInst_2_Q7, new_AGEMA_signal_2358,
         new_AGEMA_signal_2356, new_AGEMA_signal_1606,
         SubCellInst_SboxInst_2_L3, new_AGEMA_signal_2362,
         new_AGEMA_signal_2360, new_AGEMA_signal_2366, new_AGEMA_signal_2364,
         new_AGEMA_signal_1730, SubCellInst_SboxInst_3_YY_1_,
         new_AGEMA_signal_1672, SubCellInst_SboxInst_3_YY_0_,
         new_AGEMA_signal_1557, SubCellInst_SboxInst_3_T0,
         new_AGEMA_signal_1608, SubCellInst_SboxInst_3_Q2,
         new_AGEMA_signal_2370, new_AGEMA_signal_2368, new_AGEMA_signal_1558,
         SubCellInst_SboxInst_3_T2, new_AGEMA_signal_1609,
         SubCellInst_SboxInst_3_Q7, new_AGEMA_signal_2374,
         new_AGEMA_signal_2372, new_AGEMA_signal_1610,
         SubCellInst_SboxInst_3_L3, new_AGEMA_signal_2378,
         new_AGEMA_signal_2376, new_AGEMA_signal_2382, new_AGEMA_signal_2380,
         new_AGEMA_signal_1732, SubCellInst_SboxInst_4_YY_1_,
         new_AGEMA_signal_1676, SubCellInst_SboxInst_4_YY_0_,
         new_AGEMA_signal_1560, SubCellInst_SboxInst_4_T0,
         new_AGEMA_signal_1612, SubCellInst_SboxInst_4_Q2,
         new_AGEMA_signal_2386, new_AGEMA_signal_2384, new_AGEMA_signal_1561,
         SubCellInst_SboxInst_4_T2, new_AGEMA_signal_1613,
         SubCellInst_SboxInst_4_Q7, new_AGEMA_signal_2390,
         new_AGEMA_signal_2388, new_AGEMA_signal_1614,
         SubCellInst_SboxInst_4_L3, new_AGEMA_signal_2394,
         new_AGEMA_signal_2392, new_AGEMA_signal_2398, new_AGEMA_signal_2396,
         new_AGEMA_signal_1734, SubCellInst_SboxInst_5_YY_1_,
         new_AGEMA_signal_1680, SubCellInst_SboxInst_5_YY_0_,
         new_AGEMA_signal_1563, SubCellInst_SboxInst_5_T0,
         new_AGEMA_signal_1616, SubCellInst_SboxInst_5_Q2,
         new_AGEMA_signal_2402, new_AGEMA_signal_2400, new_AGEMA_signal_1564,
         SubCellInst_SboxInst_5_T2, new_AGEMA_signal_1617,
         SubCellInst_SboxInst_5_Q7, new_AGEMA_signal_2406,
         new_AGEMA_signal_2404, new_AGEMA_signal_1618,
         SubCellInst_SboxInst_5_L3, new_AGEMA_signal_2410,
         new_AGEMA_signal_2408, new_AGEMA_signal_2414, new_AGEMA_signal_2412,
         new_AGEMA_signal_1736, SubCellInst_SboxInst_6_YY_1_,
         new_AGEMA_signal_1684, SubCellInst_SboxInst_6_YY_0_,
         new_AGEMA_signal_1566, SubCellInst_SboxInst_6_T0,
         new_AGEMA_signal_1620, SubCellInst_SboxInst_6_Q2,
         new_AGEMA_signal_2418, new_AGEMA_signal_2416, new_AGEMA_signal_1567,
         SubCellInst_SboxInst_6_T2, new_AGEMA_signal_1621,
         SubCellInst_SboxInst_6_Q7, new_AGEMA_signal_2422,
         new_AGEMA_signal_2420, new_AGEMA_signal_1622,
         SubCellInst_SboxInst_6_L3, new_AGEMA_signal_2426,
         new_AGEMA_signal_2424, new_AGEMA_signal_2430, new_AGEMA_signal_2428,
         new_AGEMA_signal_1738, SubCellInst_SboxInst_7_YY_1_,
         new_AGEMA_signal_1688, SubCellInst_SboxInst_7_YY_0_,
         new_AGEMA_signal_1569, SubCellInst_SboxInst_7_T0,
         new_AGEMA_signal_1624, SubCellInst_SboxInst_7_Q2,
         new_AGEMA_signal_2434, new_AGEMA_signal_2432, new_AGEMA_signal_1570,
         SubCellInst_SboxInst_7_T2, new_AGEMA_signal_1625,
         SubCellInst_SboxInst_7_Q7, new_AGEMA_signal_2438,
         new_AGEMA_signal_2436, new_AGEMA_signal_1626,
         SubCellInst_SboxInst_7_L3, new_AGEMA_signal_2442,
         new_AGEMA_signal_2440, new_AGEMA_signal_2446, new_AGEMA_signal_2444,
         new_AGEMA_signal_1740, SubCellInst_SboxInst_8_YY_1_,
         new_AGEMA_signal_1692, SubCellInst_SboxInst_8_YY_0_,
         new_AGEMA_signal_1572, SubCellInst_SboxInst_8_T0,
         new_AGEMA_signal_1628, SubCellInst_SboxInst_8_Q2,
         new_AGEMA_signal_2450, new_AGEMA_signal_2448, new_AGEMA_signal_1573,
         SubCellInst_SboxInst_8_T2, new_AGEMA_signal_1629,
         SubCellInst_SboxInst_8_Q7, new_AGEMA_signal_2454,
         new_AGEMA_signal_2452, new_AGEMA_signal_1630,
         SubCellInst_SboxInst_8_L3, new_AGEMA_signal_2458,
         new_AGEMA_signal_2456, new_AGEMA_signal_2462, new_AGEMA_signal_2460,
         new_AGEMA_signal_1742, SubCellInst_SboxInst_9_YY_1_,
         new_AGEMA_signal_1696, SubCellInst_SboxInst_9_YY_0_,
         new_AGEMA_signal_1575, SubCellInst_SboxInst_9_T0,
         new_AGEMA_signal_1632, SubCellInst_SboxInst_9_Q2,
         new_AGEMA_signal_2466, new_AGEMA_signal_2464, new_AGEMA_signal_1576,
         SubCellInst_SboxInst_9_T2, new_AGEMA_signal_1633,
         SubCellInst_SboxInst_9_Q7, new_AGEMA_signal_2470,
         new_AGEMA_signal_2468, new_AGEMA_signal_1634,
         SubCellInst_SboxInst_9_L3, new_AGEMA_signal_2474,
         new_AGEMA_signal_2472, new_AGEMA_signal_2478, new_AGEMA_signal_2476,
         new_AGEMA_signal_1744, SubCellInst_SboxInst_10_YY_1_,
         new_AGEMA_signal_1700, SubCellInst_SboxInst_10_YY_0_,
         new_AGEMA_signal_1578, SubCellInst_SboxInst_10_T0,
         new_AGEMA_signal_1636, SubCellInst_SboxInst_10_Q2,
         new_AGEMA_signal_2482, new_AGEMA_signal_2480, new_AGEMA_signal_1579,
         SubCellInst_SboxInst_10_T2, new_AGEMA_signal_1637,
         SubCellInst_SboxInst_10_Q7, new_AGEMA_signal_2486,
         new_AGEMA_signal_2484, new_AGEMA_signal_1638,
         SubCellInst_SboxInst_10_L3, new_AGEMA_signal_2490,
         new_AGEMA_signal_2488, new_AGEMA_signal_2494, new_AGEMA_signal_2492,
         SubCellOutput_47, SubCellOutput_46, SubCellOutput_45,
         SubCellOutput_44, SubCellOutput_29, new_AGEMA_signal_1746,
         SubCellInst_SboxInst_11_YY_1_, new_AGEMA_signal_1704,
         SubCellInst_SboxInst_11_YY_0_, new_AGEMA_signal_1581,
         SubCellInst_SboxInst_11_T0, new_AGEMA_signal_1640,
         SubCellInst_SboxInst_11_Q2, new_AGEMA_signal_2498,
         new_AGEMA_signal_2496, new_AGEMA_signal_1582,
         SubCellInst_SboxInst_11_T2, new_AGEMA_signal_1641,
         SubCellInst_SboxInst_11_Q7, new_AGEMA_signal_2502,
         new_AGEMA_signal_2500, new_AGEMA_signal_1642,
         SubCellInst_SboxInst_11_L3, new_AGEMA_signal_2506,
         new_AGEMA_signal_2504, new_AGEMA_signal_2510, new_AGEMA_signal_2508,
         new_AGEMA_signal_1748, SubCellInst_SboxInst_12_YY_1_,
         new_AGEMA_signal_1708, SubCellInst_SboxInst_12_YY_0_,
         new_AGEMA_signal_1584, SubCellInst_SboxInst_12_T0,
         new_AGEMA_signal_1644, SubCellInst_SboxInst_12_Q2,
         new_AGEMA_signal_2514, new_AGEMA_signal_2512, new_AGEMA_signal_1585,
         SubCellInst_SboxInst_12_T2, new_AGEMA_signal_1645,
         SubCellInst_SboxInst_12_Q7, new_AGEMA_signal_2518,
         new_AGEMA_signal_2516, new_AGEMA_signal_1646,
         SubCellInst_SboxInst_12_L3, new_AGEMA_signal_2522,
         new_AGEMA_signal_2520, new_AGEMA_signal_2526, new_AGEMA_signal_2524,
         new_AGEMA_signal_1750, SubCellInst_SboxInst_13_YY_1_,
         new_AGEMA_signal_1712, SubCellInst_SboxInst_13_YY_0_,
         new_AGEMA_signal_1587, SubCellInst_SboxInst_13_T0,
         new_AGEMA_signal_1648, SubCellInst_SboxInst_13_Q2,
         new_AGEMA_signal_2530, new_AGEMA_signal_2528, new_AGEMA_signal_1588,
         SubCellInst_SboxInst_13_T2, new_AGEMA_signal_1649,
         SubCellInst_SboxInst_13_Q7, new_AGEMA_signal_2534,
         new_AGEMA_signal_2532, new_AGEMA_signal_1650,
         SubCellInst_SboxInst_13_L3, new_AGEMA_signal_2538,
         new_AGEMA_signal_2536, new_AGEMA_signal_2542, new_AGEMA_signal_2540,
         new_AGEMA_signal_1752, SubCellInst_SboxInst_14_YY_1_,
         new_AGEMA_signal_1716, SubCellInst_SboxInst_14_YY_0_,
         new_AGEMA_signal_1590, SubCellInst_SboxInst_14_T0,
         new_AGEMA_signal_1652, SubCellInst_SboxInst_14_Q2,
         new_AGEMA_signal_2546, new_AGEMA_signal_2544, new_AGEMA_signal_1591,
         SubCellInst_SboxInst_14_T2, new_AGEMA_signal_1653,
         SubCellInst_SboxInst_14_Q7, new_AGEMA_signal_2550,
         new_AGEMA_signal_2548, new_AGEMA_signal_1654,
         SubCellInst_SboxInst_14_L3, new_AGEMA_signal_2554,
         new_AGEMA_signal_2552, new_AGEMA_signal_2558, new_AGEMA_signal_2556,
         new_AGEMA_signal_1754, SubCellInst_SboxInst_15_YY_1_,
         new_AGEMA_signal_1720, SubCellInst_SboxInst_15_YY_0_,
         new_AGEMA_signal_1593, SubCellInst_SboxInst_15_T0,
         new_AGEMA_signal_1656, SubCellInst_SboxInst_15_Q2,
         new_AGEMA_signal_2562, new_AGEMA_signal_2560, new_AGEMA_signal_1594,
         SubCellInst_SboxInst_15_T2, new_AGEMA_signal_1657,
         SubCellInst_SboxInst_15_Q7, new_AGEMA_signal_2566,
         new_AGEMA_signal_2564, new_AGEMA_signal_1658,
         SubCellInst_SboxInst_15_L3, new_AGEMA_signal_2570,
         new_AGEMA_signal_2568, new_AGEMA_signal_2574, new_AGEMA_signal_2572,
         new_AGEMA_signal_1800, new_AGEMA_signal_2576, new_AGEMA_signal_1756,
         AddConstXOR_AddConstXOR_XORInst_0_2_n1, new_AGEMA_signal_1843,
         new_AGEMA_signal_2578, new_AGEMA_signal_1801,
         AddConstXOR_AddConstXOR_XORInst_0_3_n1, new_AGEMA_signal_1802,
         new_AGEMA_signal_1757, AddConstXOR_AddConstXOR_XORInst_1_2_n1,
         new_AGEMA_signal_1845, new_AGEMA_signal_1803,
         AddConstXOR_AddConstXOR_XORInst_1_3_n1, new_AGEMA_signal_1804,
         new_AGEMA_signal_2582, new_AGEMA_signal_2580, new_AGEMA_signal_1758,
         AddRoundTweakeyXOR_XORInst_0_2_n1, new_AGEMA_signal_1847,
         new_AGEMA_signal_2586, new_AGEMA_signal_2584, new_AGEMA_signal_1805,
         AddRoundTweakeyXOR_XORInst_0_3_n1, new_AGEMA_signal_1806,
         new_AGEMA_signal_2590, new_AGEMA_signal_2588, new_AGEMA_signal_1759,
         AddRoundTweakeyXOR_XORInst_1_2_n1, new_AGEMA_signal_1849,
         new_AGEMA_signal_2594, new_AGEMA_signal_2592, new_AGEMA_signal_1807,
         AddRoundTweakeyXOR_XORInst_1_3_n1, new_AGEMA_signal_1808,
         new_AGEMA_signal_2598, new_AGEMA_signal_2596, new_AGEMA_signal_1760,
         AddRoundTweakeyXOR_XORInst_2_2_n1, new_AGEMA_signal_1851,
         new_AGEMA_signal_2602, new_AGEMA_signal_2600, new_AGEMA_signal_1809,
         AddRoundTweakeyXOR_XORInst_2_3_n1, new_AGEMA_signal_1890,
         new_AGEMA_signal_2606, new_AGEMA_signal_2604, new_AGEMA_signal_1852,
         AddRoundTweakeyXOR_XORInst_3_2_n1, new_AGEMA_signal_1953,
         new_AGEMA_signal_2610, new_AGEMA_signal_2608, new_AGEMA_signal_1891,
         AddRoundTweakeyXOR_XORInst_3_3_n1, new_AGEMA_signal_2614,
         new_AGEMA_signal_2612, new_AGEMA_signal_1761,
         AddRoundTweakeyXOR_XORInst_4_2_n1, new_AGEMA_signal_2618,
         new_AGEMA_signal_2616, new_AGEMA_signal_1811,
         AddRoundTweakeyXOR_XORInst_4_3_n1, new_AGEMA_signal_2622,
         new_AGEMA_signal_2620, new_AGEMA_signal_1762,
         AddRoundTweakeyXOR_XORInst_5_2_n1, new_AGEMA_signal_2626,
         new_AGEMA_signal_2624, new_AGEMA_signal_1813,
         AddRoundTweakeyXOR_XORInst_5_3_n1, new_AGEMA_signal_2630,
         new_AGEMA_signal_2628, new_AGEMA_signal_1763,
         AddRoundTweakeyXOR_XORInst_6_2_n1, new_AGEMA_signal_2634,
         new_AGEMA_signal_2632, new_AGEMA_signal_1815,
         AddRoundTweakeyXOR_XORInst_6_3_n1, new_AGEMA_signal_2638,
         new_AGEMA_signal_2636, new_AGEMA_signal_1859,
         AddRoundTweakeyXOR_XORInst_7_2_n1, new_AGEMA_signal_2642,
         new_AGEMA_signal_2640, new_AGEMA_signal_1899,
         AddRoundTweakeyXOR_XORInst_7_3_n1, new_AGEMA_signal_1764,
         MCInst_MCR0_XORInst_0_2_n1, new_AGEMA_signal_1861,
         MCInst_MCR0_XORInst_0_2_n2, new_AGEMA_signal_1816,
         MCInst_MCR0_XORInst_0_3_n1, new_AGEMA_signal_1902,
         MCInst_MCR0_XORInst_0_3_n2, new_AGEMA_signal_1765,
         MCInst_MCR0_XORInst_1_2_n1, new_AGEMA_signal_1863,
         MCInst_MCR0_XORInst_1_2_n2, new_AGEMA_signal_1817,
         MCInst_MCR0_XORInst_1_3_n1, new_AGEMA_signal_1904,
         MCInst_MCR0_XORInst_1_3_n2, new_AGEMA_signal_1766,
         MCInst_MCR0_XORInst_2_2_n1, new_AGEMA_signal_1865,
         MCInst_MCR0_XORInst_2_2_n2, new_AGEMA_signal_1818,
         MCInst_MCR0_XORInst_2_3_n1, new_AGEMA_signal_1907,
         MCInst_MCR0_XORInst_2_3_n2, new_AGEMA_signal_1767,
         MCInst_MCR0_XORInst_3_2_n1, new_AGEMA_signal_1966,
         MCInst_MCR0_XORInst_3_2_n2, new_AGEMA_signal_1819,
         MCInst_MCR0_XORInst_3_3_n1, new_AGEMA_signal_2018,
         MCInst_MCR0_XORInst_3_3_n2, new_AGEMA_signal_1867,
         MCInst_MCR2_XORInst_0_2_n1, new_AGEMA_signal_1910,
         MCInst_MCR2_XORInst_0_3_n1, new_AGEMA_signal_1868,
         MCInst_MCR2_XORInst_1_2_n1, new_AGEMA_signal_1912,
         MCInst_MCR2_XORInst_1_3_n1, new_AGEMA_signal_1971,
         MCInst_MCR2_XORInst_2_2_n1, new_AGEMA_signal_2024,
         MCInst_MCR2_XORInst_2_3_n1, new_AGEMA_signal_1869,
         MCInst_MCR2_XORInst_3_2_n1, new_AGEMA_signal_1914,
         MCInst_MCR2_XORInst_3_3_n1, new_AGEMA_signal_1870,
         MCInst_MCR3_XORInst_0_2_n1, new_AGEMA_signal_1916,
         MCInst_MCR3_XORInst_0_3_n1, new_AGEMA_signal_1871,
         MCInst_MCR3_XORInst_1_2_n1, new_AGEMA_signal_1918,
         MCInst_MCR3_XORInst_1_3_n1, new_AGEMA_signal_1872,
         MCInst_MCR3_XORInst_2_2_n1, new_AGEMA_signal_1920,
         MCInst_MCR3_XORInst_2_3_n1, new_AGEMA_signal_1980,
         MCInst_MCR3_XORInst_3_2_n1, new_AGEMA_signal_2034,
         MCInst_MCR3_XORInst_3_3_n1, new_AGEMA_signal_2646,
         new_AGEMA_signal_2650, new_AGEMA_signal_2654, new_AGEMA_signal_2658,
         new_AGEMA_signal_2662, new_AGEMA_signal_2666, new_AGEMA_signal_2670,
         new_AGEMA_signal_2674, new_AGEMA_signal_2678, new_AGEMA_signal_2682,
         new_AGEMA_signal_2686, new_AGEMA_signal_2690, new_AGEMA_signal_2694,
         new_AGEMA_signal_2698, new_AGEMA_signal_2702, new_AGEMA_signal_2706,
         new_AGEMA_signal_2710, new_AGEMA_signal_2714, new_AGEMA_signal_2718,
         new_AGEMA_signal_2722, new_AGEMA_signal_2726, new_AGEMA_signal_2730,
         new_AGEMA_signal_2734, new_AGEMA_signal_2738, new_AGEMA_signal_2742,
         new_AGEMA_signal_2746, new_AGEMA_signal_2750, new_AGEMA_signal_2754,
         new_AGEMA_signal_2758, new_AGEMA_signal_2762, new_AGEMA_signal_2766,
         new_AGEMA_signal_2770, new_AGEMA_signal_2774, new_AGEMA_signal_2778,
         new_AGEMA_signal_2782, new_AGEMA_signal_2786, new_AGEMA_signal_2790,
         new_AGEMA_signal_2794, new_AGEMA_signal_2798, new_AGEMA_signal_2802,
         new_AGEMA_signal_2806, new_AGEMA_signal_2810, new_AGEMA_signal_2814,
         new_AGEMA_signal_2818, new_AGEMA_signal_2822, new_AGEMA_signal_2826,
         new_AGEMA_signal_2830, new_AGEMA_signal_2834, new_AGEMA_signal_2838,
         new_AGEMA_signal_2842, new_AGEMA_signal_2846, new_AGEMA_signal_2850,
         new_AGEMA_signal_2854, new_AGEMA_signal_2858, new_AGEMA_signal_2862,
         new_AGEMA_signal_2866, new_AGEMA_signal_2870, new_AGEMA_signal_2874,
         new_AGEMA_signal_2878, new_AGEMA_signal_2882, new_AGEMA_signal_2886,
         new_AGEMA_signal_2890, new_AGEMA_signal_2894, new_AGEMA_signal_2898,
         new_AGEMA_signal_2902, new_AGEMA_signal_2904, new_AGEMA_signal_2910,
         new_AGEMA_signal_2912, new_AGEMA_signal_2914, new_AGEMA_signal_2918,
         new_AGEMA_signal_2926, new_AGEMA_signal_2928, new_AGEMA_signal_2934,
         new_AGEMA_signal_2936, new_AGEMA_signal_2938, new_AGEMA_signal_2942,
         new_AGEMA_signal_2950, new_AGEMA_signal_2952, new_AGEMA_signal_2958,
         new_AGEMA_signal_2960, new_AGEMA_signal_2962, new_AGEMA_signal_2966,
         new_AGEMA_signal_2974, new_AGEMA_signal_2976, new_AGEMA_signal_2982,
         new_AGEMA_signal_2984, new_AGEMA_signal_2986, new_AGEMA_signal_2990,
         new_AGEMA_signal_2998, new_AGEMA_signal_3000, new_AGEMA_signal_3006,
         new_AGEMA_signal_3008, new_AGEMA_signal_3010, new_AGEMA_signal_3014,
         new_AGEMA_signal_3022, new_AGEMA_signal_3024, new_AGEMA_signal_3030,
         new_AGEMA_signal_3032, new_AGEMA_signal_3034, new_AGEMA_signal_3038,
         new_AGEMA_signal_3046, new_AGEMA_signal_3048, new_AGEMA_signal_3054,
         new_AGEMA_signal_3056, new_AGEMA_signal_3058, new_AGEMA_signal_3062,
         new_AGEMA_signal_3070, new_AGEMA_signal_3072, new_AGEMA_signal_3078,
         new_AGEMA_signal_3080, new_AGEMA_signal_3082, new_AGEMA_signal_3086,
         new_AGEMA_signal_3094, new_AGEMA_signal_3096, new_AGEMA_signal_3102,
         new_AGEMA_signal_3104, new_AGEMA_signal_3106, new_AGEMA_signal_3110,
         new_AGEMA_signal_3118, new_AGEMA_signal_3120, new_AGEMA_signal_3126,
         new_AGEMA_signal_3128, new_AGEMA_signal_3130, new_AGEMA_signal_3134,
         new_AGEMA_signal_3142, new_AGEMA_signal_3144, new_AGEMA_signal_3150,
         new_AGEMA_signal_3152, new_AGEMA_signal_3154, new_AGEMA_signal_3158,
         new_AGEMA_signal_3166, new_AGEMA_signal_3168, new_AGEMA_signal_3174,
         new_AGEMA_signal_3176, new_AGEMA_signal_3178, new_AGEMA_signal_3182,
         new_AGEMA_signal_3190, new_AGEMA_signal_3192, new_AGEMA_signal_3198,
         new_AGEMA_signal_3200, new_AGEMA_signal_3202, new_AGEMA_signal_3206,
         new_AGEMA_signal_3214, new_AGEMA_signal_3216, new_AGEMA_signal_3222,
         new_AGEMA_signal_3224, new_AGEMA_signal_3226, new_AGEMA_signal_3230,
         new_AGEMA_signal_3238, new_AGEMA_signal_3240, new_AGEMA_signal_3246,
         new_AGEMA_signal_3248, new_AGEMA_signal_3250, new_AGEMA_signal_3254,
         new_AGEMA_signal_3262, new_AGEMA_signal_3264, new_AGEMA_signal_3270,
         new_AGEMA_signal_3272, new_AGEMA_signal_3274, new_AGEMA_signal_3278,
         new_AGEMA_signal_3286, new_AGEMA_signal_3290, new_AGEMA_signal_3294,
         new_AGEMA_signal_3298, new_AGEMA_signal_3302, new_AGEMA_signal_3306,
         new_AGEMA_signal_3310, new_AGEMA_signal_3314, new_AGEMA_signal_3318,
         new_AGEMA_signal_3322, new_AGEMA_signal_3326, new_AGEMA_signal_3330,
         new_AGEMA_signal_3334, new_AGEMA_signal_3338, new_AGEMA_signal_3342,
         new_AGEMA_signal_3346, new_AGEMA_signal_3350, new_AGEMA_signal_3354,
         new_AGEMA_signal_3358, new_AGEMA_signal_3362, new_AGEMA_signal_3366,
         new_AGEMA_signal_3370, new_AGEMA_signal_3374, new_AGEMA_signal_3378,
         new_AGEMA_signal_3382, new_AGEMA_signal_3386, new_AGEMA_signal_3390,
         new_AGEMA_signal_3394, new_AGEMA_signal_3398, new_AGEMA_signal_3402,
         new_AGEMA_signal_3406, new_AGEMA_signal_3410, new_AGEMA_signal_3414,
         new_AGEMA_signal_3418, new_AGEMA_signal_3422, new_AGEMA_signal_3426,
         new_AGEMA_signal_3558, new_AGEMA_signal_3562, new_AGEMA_signal_3566,
         new_AGEMA_signal_3570, new_AGEMA_signal_3574, new_AGEMA_signal_3578,
         new_AGEMA_signal_3582, new_AGEMA_signal_3586, new_AGEMA_signal_3590,
         new_AGEMA_signal_3594, new_AGEMA_signal_3598, new_AGEMA_signal_3602,
         new_AGEMA_signal_3606, new_AGEMA_signal_3610, new_AGEMA_signal_3614,
         new_AGEMA_signal_3618, new_AGEMA_signal_3622, new_AGEMA_signal_3626,
         new_AGEMA_signal_3630, new_AGEMA_signal_3634, new_AGEMA_signal_3638,
         new_AGEMA_signal_3642, new_AGEMA_signal_3646, new_AGEMA_signal_3650,
         new_AGEMA_signal_3654, new_AGEMA_signal_3658, new_AGEMA_signal_3662,
         new_AGEMA_signal_3666, new_AGEMA_signal_3670, new_AGEMA_signal_3674,
         new_AGEMA_signal_3678, new_AGEMA_signal_3682, new_AGEMA_signal_3686,
         new_AGEMA_signal_3690, new_AGEMA_signal_3694, new_AGEMA_signal_3698,
         new_AGEMA_signal_3702, new_AGEMA_signal_3706, new_AGEMA_signal_3710,
         new_AGEMA_signal_3714, new_AGEMA_signal_3718, new_AGEMA_signal_3722,
         new_AGEMA_signal_3726, new_AGEMA_signal_3730, new_AGEMA_signal_3734,
         new_AGEMA_signal_3738, new_AGEMA_signal_3742, new_AGEMA_signal_3746,
         new_AGEMA_signal_3750, new_AGEMA_signal_3754, new_AGEMA_signal_3758,
         new_AGEMA_signal_3762, new_AGEMA_signal_3766, new_AGEMA_signal_3770,
         new_AGEMA_signal_3774, new_AGEMA_signal_3778, new_AGEMA_signal_3782,
         new_AGEMA_signal_3786, new_AGEMA_signal_3790, new_AGEMA_signal_3794,
         new_AGEMA_signal_3798, new_AGEMA_signal_3802, new_AGEMA_signal_3806,
         new_AGEMA_signal_3810, new_AGEMA_signal_3814, new_AGEMA_signal_3818,
         new_AGEMA_signal_3822, new_AGEMA_signal_3826, new_AGEMA_signal_3830,
         new_AGEMA_signal_3834, new_AGEMA_signal_3838, new_AGEMA_signal_3842,
         new_AGEMA_signal_3846, new_AGEMA_signal_3850, new_AGEMA_signal_3854,
         new_AGEMA_signal_3858, new_AGEMA_signal_3862, new_AGEMA_signal_3866,
         new_AGEMA_signal_3870, new_AGEMA_signal_3874, new_AGEMA_signal_3878,
         new_AGEMA_signal_3882, new_AGEMA_signal_3886, new_AGEMA_signal_3890,
         new_AGEMA_signal_3894, new_AGEMA_signal_3898, new_AGEMA_signal_3902,
         new_AGEMA_signal_3906, new_AGEMA_signal_3910, new_AGEMA_signal_3914,
         new_AGEMA_signal_3918, new_AGEMA_signal_3922, new_AGEMA_signal_3926,
         new_AGEMA_signal_3930, new_AGEMA_signal_3934, new_AGEMA_signal_3938,
         new_AGEMA_signal_3942, new_AGEMA_signal_3946, new_AGEMA_signal_3950,
         new_AGEMA_signal_3954, new_AGEMA_signal_3958, new_AGEMA_signal_3962,
         new_AGEMA_signal_3966, new_AGEMA_signal_3970, new_AGEMA_signal_3974,
         new_AGEMA_signal_3978, new_AGEMA_signal_3982, new_AGEMA_signal_3986,
         new_AGEMA_signal_3990, new_AGEMA_signal_3994, new_AGEMA_signal_3998,
         new_AGEMA_signal_4002, new_AGEMA_signal_4006, new_AGEMA_signal_4010,
         new_AGEMA_signal_4014, new_AGEMA_signal_4018, new_AGEMA_signal_4022,
         new_AGEMA_signal_4026, new_AGEMA_signal_4030, new_AGEMA_signal_4034,
         new_AGEMA_signal_4038, new_AGEMA_signal_4042, new_AGEMA_signal_4046,
         new_AGEMA_signal_4050, new_AGEMA_signal_4054, new_AGEMA_signal_4058,
         new_AGEMA_signal_4062, new_AGEMA_signal_4066, new_AGEMA_signal_4070,
         new_AGEMA_signal_4074, new_AGEMA_signal_4078, new_AGEMA_signal_4082,
         new_AGEMA_signal_4086, new_AGEMA_signal_4090, new_AGEMA_signal_2643,
         new_AGEMA_signal_2647, new_AGEMA_signal_2651, new_AGEMA_signal_2655,
         new_AGEMA_signal_2659, new_AGEMA_signal_2663, new_AGEMA_signal_2667,
         new_AGEMA_signal_2671, new_AGEMA_signal_2675, new_AGEMA_signal_2679,
         new_AGEMA_signal_2683, new_AGEMA_signal_2687, new_AGEMA_signal_2691,
         new_AGEMA_signal_2695, new_AGEMA_signal_2699, new_AGEMA_signal_2703,
         new_AGEMA_signal_2707, new_AGEMA_signal_2711, new_AGEMA_signal_2715,
         new_AGEMA_signal_2719, new_AGEMA_signal_2723, new_AGEMA_signal_2727,
         new_AGEMA_signal_2731, new_AGEMA_signal_2735, new_AGEMA_signal_2739,
         new_AGEMA_signal_2743, new_AGEMA_signal_2747, new_AGEMA_signal_2751,
         new_AGEMA_signal_2755, new_AGEMA_signal_2759, new_AGEMA_signal_2763,
         new_AGEMA_signal_2767, new_AGEMA_signal_2771, new_AGEMA_signal_2775,
         new_AGEMA_signal_2779, new_AGEMA_signal_2783, new_AGEMA_signal_2787,
         new_AGEMA_signal_2791, new_AGEMA_signal_2795, new_AGEMA_signal_2799,
         new_AGEMA_signal_2803, new_AGEMA_signal_2807, new_AGEMA_signal_2811,
         new_AGEMA_signal_2815, new_AGEMA_signal_2819, new_AGEMA_signal_2823,
         new_AGEMA_signal_2827, new_AGEMA_signal_2831, new_AGEMA_signal_2835,
         new_AGEMA_signal_2839, new_AGEMA_signal_2843, new_AGEMA_signal_2847,
         new_AGEMA_signal_2851, new_AGEMA_signal_2855, new_AGEMA_signal_2859,
         new_AGEMA_signal_2863, new_AGEMA_signal_2867, new_AGEMA_signal_2871,
         new_AGEMA_signal_2875, new_AGEMA_signal_2879, new_AGEMA_signal_2883,
         new_AGEMA_signal_2887, new_AGEMA_signal_2891, new_AGEMA_signal_2895,
         new_AGEMA_signal_2899, new_AGEMA_signal_2905, new_AGEMA_signal_2907,
         new_AGEMA_signal_2915, new_AGEMA_signal_2919, new_AGEMA_signal_2921,
         new_AGEMA_signal_2923, new_AGEMA_signal_2929, new_AGEMA_signal_2931,
         new_AGEMA_signal_2939, new_AGEMA_signal_2943, new_AGEMA_signal_2945,
         new_AGEMA_signal_2947, new_AGEMA_signal_2953, new_AGEMA_signal_2955,
         new_AGEMA_signal_2963, new_AGEMA_signal_2967, new_AGEMA_signal_2969,
         new_AGEMA_signal_2971, new_AGEMA_signal_2977, new_AGEMA_signal_2979,
         new_AGEMA_signal_2987, new_AGEMA_signal_2991, new_AGEMA_signal_2993,
         new_AGEMA_signal_2995, new_AGEMA_signal_3001, new_AGEMA_signal_3003,
         new_AGEMA_signal_3011, new_AGEMA_signal_3015, new_AGEMA_signal_3017,
         new_AGEMA_signal_3019, new_AGEMA_signal_3025, new_AGEMA_signal_3027,
         new_AGEMA_signal_3035, new_AGEMA_signal_3039, new_AGEMA_signal_3041,
         new_AGEMA_signal_3043, new_AGEMA_signal_3049, new_AGEMA_signal_3051,
         new_AGEMA_signal_3059, new_AGEMA_signal_3063, new_AGEMA_signal_3065,
         new_AGEMA_signal_3067, new_AGEMA_signal_3073, new_AGEMA_signal_3075,
         new_AGEMA_signal_3083, new_AGEMA_signal_3087, new_AGEMA_signal_3089,
         new_AGEMA_signal_3091, new_AGEMA_signal_3097, new_AGEMA_signal_3099,
         new_AGEMA_signal_3107, new_AGEMA_signal_3111, new_AGEMA_signal_3113,
         new_AGEMA_signal_3115, new_AGEMA_signal_3121, new_AGEMA_signal_3123,
         new_AGEMA_signal_3131, new_AGEMA_signal_3135, new_AGEMA_signal_3137,
         new_AGEMA_signal_3139, new_AGEMA_signal_3145, new_AGEMA_signal_3147,
         new_AGEMA_signal_3155, new_AGEMA_signal_3159, new_AGEMA_signal_3161,
         new_AGEMA_signal_3163, new_AGEMA_signal_3169, new_AGEMA_signal_3171,
         new_AGEMA_signal_3179, new_AGEMA_signal_3183, new_AGEMA_signal_3185,
         new_AGEMA_signal_3187, new_AGEMA_signal_3193, new_AGEMA_signal_3195,
         new_AGEMA_signal_3203, new_AGEMA_signal_3207, new_AGEMA_signal_3209,
         new_AGEMA_signal_3211, new_AGEMA_signal_3217, new_AGEMA_signal_3219,
         new_AGEMA_signal_3227, new_AGEMA_signal_3231, new_AGEMA_signal_3233,
         new_AGEMA_signal_3235, new_AGEMA_signal_3241, new_AGEMA_signal_3243,
         new_AGEMA_signal_3251, new_AGEMA_signal_3255, new_AGEMA_signal_3257,
         new_AGEMA_signal_3259, new_AGEMA_signal_3265, new_AGEMA_signal_3267,
         new_AGEMA_signal_3275, new_AGEMA_signal_3279, new_AGEMA_signal_3281,
         new_AGEMA_signal_3283, new_AGEMA_signal_3287, new_AGEMA_signal_3291,
         new_AGEMA_signal_3295, new_AGEMA_signal_3299, new_AGEMA_signal_3303,
         new_AGEMA_signal_3307, new_AGEMA_signal_3311, new_AGEMA_signal_3315,
         new_AGEMA_signal_3319, new_AGEMA_signal_3323, new_AGEMA_signal_3327,
         new_AGEMA_signal_3331, new_AGEMA_signal_3335, new_AGEMA_signal_3339,
         new_AGEMA_signal_3343, new_AGEMA_signal_3347, new_AGEMA_signal_3351,
         new_AGEMA_signal_3355, new_AGEMA_signal_3359, new_AGEMA_signal_3363,
         new_AGEMA_signal_3367, new_AGEMA_signal_3371, new_AGEMA_signal_3375,
         new_AGEMA_signal_3379, new_AGEMA_signal_3383, new_AGEMA_signal_3387,
         new_AGEMA_signal_3391, new_AGEMA_signal_3395, new_AGEMA_signal_3399,
         new_AGEMA_signal_3403, new_AGEMA_signal_3407, new_AGEMA_signal_3411,
         new_AGEMA_signal_3415, new_AGEMA_signal_3419, new_AGEMA_signal_3423,
         new_AGEMA_signal_3427, new_AGEMA_signal_3429, new_AGEMA_signal_3431,
         new_AGEMA_signal_3433, new_AGEMA_signal_3435, new_AGEMA_signal_3437,
         new_AGEMA_signal_3439, new_AGEMA_signal_3441, new_AGEMA_signal_3443,
         new_AGEMA_signal_3445, new_AGEMA_signal_3447, new_AGEMA_signal_3449,
         new_AGEMA_signal_3451, new_AGEMA_signal_3453, new_AGEMA_signal_3455,
         new_AGEMA_signal_3457, new_AGEMA_signal_3459, new_AGEMA_signal_3461,
         new_AGEMA_signal_3463, new_AGEMA_signal_3465, new_AGEMA_signal_3467,
         new_AGEMA_signal_3469, new_AGEMA_signal_3471, new_AGEMA_signal_3473,
         new_AGEMA_signal_3475, new_AGEMA_signal_3477, new_AGEMA_signal_3479,
         new_AGEMA_signal_3481, new_AGEMA_signal_3483, new_AGEMA_signal_3485,
         new_AGEMA_signal_3487, new_AGEMA_signal_3489, new_AGEMA_signal_3491,
         new_AGEMA_signal_3493, new_AGEMA_signal_3495, new_AGEMA_signal_3497,
         new_AGEMA_signal_3499, new_AGEMA_signal_3501, new_AGEMA_signal_3503,
         new_AGEMA_signal_3505, new_AGEMA_signal_3507, new_AGEMA_signal_3509,
         new_AGEMA_signal_3511, new_AGEMA_signal_3513, new_AGEMA_signal_3515,
         new_AGEMA_signal_3517, new_AGEMA_signal_3519, new_AGEMA_signal_3521,
         new_AGEMA_signal_3523, new_AGEMA_signal_3525, new_AGEMA_signal_3527,
         new_AGEMA_signal_3529, new_AGEMA_signal_3531, new_AGEMA_signal_3533,
         new_AGEMA_signal_3535, new_AGEMA_signal_3537, new_AGEMA_signal_3539,
         new_AGEMA_signal_3541, new_AGEMA_signal_3543, new_AGEMA_signal_3545,
         new_AGEMA_signal_3547, new_AGEMA_signal_3549, new_AGEMA_signal_3551,
         new_AGEMA_signal_3553, new_AGEMA_signal_3555, new_AGEMA_signal_3559,
         new_AGEMA_signal_3563, new_AGEMA_signal_3567, new_AGEMA_signal_3571,
         new_AGEMA_signal_3575, new_AGEMA_signal_3579, new_AGEMA_signal_3583,
         new_AGEMA_signal_3587, new_AGEMA_signal_3591, new_AGEMA_signal_3595,
         new_AGEMA_signal_3599, new_AGEMA_signal_3603, new_AGEMA_signal_3607,
         new_AGEMA_signal_3611, new_AGEMA_signal_3615, new_AGEMA_signal_3619,
         new_AGEMA_signal_3623, new_AGEMA_signal_3627, new_AGEMA_signal_3631,
         new_AGEMA_signal_3635, new_AGEMA_signal_3639, new_AGEMA_signal_3643,
         new_AGEMA_signal_3647, new_AGEMA_signal_3651, new_AGEMA_signal_3655,
         new_AGEMA_signal_3659, new_AGEMA_signal_3663, new_AGEMA_signal_3667,
         new_AGEMA_signal_3671, new_AGEMA_signal_3675, new_AGEMA_signal_3679,
         new_AGEMA_signal_3683, new_AGEMA_signal_3687, new_AGEMA_signal_3691,
         new_AGEMA_signal_3695, new_AGEMA_signal_3699, new_AGEMA_signal_3703,
         new_AGEMA_signal_3707, new_AGEMA_signal_3711, new_AGEMA_signal_3715,
         new_AGEMA_signal_3719, new_AGEMA_signal_3723, new_AGEMA_signal_3727,
         new_AGEMA_signal_3731, new_AGEMA_signal_3735, new_AGEMA_signal_3739,
         new_AGEMA_signal_3743, new_AGEMA_signal_3747, new_AGEMA_signal_3751,
         new_AGEMA_signal_3755, new_AGEMA_signal_3759, new_AGEMA_signal_3763,
         new_AGEMA_signal_3767, new_AGEMA_signal_3771, new_AGEMA_signal_3775,
         new_AGEMA_signal_3779, new_AGEMA_signal_3783, new_AGEMA_signal_3787,
         new_AGEMA_signal_3791, new_AGEMA_signal_3795, new_AGEMA_signal_3799,
         new_AGEMA_signal_3803, new_AGEMA_signal_3807, new_AGEMA_signal_3811,
         new_AGEMA_signal_3815, new_AGEMA_signal_3819, new_AGEMA_signal_3823,
         new_AGEMA_signal_3827, new_AGEMA_signal_3831, new_AGEMA_signal_3835,
         new_AGEMA_signal_3839, new_AGEMA_signal_3843, new_AGEMA_signal_3847,
         new_AGEMA_signal_3851, new_AGEMA_signal_3855, new_AGEMA_signal_3859,
         new_AGEMA_signal_3863, new_AGEMA_signal_3867, new_AGEMA_signal_3871,
         new_AGEMA_signal_3875, new_AGEMA_signal_3879, new_AGEMA_signal_3883,
         new_AGEMA_signal_3887, new_AGEMA_signal_3891, new_AGEMA_signal_3895,
         new_AGEMA_signal_3899, new_AGEMA_signal_3903, new_AGEMA_signal_3907,
         new_AGEMA_signal_3911, new_AGEMA_signal_3915, new_AGEMA_signal_3919,
         new_AGEMA_signal_3923, new_AGEMA_signal_3927, new_AGEMA_signal_3931,
         new_AGEMA_signal_3935, new_AGEMA_signal_3939, new_AGEMA_signal_3943,
         new_AGEMA_signal_3947, new_AGEMA_signal_3951, new_AGEMA_signal_3955,
         new_AGEMA_signal_3959, new_AGEMA_signal_3963, new_AGEMA_signal_3967,
         new_AGEMA_signal_3971, new_AGEMA_signal_3975, new_AGEMA_signal_3979,
         new_AGEMA_signal_3983, new_AGEMA_signal_3987, new_AGEMA_signal_3991,
         new_AGEMA_signal_3995, new_AGEMA_signal_3999, new_AGEMA_signal_4003,
         new_AGEMA_signal_4007, new_AGEMA_signal_4011, new_AGEMA_signal_4015,
         new_AGEMA_signal_4019, new_AGEMA_signal_4023, new_AGEMA_signal_4027,
         new_AGEMA_signal_4031, new_AGEMA_signal_4035, new_AGEMA_signal_4039,
         new_AGEMA_signal_4043, new_AGEMA_signal_4047, new_AGEMA_signal_4051,
         new_AGEMA_signal_4055, new_AGEMA_signal_4059, new_AGEMA_signal_4063,
         new_AGEMA_signal_4067, new_AGEMA_signal_4071, new_AGEMA_signal_4075,
         new_AGEMA_signal_4079, new_AGEMA_signal_4083, new_AGEMA_signal_4087,
         new_AGEMA_signal_4091, new_AGEMA_signal_2644, new_AGEMA_signal_2036,
         new_AGEMA_signal_2652, new_AGEMA_signal_2648, new_AGEMA_signal_2027,
         new_AGEMA_signal_2079, new_AGEMA_signal_2660, new_AGEMA_signal_2656,
         new_AGEMA_signal_2073, new_AGEMA_signal_2038, new_AGEMA_signal_2668,
         new_AGEMA_signal_2664, new_AGEMA_signal_2029, new_AGEMA_signal_2081,
         new_AGEMA_signal_2676, new_AGEMA_signal_2672, new_AGEMA_signal_2074,
         new_AGEMA_signal_2040, new_AGEMA_signal_2684, new_AGEMA_signal_2680,
         new_AGEMA_signal_2031, new_AGEMA_signal_2083, new_AGEMA_signal_2692,
         new_AGEMA_signal_2688, new_AGEMA_signal_2075, new_AGEMA_signal_2111,
         new_AGEMA_signal_2700, new_AGEMA_signal_2696, new_AGEMA_signal_2108,
         new_AGEMA_signal_2120, new_AGEMA_signal_2708, new_AGEMA_signal_2704,
         new_AGEMA_signal_2118, new_AGEMA_signal_2044, new_AGEMA_signal_2716,
         new_AGEMA_signal_2712, new_AGEMA_signal_2019, new_AGEMA_signal_2087,
         new_AGEMA_signal_2724, new_AGEMA_signal_2720, new_AGEMA_signal_2068,
         new_AGEMA_signal_2046, new_AGEMA_signal_2732, new_AGEMA_signal_2728,
         new_AGEMA_signal_2021, new_AGEMA_signal_2089, new_AGEMA_signal_2740,
         new_AGEMA_signal_2736, new_AGEMA_signal_2069, new_AGEMA_signal_2113,
         new_AGEMA_signal_2748, new_AGEMA_signal_2744, new_AGEMA_signal_2106,
         new_AGEMA_signal_2122, new_AGEMA_signal_2756, new_AGEMA_signal_2752,
         new_AGEMA_signal_2117, new_AGEMA_signal_2050, new_AGEMA_signal_2764,
         new_AGEMA_signal_2760, new_AGEMA_signal_2025, new_AGEMA_signal_2093,
         new_AGEMA_signal_2772, new_AGEMA_signal_2768, new_AGEMA_signal_2072,
         new_AGEMA_signal_1934, new_AGEMA_signal_2780, new_AGEMA_signal_2776,
         new_AGEMA_signal_1892, new_AGEMA_signal_1994, new_AGEMA_signal_2788,
         new_AGEMA_signal_2784, new_AGEMA_signal_1954, new_AGEMA_signal_1936,
         new_AGEMA_signal_2796, new_AGEMA_signal_2792, new_AGEMA_signal_1894,
         new_AGEMA_signal_1996, new_AGEMA_signal_2804, new_AGEMA_signal_2800,
         new_AGEMA_signal_1955, new_AGEMA_signal_1938, new_AGEMA_signal_2812,
         new_AGEMA_signal_2808, new_AGEMA_signal_1896, new_AGEMA_signal_1998,
         new_AGEMA_signal_2820, new_AGEMA_signal_2816, new_AGEMA_signal_1956,
         new_AGEMA_signal_2052, new_AGEMA_signal_2828, new_AGEMA_signal_2824,
         new_AGEMA_signal_2009, new_AGEMA_signal_2095, new_AGEMA_signal_2836,
         new_AGEMA_signal_2832, new_AGEMA_signal_2062, new_AGEMA_signal_2054,
         new_AGEMA_signal_2844, new_AGEMA_signal_2840, new_AGEMA_signal_2011,
         new_AGEMA_signal_2097, new_AGEMA_signal_2852, new_AGEMA_signal_2848,
         new_AGEMA_signal_2063, new_AGEMA_signal_2056, new_AGEMA_signal_2860,
         new_AGEMA_signal_2856, new_AGEMA_signal_2013, new_AGEMA_signal_2099,
         new_AGEMA_signal_2868, new_AGEMA_signal_2864, new_AGEMA_signal_2064,
         new_AGEMA_signal_2058, new_AGEMA_signal_2876, new_AGEMA_signal_2872,
         new_AGEMA_signal_2015, new_AGEMA_signal_2101, new_AGEMA_signal_2884,
         new_AGEMA_signal_2880, new_AGEMA_signal_2065, new_AGEMA_signal_2115,
         new_AGEMA_signal_2892, new_AGEMA_signal_2888, new_AGEMA_signal_2104,
         new_AGEMA_signal_2124, new_AGEMA_signal_2900, new_AGEMA_signal_2896,
         new_AGEMA_signal_2116, new_AGEMA_signal_1661,
         SubCellInst_SboxInst_0_T1, new_AGEMA_signal_1725,
         SubCellInst_SboxInst_0_L0, new_AGEMA_signal_2908,
         new_AGEMA_signal_2906, new_AGEMA_signal_1662,
         SubCellInst_SboxInst_0_T3, new_AGEMA_signal_1768,
         SubCellInst_SboxInst_0_YY_3, new_AGEMA_signal_2920,
         new_AGEMA_signal_2916, new_AGEMA_signal_1769, new_AGEMA_signal_1826,
         new_AGEMA_signal_2924, new_AGEMA_signal_2922, new_AGEMA_signal_1665,
         SubCellInst_SboxInst_1_T1, new_AGEMA_signal_1727,
         SubCellInst_SboxInst_1_L0, new_AGEMA_signal_2932,
         new_AGEMA_signal_2930, new_AGEMA_signal_1666,
         SubCellInst_SboxInst_1_T3, new_AGEMA_signal_1770,
         SubCellInst_SboxInst_1_YY_3, new_AGEMA_signal_2944,
         new_AGEMA_signal_2940, new_AGEMA_signal_1771, new_AGEMA_signal_1827,
         new_AGEMA_signal_2948, new_AGEMA_signal_2946, new_AGEMA_signal_1669,
         SubCellInst_SboxInst_2_T1, new_AGEMA_signal_1729,
         SubCellInst_SboxInst_2_L0, new_AGEMA_signal_2956,
         new_AGEMA_signal_2954, new_AGEMA_signal_1670,
         SubCellInst_SboxInst_2_T3, new_AGEMA_signal_1772,
         SubCellInst_SboxInst_2_YY_3, new_AGEMA_signal_2968,
         new_AGEMA_signal_2964, new_AGEMA_signal_1773, new_AGEMA_signal_1828,
         new_AGEMA_signal_2972, new_AGEMA_signal_2970, new_AGEMA_signal_1673,
         SubCellInst_SboxInst_3_T1, new_AGEMA_signal_1731,
         SubCellInst_SboxInst_3_L0, new_AGEMA_signal_2980,
         new_AGEMA_signal_2978, new_AGEMA_signal_1674,
         SubCellInst_SboxInst_3_T3, new_AGEMA_signal_1774,
         SubCellInst_SboxInst_3_YY_3, new_AGEMA_signal_2992,
         new_AGEMA_signal_2988, new_AGEMA_signal_1775, new_AGEMA_signal_1829,
         new_AGEMA_signal_2996, new_AGEMA_signal_2994, new_AGEMA_signal_1677,
         SubCellInst_SboxInst_4_T1, new_AGEMA_signal_1733,
         SubCellInst_SboxInst_4_L0, new_AGEMA_signal_3004,
         new_AGEMA_signal_3002, new_AGEMA_signal_1678,
         SubCellInst_SboxInst_4_T3, new_AGEMA_signal_1776,
         SubCellInst_SboxInst_4_YY_3, new_AGEMA_signal_3016,
         new_AGEMA_signal_3012, new_AGEMA_signal_1777, new_AGEMA_signal_1830,
         new_AGEMA_signal_3020, new_AGEMA_signal_3018, new_AGEMA_signal_1681,
         SubCellInst_SboxInst_5_T1, new_AGEMA_signal_1735,
         SubCellInst_SboxInst_5_L0, new_AGEMA_signal_3028,
         new_AGEMA_signal_3026, new_AGEMA_signal_1682,
         SubCellInst_SboxInst_5_T3, new_AGEMA_signal_1778,
         SubCellInst_SboxInst_5_YY_3, new_AGEMA_signal_3040,
         new_AGEMA_signal_3036, new_AGEMA_signal_1779, new_AGEMA_signal_1831,
         new_AGEMA_signal_3044, new_AGEMA_signal_3042, new_AGEMA_signal_1685,
         SubCellInst_SboxInst_6_T1, new_AGEMA_signal_1737,
         SubCellInst_SboxInst_6_L0, new_AGEMA_signal_3052,
         new_AGEMA_signal_3050, new_AGEMA_signal_1686,
         SubCellInst_SboxInst_6_T3, new_AGEMA_signal_1780,
         SubCellInst_SboxInst_6_YY_3, new_AGEMA_signal_3064,
         new_AGEMA_signal_3060, new_AGEMA_signal_1781, new_AGEMA_signal_1832,
         new_AGEMA_signal_3068, new_AGEMA_signal_3066, new_AGEMA_signal_1689,
         SubCellInst_SboxInst_7_T1, new_AGEMA_signal_1739,
         SubCellInst_SboxInst_7_L0, new_AGEMA_signal_3076,
         new_AGEMA_signal_3074, new_AGEMA_signal_1690,
         SubCellInst_SboxInst_7_T3, new_AGEMA_signal_1782,
         SubCellInst_SboxInst_7_YY_3, new_AGEMA_signal_3088,
         new_AGEMA_signal_3084, new_AGEMA_signal_1783, new_AGEMA_signal_3092,
         new_AGEMA_signal_3090, new_AGEMA_signal_1693,
         SubCellInst_SboxInst_8_T1, new_AGEMA_signal_1741,
         SubCellInst_SboxInst_8_L0, new_AGEMA_signal_3100,
         new_AGEMA_signal_3098, new_AGEMA_signal_1694,
         SubCellInst_SboxInst_8_T3, new_AGEMA_signal_1784,
         SubCellInst_SboxInst_8_YY_3, new_AGEMA_signal_3112,
         new_AGEMA_signal_3108, new_AGEMA_signal_1785, new_AGEMA_signal_1834,
         new_AGEMA_signal_3116, new_AGEMA_signal_3114, new_AGEMA_signal_1697,
         SubCellInst_SboxInst_9_T1, new_AGEMA_signal_1743,
         SubCellInst_SboxInst_9_L0, new_AGEMA_signal_3124,
         new_AGEMA_signal_3122, new_AGEMA_signal_1698,
         SubCellInst_SboxInst_9_T3, new_AGEMA_signal_1786,
         SubCellInst_SboxInst_9_YY_3, new_AGEMA_signal_3136,
         new_AGEMA_signal_3132, new_AGEMA_signal_1787, new_AGEMA_signal_1835,
         new_AGEMA_signal_3140, new_AGEMA_signal_3138, new_AGEMA_signal_1701,
         SubCellInst_SboxInst_10_T1, new_AGEMA_signal_1745,
         SubCellInst_SboxInst_10_L0, new_AGEMA_signal_3148,
         new_AGEMA_signal_3146, new_AGEMA_signal_1702,
         SubCellInst_SboxInst_10_T3, new_AGEMA_signal_1788,
         SubCellInst_SboxInst_10_YY_3, new_AGEMA_signal_3160,
         new_AGEMA_signal_3156, new_AGEMA_signal_1789, new_AGEMA_signal_1836,
         new_AGEMA_signal_3164, new_AGEMA_signal_3162, new_AGEMA_signal_1705,
         SubCellInst_SboxInst_11_T1, new_AGEMA_signal_1747,
         SubCellInst_SboxInst_11_L0, new_AGEMA_signal_3172,
         new_AGEMA_signal_3170, new_AGEMA_signal_1706,
         SubCellInst_SboxInst_11_T3, new_AGEMA_signal_1790,
         SubCellInst_SboxInst_11_YY_3, new_AGEMA_signal_3184,
         new_AGEMA_signal_3180, new_AGEMA_signal_1791, new_AGEMA_signal_1837,
         new_AGEMA_signal_3188, new_AGEMA_signal_3186, new_AGEMA_signal_1709,
         SubCellInst_SboxInst_12_T1, new_AGEMA_signal_1749,
         SubCellInst_SboxInst_12_L0, new_AGEMA_signal_3196,
         new_AGEMA_signal_3194, new_AGEMA_signal_1710,
         SubCellInst_SboxInst_12_T3, new_AGEMA_signal_1792,
         SubCellInst_SboxInst_12_YY_3, new_AGEMA_signal_3208,
         new_AGEMA_signal_3204, new_AGEMA_signal_1793, new_AGEMA_signal_1838,
         new_AGEMA_signal_3212, new_AGEMA_signal_3210, new_AGEMA_signal_1713,
         SubCellInst_SboxInst_13_T1, new_AGEMA_signal_1751,
         SubCellInst_SboxInst_13_L0, new_AGEMA_signal_3220,
         new_AGEMA_signal_3218, new_AGEMA_signal_1714,
         SubCellInst_SboxInst_13_T3, new_AGEMA_signal_1794,
         SubCellInst_SboxInst_13_YY_3, new_AGEMA_signal_3232,
         new_AGEMA_signal_3228, new_AGEMA_signal_1795, new_AGEMA_signal_1839,
         new_AGEMA_signal_3236, new_AGEMA_signal_3234, new_AGEMA_signal_1717,
         SubCellInst_SboxInst_14_T1, new_AGEMA_signal_1753,
         SubCellInst_SboxInst_14_L0, new_AGEMA_signal_3244,
         new_AGEMA_signal_3242, new_AGEMA_signal_1718,
         SubCellInst_SboxInst_14_T3, new_AGEMA_signal_1796,
         SubCellInst_SboxInst_14_YY_3, new_AGEMA_signal_3256,
         new_AGEMA_signal_3252, new_AGEMA_signal_1797, new_AGEMA_signal_1840,
         new_AGEMA_signal_3260, new_AGEMA_signal_3258, new_AGEMA_signal_1721,
         SubCellInst_SboxInst_15_T1, new_AGEMA_signal_1755,
         SubCellInst_SboxInst_15_L0, new_AGEMA_signal_3268,
         new_AGEMA_signal_3266, new_AGEMA_signal_1722,
         SubCellInst_SboxInst_15_T3, new_AGEMA_signal_1798,
         SubCellInst_SboxInst_15_YY_3, new_AGEMA_signal_3280,
         new_AGEMA_signal_3276, new_AGEMA_signal_1799, new_AGEMA_signal_1841,
         new_AGEMA_signal_3284, new_AGEMA_signal_3282, new_AGEMA_signal_1879,
         new_AGEMA_signal_1880, new_AGEMA_signal_3288, new_AGEMA_signal_1842,
         AddConstXOR_AddConstXOR_XORInst_0_0_n1, new_AGEMA_signal_1947,
         new_AGEMA_signal_3292, new_AGEMA_signal_1881,
         AddConstXOR_AddConstXOR_XORInst_0_1_n1, new_AGEMA_signal_1882,
         new_AGEMA_signal_3296, new_AGEMA_signal_1844,
         AddConstXOR_AddConstXOR_XORInst_1_0_n1, new_AGEMA_signal_1948,
         new_AGEMA_signal_3300, new_AGEMA_signal_1883,
         AddConstXOR_AddConstXOR_XORInst_1_1_n1, new_AGEMA_signal_1884,
         new_AGEMA_signal_3308, new_AGEMA_signal_3304, new_AGEMA_signal_1846,
         AddRoundTweakeyXOR_XORInst_0_0_n1, new_AGEMA_signal_1949,
         new_AGEMA_signal_3316, new_AGEMA_signal_3312, new_AGEMA_signal_1885,
         AddRoundTweakeyXOR_XORInst_0_1_n1, new_AGEMA_signal_1886,
         new_AGEMA_signal_3324, new_AGEMA_signal_3320, new_AGEMA_signal_1848,
         AddRoundTweakeyXOR_XORInst_1_0_n1, new_AGEMA_signal_1950,
         new_AGEMA_signal_3332, new_AGEMA_signal_3328, new_AGEMA_signal_1887,
         AddRoundTweakeyXOR_XORInst_1_1_n1, new_AGEMA_signal_1888,
         new_AGEMA_signal_3340, new_AGEMA_signal_3336, new_AGEMA_signal_1850,
         AddRoundTweakeyXOR_XORInst_2_0_n1, new_AGEMA_signal_1951,
         new_AGEMA_signal_3348, new_AGEMA_signal_3344, new_AGEMA_signal_1889,
         AddRoundTweakeyXOR_XORInst_2_1_n1, new_AGEMA_signal_2007,
         new_AGEMA_signal_3356, new_AGEMA_signal_3352, new_AGEMA_signal_1952,
         AddRoundTweakeyXOR_XORInst_3_0_n1, new_AGEMA_signal_2061,
         new_AGEMA_signal_3364, new_AGEMA_signal_3360, new_AGEMA_signal_2008,
         AddRoundTweakeyXOR_XORInst_3_1_n1, new_AGEMA_signal_3372,
         new_AGEMA_signal_3368, new_AGEMA_signal_1853,
         AddRoundTweakeyXOR_XORInst_4_0_n1, new_AGEMA_signal_3380,
         new_AGEMA_signal_3376, new_AGEMA_signal_1893,
         AddRoundTweakeyXOR_XORInst_4_1_n1, new_AGEMA_signal_3388,
         new_AGEMA_signal_3384, new_AGEMA_signal_1855,
         AddRoundTweakeyXOR_XORInst_5_0_n1, new_AGEMA_signal_3396,
         new_AGEMA_signal_3392, new_AGEMA_signal_1895,
         AddRoundTweakeyXOR_XORInst_5_1_n1, new_AGEMA_signal_3404,
         new_AGEMA_signal_3400, new_AGEMA_signal_1857,
         AddRoundTweakeyXOR_XORInst_6_0_n1, new_AGEMA_signal_3412,
         new_AGEMA_signal_3408, new_AGEMA_signal_1897,
         AddRoundTweakeyXOR_XORInst_6_1_n1, new_AGEMA_signal_3420,
         new_AGEMA_signal_3416, new_AGEMA_signal_1957,
         AddRoundTweakeyXOR_XORInst_7_0_n1, new_AGEMA_signal_3428,
         new_AGEMA_signal_3424, new_AGEMA_signal_2010,
         AddRoundTweakeyXOR_XORInst_7_1_n1, new_AGEMA_signal_1860,
         MCInst_MCR0_XORInst_0_0_n1, new_AGEMA_signal_1959,
         MCInst_MCR0_XORInst_0_0_n2, new_AGEMA_signal_1900,
         MCInst_MCR0_XORInst_0_1_n1, new_AGEMA_signal_2012,
         MCInst_MCR0_XORInst_0_1_n2, new_AGEMA_signal_1862,
         MCInst_MCR0_XORInst_1_0_n1, new_AGEMA_signal_1961,
         MCInst_MCR0_XORInst_1_0_n2, new_AGEMA_signal_1962,
         MCInst_MCR0_XORInst_1_1_n1, new_AGEMA_signal_2014,
         MCInst_MCR0_XORInst_1_1_n2, new_AGEMA_signal_1864,
         MCInst_MCR0_XORInst_2_0_n1, new_AGEMA_signal_1964,
         MCInst_MCR0_XORInst_2_0_n2, new_AGEMA_signal_1905,
         MCInst_MCR0_XORInst_2_1_n1, new_AGEMA_signal_2016,
         MCInst_MCR0_XORInst_2_1_n2, new_AGEMA_signal_1866,
         MCInst_MCR0_XORInst_3_0_n1, new_AGEMA_signal_2066,
         MCInst_MCR0_XORInst_3_0_n2, new_AGEMA_signal_1908,
         MCInst_MCR0_XORInst_3_1_n1, new_AGEMA_signal_2105,
         MCInst_MCR0_XORInst_3_1_n2, new_AGEMA_signal_1967,
         MCInst_MCR2_XORInst_0_0_n1, new_AGEMA_signal_2020,
         MCInst_MCR2_XORInst_0_1_n1, new_AGEMA_signal_1969,
         MCInst_MCR2_XORInst_1_0_n1, new_AGEMA_signal_2022,
         MCInst_MCR2_XORInst_1_1_n1, new_AGEMA_signal_2070,
         MCInst_MCR2_XORInst_2_0_n1, new_AGEMA_signal_2107,
         MCInst_MCR2_XORInst_2_1_n1, new_AGEMA_signal_1972,
         MCInst_MCR2_XORInst_3_0_n1, new_AGEMA_signal_2026,
         MCInst_MCR2_XORInst_3_1_n1, new_AGEMA_signal_1974,
         MCInst_MCR3_XORInst_0_0_n1, new_AGEMA_signal_2028,
         MCInst_MCR3_XORInst_0_1_n1, new_AGEMA_signal_1976,
         MCInst_MCR3_XORInst_1_0_n1, new_AGEMA_signal_2030,
         MCInst_MCR3_XORInst_1_1_n1, new_AGEMA_signal_1978,
         MCInst_MCR3_XORInst_2_0_n1, new_AGEMA_signal_2032,
         MCInst_MCR3_XORInst_2_1_n1, new_AGEMA_signal_2076,
         MCInst_MCR3_XORInst_3_0_n1, new_AGEMA_signal_2109,
         MCInst_MCR3_XORInst_3_1_n1, new_AGEMA_signal_3430,
         new_AGEMA_signal_3432, new_AGEMA_signal_3434, new_AGEMA_signal_3436,
         new_AGEMA_signal_3438, new_AGEMA_signal_3440, new_AGEMA_signal_3442,
         new_AGEMA_signal_3444, new_AGEMA_signal_3446, new_AGEMA_signal_3448,
         new_AGEMA_signal_3450, new_AGEMA_signal_3452, new_AGEMA_signal_3454,
         new_AGEMA_signal_3456, new_AGEMA_signal_3458, new_AGEMA_signal_3460,
         new_AGEMA_signal_3462, new_AGEMA_signal_3464, new_AGEMA_signal_3466,
         new_AGEMA_signal_3468, new_AGEMA_signal_3470, new_AGEMA_signal_3472,
         new_AGEMA_signal_3474, new_AGEMA_signal_3476, new_AGEMA_signal_3478,
         new_AGEMA_signal_3480, new_AGEMA_signal_3482, new_AGEMA_signal_3484,
         new_AGEMA_signal_3486, new_AGEMA_signal_3488, new_AGEMA_signal_3490,
         new_AGEMA_signal_3492, new_AGEMA_signal_3494, new_AGEMA_signal_3496,
         new_AGEMA_signal_3498, new_AGEMA_signal_3500, new_AGEMA_signal_3502,
         new_AGEMA_signal_3504, new_AGEMA_signal_3506, new_AGEMA_signal_3508,
         new_AGEMA_signal_3510, new_AGEMA_signal_3512, new_AGEMA_signal_3514,
         new_AGEMA_signal_3516, new_AGEMA_signal_3518, new_AGEMA_signal_3520,
         new_AGEMA_signal_3522, new_AGEMA_signal_3524, new_AGEMA_signal_3526,
         new_AGEMA_signal_3528, new_AGEMA_signal_3530, new_AGEMA_signal_3532,
         new_AGEMA_signal_3534, new_AGEMA_signal_3536, new_AGEMA_signal_3538,
         new_AGEMA_signal_3540, new_AGEMA_signal_3542, new_AGEMA_signal_3544,
         new_AGEMA_signal_3546, new_AGEMA_signal_3548, new_AGEMA_signal_3550,
         new_AGEMA_signal_3552, new_AGEMA_signal_3554, new_AGEMA_signal_3556,
         new_AGEMA_signal_3560, new_AGEMA_signal_3564, new_AGEMA_signal_3568,
         new_AGEMA_signal_3572, new_AGEMA_signal_3576, new_AGEMA_signal_3580,
         new_AGEMA_signal_3584, new_AGEMA_signal_3588, new_AGEMA_signal_3592,
         new_AGEMA_signal_3596, new_AGEMA_signal_3600, new_AGEMA_signal_3604,
         new_AGEMA_signal_3608, new_AGEMA_signal_3612, new_AGEMA_signal_3616,
         new_AGEMA_signal_3620, new_AGEMA_signal_3624, new_AGEMA_signal_3628,
         new_AGEMA_signal_3632, new_AGEMA_signal_3636, new_AGEMA_signal_3640,
         new_AGEMA_signal_3644, new_AGEMA_signal_3648, new_AGEMA_signal_3652,
         new_AGEMA_signal_3656, new_AGEMA_signal_3660, new_AGEMA_signal_3664,
         new_AGEMA_signal_3668, new_AGEMA_signal_3672, new_AGEMA_signal_3676,
         new_AGEMA_signal_3680, new_AGEMA_signal_3684, new_AGEMA_signal_3688,
         new_AGEMA_signal_3692, new_AGEMA_signal_3696, new_AGEMA_signal_3700,
         new_AGEMA_signal_3704, new_AGEMA_signal_3708, new_AGEMA_signal_3712,
         new_AGEMA_signal_3716, new_AGEMA_signal_3720, new_AGEMA_signal_3724,
         new_AGEMA_signal_3728, new_AGEMA_signal_3732, new_AGEMA_signal_3736,
         new_AGEMA_signal_3740, new_AGEMA_signal_3744, new_AGEMA_signal_3748,
         new_AGEMA_signal_3752, new_AGEMA_signal_3756, new_AGEMA_signal_3760,
         new_AGEMA_signal_3764, new_AGEMA_signal_3768, new_AGEMA_signal_3772,
         new_AGEMA_signal_3776, new_AGEMA_signal_3780, new_AGEMA_signal_3784,
         new_AGEMA_signal_3788, new_AGEMA_signal_3792, new_AGEMA_signal_3796,
         new_AGEMA_signal_3800, new_AGEMA_signal_3804, new_AGEMA_signal_3808,
         new_AGEMA_signal_3812, new_AGEMA_signal_3816, new_AGEMA_signal_3820,
         new_AGEMA_signal_3824, new_AGEMA_signal_3828, new_AGEMA_signal_3832,
         new_AGEMA_signal_3836, new_AGEMA_signal_3840, new_AGEMA_signal_3844,
         new_AGEMA_signal_3848, new_AGEMA_signal_3852, new_AGEMA_signal_3856,
         new_AGEMA_signal_3860, new_AGEMA_signal_3864, new_AGEMA_signal_3868,
         new_AGEMA_signal_3872, new_AGEMA_signal_3876, new_AGEMA_signal_3880,
         new_AGEMA_signal_3884, new_AGEMA_signal_3888, new_AGEMA_signal_3892,
         new_AGEMA_signal_3896, new_AGEMA_signal_3900, new_AGEMA_signal_3904,
         new_AGEMA_signal_3908, new_AGEMA_signal_3912, new_AGEMA_signal_3916,
         new_AGEMA_signal_3920, new_AGEMA_signal_3924, new_AGEMA_signal_3928,
         new_AGEMA_signal_3932, new_AGEMA_signal_3936, new_AGEMA_signal_3940,
         new_AGEMA_signal_3944, new_AGEMA_signal_3948, new_AGEMA_signal_3952,
         new_AGEMA_signal_3956, new_AGEMA_signal_3960, new_AGEMA_signal_3964,
         new_AGEMA_signal_3968, new_AGEMA_signal_3972, new_AGEMA_signal_3976,
         new_AGEMA_signal_3980, new_AGEMA_signal_3984, new_AGEMA_signal_3988,
         new_AGEMA_signal_3992, new_AGEMA_signal_3996, new_AGEMA_signal_4000,
         new_AGEMA_signal_4004, new_AGEMA_signal_4008, new_AGEMA_signal_4012,
         new_AGEMA_signal_4016, new_AGEMA_signal_4020, new_AGEMA_signal_4024,
         new_AGEMA_signal_4028, new_AGEMA_signal_4032, new_AGEMA_signal_4036,
         new_AGEMA_signal_4040, new_AGEMA_signal_4044, new_AGEMA_signal_4048,
         new_AGEMA_signal_4052, new_AGEMA_signal_4056, new_AGEMA_signal_4060,
         new_AGEMA_signal_4064, new_AGEMA_signal_4068, new_AGEMA_signal_4072,
         new_AGEMA_signal_4076, new_AGEMA_signal_4080, new_AGEMA_signal_4084,
         new_AGEMA_signal_4088, new_AGEMA_signal_4092, n13, n14, n15, n16, n17,
         n18, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, SubCellInst_SboxInst_0_AND1_U1_n9,
         SubCellInst_SboxInst_0_AND1_U1_n8, SubCellInst_SboxInst_0_AND1_U1_n7,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_0_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_0_AND3_U1_n9, SubCellInst_SboxInst_0_AND3_U1_n8,
         SubCellInst_SboxInst_0_AND3_U1_n7,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_0_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_1_AND1_U1_n9, SubCellInst_SboxInst_1_AND1_U1_n8,
         SubCellInst_SboxInst_1_AND1_U1_n7,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_1_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_1_AND3_U1_n9, SubCellInst_SboxInst_1_AND3_U1_n8,
         SubCellInst_SboxInst_1_AND3_U1_n7,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_1_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_2_AND1_U1_n9, SubCellInst_SboxInst_2_AND1_U1_n8,
         SubCellInst_SboxInst_2_AND1_U1_n7,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_2_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_2_AND3_U1_n9, SubCellInst_SboxInst_2_AND3_U1_n8,
         SubCellInst_SboxInst_2_AND3_U1_n7,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_2_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_3_AND1_U1_n9, SubCellInst_SboxInst_3_AND1_U1_n8,
         SubCellInst_SboxInst_3_AND1_U1_n7,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_3_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_3_AND3_U1_n9, SubCellInst_SboxInst_3_AND3_U1_n8,
         SubCellInst_SboxInst_3_AND3_U1_n7,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_3_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_4_AND1_U1_n9, SubCellInst_SboxInst_4_AND1_U1_n8,
         SubCellInst_SboxInst_4_AND1_U1_n7,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_4_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_4_AND3_U1_n9, SubCellInst_SboxInst_4_AND3_U1_n8,
         SubCellInst_SboxInst_4_AND3_U1_n7,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_4_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_5_AND1_U1_n9, SubCellInst_SboxInst_5_AND1_U1_n8,
         SubCellInst_SboxInst_5_AND1_U1_n7,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_5_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_5_AND3_U1_n9, SubCellInst_SboxInst_5_AND3_U1_n8,
         SubCellInst_SboxInst_5_AND3_U1_n7,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_5_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_6_AND1_U1_n9, SubCellInst_SboxInst_6_AND1_U1_n8,
         SubCellInst_SboxInst_6_AND1_U1_n7,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_6_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_6_AND3_U1_n9, SubCellInst_SboxInst_6_AND3_U1_n8,
         SubCellInst_SboxInst_6_AND3_U1_n7,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_6_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_7_AND1_U1_n9, SubCellInst_SboxInst_7_AND1_U1_n8,
         SubCellInst_SboxInst_7_AND1_U1_n7,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_7_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_7_AND3_U1_n9, SubCellInst_SboxInst_7_AND3_U1_n8,
         SubCellInst_SboxInst_7_AND3_U1_n7,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_7_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_8_AND1_U1_n9, SubCellInst_SboxInst_8_AND1_U1_n8,
         SubCellInst_SboxInst_8_AND1_U1_n7,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_8_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_8_AND3_U1_n9, SubCellInst_SboxInst_8_AND3_U1_n8,
         SubCellInst_SboxInst_8_AND3_U1_n7,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_8_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_9_AND1_U1_n9, SubCellInst_SboxInst_9_AND1_U1_n8,
         SubCellInst_SboxInst_9_AND1_U1_n7,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_9_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_9_AND3_U1_n9, SubCellInst_SboxInst_9_AND3_U1_n8,
         SubCellInst_SboxInst_9_AND3_U1_n7,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_9_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_10_AND1_U1_n9,
         SubCellInst_SboxInst_10_AND1_U1_n8,
         SubCellInst_SboxInst_10_AND1_U1_n7,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_10_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_10_AND3_U1_n9,
         SubCellInst_SboxInst_10_AND3_U1_n8,
         SubCellInst_SboxInst_10_AND3_U1_n7,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_10_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_11_AND1_U1_n9,
         SubCellInst_SboxInst_11_AND1_U1_n8,
         SubCellInst_SboxInst_11_AND1_U1_n7,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_11_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_11_AND3_U1_n9,
         SubCellInst_SboxInst_11_AND3_U1_n8,
         SubCellInst_SboxInst_11_AND3_U1_n7,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_11_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_12_AND1_U1_n9,
         SubCellInst_SboxInst_12_AND1_U1_n8,
         SubCellInst_SboxInst_12_AND1_U1_n7,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_12_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_12_AND3_U1_n9,
         SubCellInst_SboxInst_12_AND3_U1_n8,
         SubCellInst_SboxInst_12_AND3_U1_n7,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_12_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_13_AND1_U1_n9,
         SubCellInst_SboxInst_13_AND1_U1_n8,
         SubCellInst_SboxInst_13_AND1_U1_n7,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_13_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_13_AND3_U1_n9,
         SubCellInst_SboxInst_13_AND3_U1_n8,
         SubCellInst_SboxInst_13_AND3_U1_n7,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_13_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_14_AND1_U1_n9,
         SubCellInst_SboxInst_14_AND1_U1_n8,
         SubCellInst_SboxInst_14_AND1_U1_n7,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_14_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_14_AND3_U1_n9,
         SubCellInst_SboxInst_14_AND3_U1_n8,
         SubCellInst_SboxInst_14_AND3_U1_n7,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_14_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_15_AND1_U1_n9,
         SubCellInst_SboxInst_15_AND1_U1_n8,
         SubCellInst_SboxInst_15_AND1_U1_n7,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_15_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_15_AND3_U1_n9,
         SubCellInst_SboxInst_15_AND3_U1_n8,
         SubCellInst_SboxInst_15_AND3_U1_n7,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_15_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_0_AND2_U1_n9, SubCellInst_SboxInst_0_AND2_U1_n8,
         SubCellInst_SboxInst_0_AND2_U1_n7,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_0_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_0_AND4_U1_n9, SubCellInst_SboxInst_0_AND4_U1_n8,
         SubCellInst_SboxInst_0_AND4_U1_n7,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_0_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_1_AND2_U1_n9, SubCellInst_SboxInst_1_AND2_U1_n8,
         SubCellInst_SboxInst_1_AND2_U1_n7,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_1_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_1_AND4_U1_n9, SubCellInst_SboxInst_1_AND4_U1_n8,
         SubCellInst_SboxInst_1_AND4_U1_n7,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_1_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_2_AND2_U1_n9, SubCellInst_SboxInst_2_AND2_U1_n8,
         SubCellInst_SboxInst_2_AND2_U1_n7,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_2_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_2_AND4_U1_n9, SubCellInst_SboxInst_2_AND4_U1_n8,
         SubCellInst_SboxInst_2_AND4_U1_n7,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_2_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_3_AND2_U1_n9, SubCellInst_SboxInst_3_AND2_U1_n8,
         SubCellInst_SboxInst_3_AND2_U1_n7,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_3_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_3_AND4_U1_n9, SubCellInst_SboxInst_3_AND4_U1_n8,
         SubCellInst_SboxInst_3_AND4_U1_n7,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_3_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_4_AND2_U1_n9, SubCellInst_SboxInst_4_AND2_U1_n8,
         SubCellInst_SboxInst_4_AND2_U1_n7,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_4_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_4_AND4_U1_n9, SubCellInst_SboxInst_4_AND4_U1_n8,
         SubCellInst_SboxInst_4_AND4_U1_n7,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_4_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_5_AND2_U1_n9, SubCellInst_SboxInst_5_AND2_U1_n8,
         SubCellInst_SboxInst_5_AND2_U1_n7,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_5_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_5_AND4_U1_n9, SubCellInst_SboxInst_5_AND4_U1_n8,
         SubCellInst_SboxInst_5_AND4_U1_n7,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_5_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_6_AND2_U1_n9, SubCellInst_SboxInst_6_AND2_U1_n8,
         SubCellInst_SboxInst_6_AND2_U1_n7,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_6_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_6_AND4_U1_n9, SubCellInst_SboxInst_6_AND4_U1_n8,
         SubCellInst_SboxInst_6_AND4_U1_n7,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_6_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_7_AND2_U1_n9, SubCellInst_SboxInst_7_AND2_U1_n8,
         SubCellInst_SboxInst_7_AND2_U1_n7,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_7_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_7_AND4_U1_n9, SubCellInst_SboxInst_7_AND4_U1_n8,
         SubCellInst_SboxInst_7_AND4_U1_n7,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_7_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_8_AND2_U1_n9, SubCellInst_SboxInst_8_AND2_U1_n8,
         SubCellInst_SboxInst_8_AND2_U1_n7,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_8_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_8_AND4_U1_n9, SubCellInst_SboxInst_8_AND4_U1_n8,
         SubCellInst_SboxInst_8_AND4_U1_n7,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_8_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_9_AND2_U1_n9, SubCellInst_SboxInst_9_AND2_U1_n8,
         SubCellInst_SboxInst_9_AND2_U1_n7,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_9_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_9_AND4_U1_n9, SubCellInst_SboxInst_9_AND4_U1_n8,
         SubCellInst_SboxInst_9_AND4_U1_n7,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_9_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_10_AND2_U1_n9,
         SubCellInst_SboxInst_10_AND2_U1_n8,
         SubCellInst_SboxInst_10_AND2_U1_n7,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_10_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_10_AND4_U1_n9,
         SubCellInst_SboxInst_10_AND4_U1_n8,
         SubCellInst_SboxInst_10_AND4_U1_n7,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_10_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_11_AND2_U1_n9,
         SubCellInst_SboxInst_11_AND2_U1_n8,
         SubCellInst_SboxInst_11_AND2_U1_n7,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_11_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_11_AND4_U1_n9,
         SubCellInst_SboxInst_11_AND4_U1_n8,
         SubCellInst_SboxInst_11_AND4_U1_n7,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_11_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_12_AND2_U1_n9,
         SubCellInst_SboxInst_12_AND2_U1_n8,
         SubCellInst_SboxInst_12_AND2_U1_n7,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_12_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_12_AND4_U1_n9,
         SubCellInst_SboxInst_12_AND4_U1_n8,
         SubCellInst_SboxInst_12_AND4_U1_n7,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_12_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_13_AND2_U1_n9,
         SubCellInst_SboxInst_13_AND2_U1_n8,
         SubCellInst_SboxInst_13_AND2_U1_n7,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_13_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_13_AND4_U1_n9,
         SubCellInst_SboxInst_13_AND4_U1_n8,
         SubCellInst_SboxInst_13_AND4_U1_n7,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_13_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_14_AND2_U1_n9,
         SubCellInst_SboxInst_14_AND2_U1_n8,
         SubCellInst_SboxInst_14_AND2_U1_n7,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_14_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_14_AND4_U1_n9,
         SubCellInst_SboxInst_14_AND4_U1_n8,
         SubCellInst_SboxInst_14_AND4_U1_n7,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_14_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_15_AND2_U1_n9,
         SubCellInst_SboxInst_15_AND2_U1_n8,
         SubCellInst_SboxInst_15_AND2_U1_n7,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_15_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_15_AND4_U1_n9,
         SubCellInst_SboxInst_15_AND4_U1_n8,
         SubCellInst_SboxInst_15_AND4_U1_n7,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_15_AND4_U1_z_1__1_;
  wire   [63:0] TweakeyGeneration_StateRegInput;
  wire   [63:0] TweakeyGeneration_key_Feedback;
  wire   [4:1] FSMUpdate;
  wire   [5:0] FSMSelected;
  wire   [5:4] FSM;
  wire   [63:0] StateRegInput;
  wire   [63:0] MCOutput;
  wire   [47:0] ShiftRowsOutput;
  wire   [63:32] AddRoundConstantOutput;
  wire   [63:60] SubCellOutput;
  wire   [1:0] SubCellInst_SboxInst_0_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_0_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_0_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_0_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_0_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_0_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_1_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_1_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_1_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_1_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_1_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_1_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_2_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_2_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_2_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_2_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_2_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_2_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_3_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_3_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_3_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_3_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_3_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_3_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_4_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_4_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_4_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_4_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_4_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_4_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_5_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_5_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_5_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_5_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_5_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_5_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_6_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_6_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_6_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_6_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_6_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_6_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_7_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_7_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_7_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_7_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_7_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_7_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_8_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_8_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_8_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_8_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_8_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_8_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_9_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_9_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_9_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_9_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_9_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_9_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_10_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_10_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_10_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_10_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_10_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_10_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_11_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_11_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_11_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_11_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_11_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_11_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_12_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_12_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_12_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_12_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_12_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_12_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_13_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_13_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_13_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_13_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_13_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_13_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_14_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_14_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_14_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_14_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_14_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_14_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_15_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_15_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_15_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_15_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_15_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_15_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_0_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_0_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_0_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_0_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_0_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_0_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_1_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_1_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_1_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_1_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_1_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_1_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_2_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_2_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_2_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_2_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_2_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_2_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_3_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_3_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_3_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_3_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_3_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_3_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_4_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_4_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_4_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_4_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_4_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_4_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_5_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_5_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_5_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_5_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_5_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_5_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_6_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_6_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_6_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_6_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_6_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_6_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_7_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_7_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_7_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_7_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_7_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_7_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_8_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_8_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_8_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_8_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_8_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_8_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_9_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_9_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_9_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_9_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_9_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_9_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_10_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_10_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_10_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_10_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_10_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_10_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_11_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_11_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_11_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_11_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_11_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_11_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_12_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_12_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_12_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_12_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_12_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_12_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_13_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_13_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_13_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_13_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_13_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_13_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_14_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_14_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_14_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_14_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_14_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_14_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_15_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_15_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_15_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_15_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_15_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_15_AND4_U1_mul;

  DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .D(new_AGEMA_signal_4072), .CK(
        clk), .Q(FSM[5]), .QN(n13) );
  DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .D(new_AGEMA_signal_4076), .CK(
        clk), .Q(FSM[4]), .QN(n14) );
  DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .D(new_AGEMA_signal_4080), .CK(
        clk), .Q(FSMUpdate[4]), .QN(n16) );
  DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .D(new_AGEMA_signal_4084), .CK(
        clk), .Q(FSMUpdate[3]), .QN(n17) );
  DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .D(new_AGEMA_signal_4088), .CK(
        clk), .Q(FSM_1), .QN(n15) );
  DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .D(new_AGEMA_signal_4092), .CK(
        clk), .Q(FSMUpdate[1]), .QN(n18) );
  BUF_X1 U39 ( .A(new_AGEMA_signal_2644), .Z(n35) );
  BUF_X1 U40 ( .A(new_AGEMA_signal_2644), .Z(n36) );
  BUF_X1 U41 ( .A(new_AGEMA_signal_2190), .Z(n38) );
  BUF_X1 U42 ( .A(new_AGEMA_signal_2190), .Z(n39) );
  BUF_X1 U43 ( .A(new_AGEMA_signal_2190), .Z(n37) );
  BUF_X1 U44 ( .A(new_AGEMA_signal_2644), .Z(n34) );
  INV_X1 U45 ( .A(rst), .ZN(n40) );
  NAND3_X1 U46 ( .A1(n16), .A2(n17), .A3(FSM_1), .ZN(n46) );
  NOR2_X1 U47 ( .A1(n18), .A2(n46), .ZN(n41) );
  OAI21_X1 U48 ( .B1(n13), .B2(n41), .A(n14), .ZN(n42) );
  OAI211_X1 U49 ( .C1(n13), .C2(n14), .A(n40), .B(n42), .ZN(FSMSelected[0]) );
  NOR2_X1 U50 ( .A1(rst), .A2(n18), .ZN(FSMSelected[1]) );
  NOR2_X1 U51 ( .A1(rst), .A2(n16), .ZN(FSMSelected[4]) );
  NOR2_X1 U52 ( .A1(rst), .A2(n17), .ZN(FSMSelected[3]) );
  NOR2_X1 U53 ( .A1(FSMSelected[4]), .A2(FSMSelected[3]), .ZN(n45) );
  NAND2_X1 U54 ( .A1(n14), .A2(FSM[5]), .ZN(n43) );
  OAI21_X1 U55 ( .B1(n18), .B2(n43), .A(n40), .ZN(n44) );
  AOI21_X1 U56 ( .B1(n45), .B2(n44), .A(n15), .ZN(FSMSelected[2]) );
  NAND2_X1 U57 ( .A1(FSMSelected[1]), .A2(FSM[5]), .ZN(n47) );
  OAI22_X1 U58 ( .A1(rst), .A2(n14), .B1(n47), .B2(n46), .ZN(FSMSelected[5])
         );
  NAND4_X1 U59 ( .A1(n15), .A2(n16), .A3(n17), .A4(FSM[5]), .ZN(n48) );
  NOR3_X1 U60 ( .A1(n14), .A2(n18), .A3(n48), .ZN(done) );
  INV_X1 SubCellInst_SboxInst_0_U1_U1 ( .A(Ciphertext_s0[2]), .ZN(
        SubCellInst_SboxInst_0_n3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[2]), 
        .B(Ciphertext_s0[3]), .Z(SubCellInst_SboxInst_0_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[2]), 
        .B(Ciphertext_s1[3]), .Z(new_AGEMA_signal_1167) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[0]), 
        .B(Ciphertext_s0[2]), .Z(SubCellInst_SboxInst_0_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[0]), 
        .B(Ciphertext_s1[2]), .Z(new_AGEMA_signal_1169) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_XX_2_), .Z(SubCellInst_SboxInst_0_Q0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        new_AGEMA_signal_1169), .Z(new_AGEMA_signal_1453) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_XX_1_), .Z(SubCellInst_SboxInst_0_Q1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        new_AGEMA_signal_1167), .Z(new_AGEMA_signal_1454) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_n3), .ZN(SubCellInst_SboxInst_0_Q4) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        Ciphertext_s1[2]), .Z(new_AGEMA_signal_1455) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_XX_2_), .B(SubCellInst_SboxInst_0_n3), .Z(
        SubCellInst_SboxInst_0_Q6) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1169), 
        .B(Ciphertext_s1[2]), .Z(new_AGEMA_signal_1456) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_0_Q1), .B(SubCellInst_SboxInst_0_Q6), .ZN(
        SubCellInst_SboxInst_0_L1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1454), 
        .B(new_AGEMA_signal_1456), .Z(new_AGEMA_signal_1550) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_n3), .Z(SubCellInst_SboxInst_0_L2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        Ciphertext_s1[2]), .Z(new_AGEMA_signal_1457) );
  INV_X1 SubCellInst_SboxInst_1_U1_U1 ( .A(Ciphertext_s0[6]), .ZN(
        SubCellInst_SboxInst_1_n3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[6]), 
        .B(Ciphertext_s0[7]), .Z(SubCellInst_SboxInst_1_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[6]), 
        .B(Ciphertext_s1[7]), .Z(new_AGEMA_signal_1173) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[4]), 
        .B(Ciphertext_s0[6]), .Z(SubCellInst_SboxInst_1_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[4]), 
        .B(Ciphertext_s1[6]), .Z(new_AGEMA_signal_1175) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_XX_2_), .Z(SubCellInst_SboxInst_1_Q0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        new_AGEMA_signal_1175), .Z(new_AGEMA_signal_1459) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_XX_1_), .Z(SubCellInst_SboxInst_1_Q1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        new_AGEMA_signal_1173), .Z(new_AGEMA_signal_1460) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_n3), .ZN(SubCellInst_SboxInst_1_Q4) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        Ciphertext_s1[6]), .Z(new_AGEMA_signal_1461) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_XX_2_), .B(SubCellInst_SboxInst_1_n3), .Z(
        SubCellInst_SboxInst_1_Q6) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1175), 
        .B(Ciphertext_s1[6]), .Z(new_AGEMA_signal_1462) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_1_Q1), .B(SubCellInst_SboxInst_1_Q6), .ZN(
        SubCellInst_SboxInst_1_L1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1460), 
        .B(new_AGEMA_signal_1462), .Z(new_AGEMA_signal_1553) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_n3), .Z(SubCellInst_SboxInst_1_L2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        Ciphertext_s1[6]), .Z(new_AGEMA_signal_1463) );
  INV_X1 SubCellInst_SboxInst_2_U1_U1 ( .A(Ciphertext_s0[10]), .ZN(
        SubCellInst_SboxInst_2_n3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[10]), 
        .B(Ciphertext_s0[11]), .Z(SubCellInst_SboxInst_2_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[10]), 
        .B(Ciphertext_s1[11]), .Z(new_AGEMA_signal_1179) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[8]), 
        .B(Ciphertext_s0[10]), .Z(SubCellInst_SboxInst_2_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[8]), 
        .B(Ciphertext_s1[10]), .Z(new_AGEMA_signal_1181) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_XX_2_), .Z(SubCellInst_SboxInst_2_Q0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        new_AGEMA_signal_1181), .Z(new_AGEMA_signal_1465) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_XX_1_), .Z(SubCellInst_SboxInst_2_Q1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        new_AGEMA_signal_1179), .Z(new_AGEMA_signal_1466) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_n3), .ZN(SubCellInst_SboxInst_2_Q4) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        Ciphertext_s1[10]), .Z(new_AGEMA_signal_1467) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_XX_2_), .B(SubCellInst_SboxInst_2_n3), .Z(
        SubCellInst_SboxInst_2_Q6) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1181), 
        .B(Ciphertext_s1[10]), .Z(new_AGEMA_signal_1468) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_2_Q1), .B(SubCellInst_SboxInst_2_Q6), .ZN(
        SubCellInst_SboxInst_2_L1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1466), 
        .B(new_AGEMA_signal_1468), .Z(new_AGEMA_signal_1556) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_n3), .Z(SubCellInst_SboxInst_2_L2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        Ciphertext_s1[10]), .Z(new_AGEMA_signal_1469) );
  INV_X1 SubCellInst_SboxInst_3_U1_U1 ( .A(Ciphertext_s0[14]), .ZN(
        SubCellInst_SboxInst_3_n3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[14]), 
        .B(Ciphertext_s0[15]), .Z(SubCellInst_SboxInst_3_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[14]), 
        .B(Ciphertext_s1[15]), .Z(new_AGEMA_signal_1185) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[12]), 
        .B(Ciphertext_s0[14]), .Z(SubCellInst_SboxInst_3_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[12]), 
        .B(Ciphertext_s1[14]), .Z(new_AGEMA_signal_1187) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_XX_2_), .Z(SubCellInst_SboxInst_3_Q0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        new_AGEMA_signal_1187), .Z(new_AGEMA_signal_1471) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_XX_1_), .Z(SubCellInst_SboxInst_3_Q1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        new_AGEMA_signal_1185), .Z(new_AGEMA_signal_1472) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_n3), .ZN(SubCellInst_SboxInst_3_Q4) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        Ciphertext_s1[14]), .Z(new_AGEMA_signal_1473) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_XX_2_), .B(SubCellInst_SboxInst_3_n3), .Z(
        SubCellInst_SboxInst_3_Q6) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1187), 
        .B(Ciphertext_s1[14]), .Z(new_AGEMA_signal_1474) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_3_Q1), .B(SubCellInst_SboxInst_3_Q6), .ZN(
        SubCellInst_SboxInst_3_L1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1472), 
        .B(new_AGEMA_signal_1474), .Z(new_AGEMA_signal_1559) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_n3), .Z(SubCellInst_SboxInst_3_L2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        Ciphertext_s1[14]), .Z(new_AGEMA_signal_1475) );
  INV_X1 SubCellInst_SboxInst_4_U1_U1 ( .A(Ciphertext_s0[18]), .ZN(
        SubCellInst_SboxInst_4_n3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[18]), 
        .B(Ciphertext_s0[19]), .Z(SubCellInst_SboxInst_4_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[18]), 
        .B(Ciphertext_s1[19]), .Z(new_AGEMA_signal_1191) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[16]), 
        .B(Ciphertext_s0[18]), .Z(SubCellInst_SboxInst_4_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[16]), 
        .B(Ciphertext_s1[18]), .Z(new_AGEMA_signal_1193) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_XX_2_), .Z(SubCellInst_SboxInst_4_Q0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        new_AGEMA_signal_1193), .Z(new_AGEMA_signal_1477) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_XX_1_), .Z(SubCellInst_SboxInst_4_Q1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        new_AGEMA_signal_1191), .Z(new_AGEMA_signal_1478) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_n3), .ZN(SubCellInst_SboxInst_4_Q4) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        Ciphertext_s1[18]), .Z(new_AGEMA_signal_1479) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_XX_2_), .B(SubCellInst_SboxInst_4_n3), .Z(
        SubCellInst_SboxInst_4_Q6) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1193), 
        .B(Ciphertext_s1[18]), .Z(new_AGEMA_signal_1480) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_4_Q1), .B(SubCellInst_SboxInst_4_Q6), .ZN(
        SubCellInst_SboxInst_4_L1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1478), 
        .B(new_AGEMA_signal_1480), .Z(new_AGEMA_signal_1562) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_n3), .Z(SubCellInst_SboxInst_4_L2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        Ciphertext_s1[18]), .Z(new_AGEMA_signal_1481) );
  INV_X1 SubCellInst_SboxInst_5_U1_U1 ( .A(Ciphertext_s0[22]), .ZN(
        SubCellInst_SboxInst_5_n3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[22]), 
        .B(Ciphertext_s0[23]), .Z(SubCellInst_SboxInst_5_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[22]), 
        .B(Ciphertext_s1[23]), .Z(new_AGEMA_signal_1197) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[20]), 
        .B(Ciphertext_s0[22]), .Z(SubCellInst_SboxInst_5_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[20]), 
        .B(Ciphertext_s1[22]), .Z(new_AGEMA_signal_1199) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_XX_2_), .Z(SubCellInst_SboxInst_5_Q0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        new_AGEMA_signal_1199), .Z(new_AGEMA_signal_1483) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_XX_1_), .Z(SubCellInst_SboxInst_5_Q1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        new_AGEMA_signal_1197), .Z(new_AGEMA_signal_1484) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_n3), .ZN(SubCellInst_SboxInst_5_Q4) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        Ciphertext_s1[22]), .Z(new_AGEMA_signal_1485) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_XX_2_), .B(SubCellInst_SboxInst_5_n3), .Z(
        SubCellInst_SboxInst_5_Q6) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1199), 
        .B(Ciphertext_s1[22]), .Z(new_AGEMA_signal_1486) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_5_Q1), .B(SubCellInst_SboxInst_5_Q6), .ZN(
        SubCellInst_SboxInst_5_L1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1484), 
        .B(new_AGEMA_signal_1486), .Z(new_AGEMA_signal_1565) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_n3), .Z(SubCellInst_SboxInst_5_L2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        Ciphertext_s1[22]), .Z(new_AGEMA_signal_1487) );
  INV_X1 SubCellInst_SboxInst_6_U1_U1 ( .A(Ciphertext_s0[26]), .ZN(
        SubCellInst_SboxInst_6_n3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[26]), 
        .B(Ciphertext_s0[27]), .Z(SubCellInst_SboxInst_6_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[26]), 
        .B(Ciphertext_s1[27]), .Z(new_AGEMA_signal_1203) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[24]), 
        .B(Ciphertext_s0[26]), .Z(SubCellInst_SboxInst_6_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[24]), 
        .B(Ciphertext_s1[26]), .Z(new_AGEMA_signal_1205) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_XX_2_), .Z(SubCellInst_SboxInst_6_Q0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        new_AGEMA_signal_1205), .Z(new_AGEMA_signal_1489) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_XX_1_), .Z(SubCellInst_SboxInst_6_Q1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        new_AGEMA_signal_1203), .Z(new_AGEMA_signal_1490) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_n3), .ZN(SubCellInst_SboxInst_6_Q4) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        Ciphertext_s1[26]), .Z(new_AGEMA_signal_1491) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_XX_2_), .B(SubCellInst_SboxInst_6_n3), .Z(
        SubCellInst_SboxInst_6_Q6) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1205), 
        .B(Ciphertext_s1[26]), .Z(new_AGEMA_signal_1492) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_6_Q1), .B(SubCellInst_SboxInst_6_Q6), .ZN(
        SubCellInst_SboxInst_6_L1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1490), 
        .B(new_AGEMA_signal_1492), .Z(new_AGEMA_signal_1568) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_n3), .Z(SubCellInst_SboxInst_6_L2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        Ciphertext_s1[26]), .Z(new_AGEMA_signal_1493) );
  INV_X1 SubCellInst_SboxInst_7_U1_U1 ( .A(Ciphertext_s0[30]), .ZN(
        SubCellInst_SboxInst_7_n3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[30]), 
        .B(Ciphertext_s0[31]), .Z(SubCellInst_SboxInst_7_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[30]), 
        .B(Ciphertext_s1[31]), .Z(new_AGEMA_signal_1209) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[28]), 
        .B(Ciphertext_s0[30]), .Z(SubCellInst_SboxInst_7_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[28]), 
        .B(Ciphertext_s1[30]), .Z(new_AGEMA_signal_1211) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_XX_2_), .Z(SubCellInst_SboxInst_7_Q0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        new_AGEMA_signal_1211), .Z(new_AGEMA_signal_1495) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_XX_1_), .Z(SubCellInst_SboxInst_7_Q1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        new_AGEMA_signal_1209), .Z(new_AGEMA_signal_1496) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_n3), .ZN(SubCellInst_SboxInst_7_Q4) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        Ciphertext_s1[30]), .Z(new_AGEMA_signal_1497) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_XX_2_), .B(SubCellInst_SboxInst_7_n3), .Z(
        SubCellInst_SboxInst_7_Q6) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1211), 
        .B(Ciphertext_s1[30]), .Z(new_AGEMA_signal_1498) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_7_Q1), .B(SubCellInst_SboxInst_7_Q6), .ZN(
        SubCellInst_SboxInst_7_L1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1496), 
        .B(new_AGEMA_signal_1498), .Z(new_AGEMA_signal_1571) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_n3), .Z(SubCellInst_SboxInst_7_L2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        Ciphertext_s1[30]), .Z(new_AGEMA_signal_1499) );
  INV_X1 SubCellInst_SboxInst_8_U1_U1 ( .A(Ciphertext_s0[34]), .ZN(
        SubCellInst_SboxInst_8_n3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[34]), 
        .B(Ciphertext_s0[35]), .Z(SubCellInst_SboxInst_8_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[34]), 
        .B(Ciphertext_s1[35]), .Z(new_AGEMA_signal_1215) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[32]), 
        .B(Ciphertext_s0[34]), .Z(SubCellInst_SboxInst_8_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[32]), 
        .B(Ciphertext_s1[34]), .Z(new_AGEMA_signal_1217) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_XX_2_), .Z(SubCellInst_SboxInst_8_Q0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        new_AGEMA_signal_1217), .Z(new_AGEMA_signal_1501) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_XX_1_), .Z(SubCellInst_SboxInst_8_Q1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        new_AGEMA_signal_1215), .Z(new_AGEMA_signal_1502) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_n3), .ZN(SubCellInst_SboxInst_8_Q4) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        Ciphertext_s1[34]), .Z(new_AGEMA_signal_1503) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_XX_2_), .B(SubCellInst_SboxInst_8_n3), .Z(
        SubCellInst_SboxInst_8_Q6) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1217), 
        .B(Ciphertext_s1[34]), .Z(new_AGEMA_signal_1504) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_8_Q1), .B(SubCellInst_SboxInst_8_Q6), .ZN(
        SubCellInst_SboxInst_8_L1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1502), 
        .B(new_AGEMA_signal_1504), .Z(new_AGEMA_signal_1574) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_n3), .Z(SubCellInst_SboxInst_8_L2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        Ciphertext_s1[34]), .Z(new_AGEMA_signal_1505) );
  INV_X1 SubCellInst_SboxInst_9_U1_U1 ( .A(Ciphertext_s0[38]), .ZN(
        SubCellInst_SboxInst_9_n3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[38]), 
        .B(Ciphertext_s0[39]), .Z(SubCellInst_SboxInst_9_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[38]), 
        .B(Ciphertext_s1[39]), .Z(new_AGEMA_signal_1221) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[36]), 
        .B(Ciphertext_s0[38]), .Z(SubCellInst_SboxInst_9_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[36]), 
        .B(Ciphertext_s1[38]), .Z(new_AGEMA_signal_1223) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_XX_2_), .Z(SubCellInst_SboxInst_9_Q0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        new_AGEMA_signal_1223), .Z(new_AGEMA_signal_1507) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_XX_1_), .Z(SubCellInst_SboxInst_9_Q1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        new_AGEMA_signal_1221), .Z(new_AGEMA_signal_1508) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_n3), .ZN(SubCellInst_SboxInst_9_Q4) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        Ciphertext_s1[38]), .Z(new_AGEMA_signal_1509) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_XX_2_), .B(SubCellInst_SboxInst_9_n3), .Z(
        SubCellInst_SboxInst_9_Q6) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1223), 
        .B(Ciphertext_s1[38]), .Z(new_AGEMA_signal_1510) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_9_Q1), .B(SubCellInst_SboxInst_9_Q6), .ZN(
        SubCellInst_SboxInst_9_L1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1508), 
        .B(new_AGEMA_signal_1510), .Z(new_AGEMA_signal_1577) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_n3), .Z(SubCellInst_SboxInst_9_L2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        Ciphertext_s1[38]), .Z(new_AGEMA_signal_1511) );
  INV_X1 SubCellInst_SboxInst_10_U1_U1 ( .A(Ciphertext_s0[42]), .ZN(
        SubCellInst_SboxInst_10_n3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[42]), 
        .B(Ciphertext_s0[43]), .Z(SubCellInst_SboxInst_10_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[42]), 
        .B(Ciphertext_s1[43]), .Z(new_AGEMA_signal_1227) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[40]), 
        .B(Ciphertext_s0[42]), .Z(SubCellInst_SboxInst_10_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[40]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1229) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_XX_2_), .Z(SubCellInst_SboxInst_10_Q0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(new_AGEMA_signal_1229), .Z(new_AGEMA_signal_1513) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_XX_1_), .Z(SubCellInst_SboxInst_10_Q1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(new_AGEMA_signal_1227), .Z(new_AGEMA_signal_1514) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_Q4) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1515) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_XX_2_), .B(SubCellInst_SboxInst_10_n3), .Z(
        SubCellInst_SboxInst_10_Q6) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1229), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1516) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_10_Q1), .B(SubCellInst_SboxInst_10_Q6), .ZN(
        SubCellInst_SboxInst_10_L1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1514), 
        .B(new_AGEMA_signal_1516), .Z(new_AGEMA_signal_1580) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_n3), .Z(SubCellInst_SboxInst_10_L2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1517) );
  INV_X1 SubCellInst_SboxInst_11_U1_U1 ( .A(Ciphertext_s0[46]), .ZN(
        SubCellInst_SboxInst_11_n3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[46]), 
        .B(Ciphertext_s0[47]), .Z(SubCellInst_SboxInst_11_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[46]), 
        .B(Ciphertext_s1[47]), .Z(new_AGEMA_signal_1233) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[44]), 
        .B(Ciphertext_s0[46]), .Z(SubCellInst_SboxInst_11_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[44]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1235) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_XX_2_), .Z(SubCellInst_SboxInst_11_Q0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(new_AGEMA_signal_1235), .Z(new_AGEMA_signal_1519) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_XX_1_), .Z(SubCellInst_SboxInst_11_Q1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(new_AGEMA_signal_1233), .Z(new_AGEMA_signal_1520) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_Q4) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1521) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_XX_2_), .B(SubCellInst_SboxInst_11_n3), .Z(
        SubCellInst_SboxInst_11_Q6) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1235), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1522) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_11_Q1), .B(SubCellInst_SboxInst_11_Q6), .ZN(
        SubCellInst_SboxInst_11_L1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1520), 
        .B(new_AGEMA_signal_1522), .Z(new_AGEMA_signal_1583) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_n3), .Z(SubCellInst_SboxInst_11_L2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1523) );
  INV_X1 SubCellInst_SboxInst_12_U1_U1 ( .A(Ciphertext_s0[50]), .ZN(
        SubCellInst_SboxInst_12_n3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[50]), 
        .B(Ciphertext_s0[51]), .Z(SubCellInst_SboxInst_12_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[50]), 
        .B(Ciphertext_s1[51]), .Z(new_AGEMA_signal_1239) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[48]), 
        .B(Ciphertext_s0[50]), .Z(SubCellInst_SboxInst_12_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[48]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1241) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_XX_2_), .Z(SubCellInst_SboxInst_12_Q0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(new_AGEMA_signal_1241), .Z(new_AGEMA_signal_1525) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_XX_1_), .Z(SubCellInst_SboxInst_12_Q1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(new_AGEMA_signal_1239), .Z(new_AGEMA_signal_1526) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_Q4) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1527) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_XX_2_), .B(SubCellInst_SboxInst_12_n3), .Z(
        SubCellInst_SboxInst_12_Q6) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1241), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1528) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_12_Q1), .B(SubCellInst_SboxInst_12_Q6), .ZN(
        SubCellInst_SboxInst_12_L1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1526), 
        .B(new_AGEMA_signal_1528), .Z(new_AGEMA_signal_1586) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_n3), .Z(SubCellInst_SboxInst_12_L2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1529) );
  INV_X1 SubCellInst_SboxInst_13_U1_U1 ( .A(Ciphertext_s0[54]), .ZN(
        SubCellInst_SboxInst_13_n3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[54]), 
        .B(Ciphertext_s0[55]), .Z(SubCellInst_SboxInst_13_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[54]), 
        .B(Ciphertext_s1[55]), .Z(new_AGEMA_signal_1245) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[52]), 
        .B(Ciphertext_s0[54]), .Z(SubCellInst_SboxInst_13_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[52]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1247) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_XX_2_), .Z(SubCellInst_SboxInst_13_Q0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(new_AGEMA_signal_1247), .Z(new_AGEMA_signal_1531) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_XX_1_), .Z(SubCellInst_SboxInst_13_Q1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(new_AGEMA_signal_1245), .Z(new_AGEMA_signal_1532) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_Q4) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1533) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_XX_2_), .B(SubCellInst_SboxInst_13_n3), .Z(
        SubCellInst_SboxInst_13_Q6) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1247), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1534) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_13_Q1), .B(SubCellInst_SboxInst_13_Q6), .ZN(
        SubCellInst_SboxInst_13_L1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1532), 
        .B(new_AGEMA_signal_1534), .Z(new_AGEMA_signal_1589) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_n3), .Z(SubCellInst_SboxInst_13_L2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1535) );
  INV_X1 SubCellInst_SboxInst_14_U1_U1 ( .A(Ciphertext_s0[58]), .ZN(
        SubCellInst_SboxInst_14_n3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[58]), 
        .B(Ciphertext_s0[59]), .Z(SubCellInst_SboxInst_14_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[58]), 
        .B(Ciphertext_s1[59]), .Z(new_AGEMA_signal_1251) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[56]), 
        .B(Ciphertext_s0[58]), .Z(SubCellInst_SboxInst_14_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[56]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1253) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_XX_2_), .Z(SubCellInst_SboxInst_14_Q0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(new_AGEMA_signal_1253), .Z(new_AGEMA_signal_1537) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_XX_1_), .Z(SubCellInst_SboxInst_14_Q1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(new_AGEMA_signal_1251), .Z(new_AGEMA_signal_1538) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_Q4) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1539) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_XX_2_), .B(SubCellInst_SboxInst_14_n3), .Z(
        SubCellInst_SboxInst_14_Q6) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1253), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1540) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_14_Q1), .B(SubCellInst_SboxInst_14_Q6), .ZN(
        SubCellInst_SboxInst_14_L1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1538), 
        .B(new_AGEMA_signal_1540), .Z(new_AGEMA_signal_1592) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_n3), .Z(SubCellInst_SboxInst_14_L2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1541) );
  INV_X1 SubCellInst_SboxInst_15_U1_U1 ( .A(Ciphertext_s0[62]), .ZN(
        SubCellInst_SboxInst_15_n3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[62]), 
        .B(Ciphertext_s0[63]), .Z(SubCellInst_SboxInst_15_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[62]), 
        .B(Ciphertext_s1[63]), .Z(new_AGEMA_signal_1257) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[60]), 
        .B(Ciphertext_s0[62]), .Z(SubCellInst_SboxInst_15_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[60]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1259) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_XX_2_), .Z(SubCellInst_SboxInst_15_Q0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(new_AGEMA_signal_1259), .Z(new_AGEMA_signal_1543) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_XX_1_), .Z(SubCellInst_SboxInst_15_Q1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(new_AGEMA_signal_1257), .Z(new_AGEMA_signal_1544) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_Q4) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1545) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_XX_2_), .B(SubCellInst_SboxInst_15_n3), .Z(
        SubCellInst_SboxInst_15_Q6) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1259), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1546) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_15_Q1), .B(SubCellInst_SboxInst_15_Q6), .ZN(
        SubCellInst_SboxInst_15_L1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1544), 
        .B(new_AGEMA_signal_1546), .Z(new_AGEMA_signal_1595) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_n3), .Z(SubCellInst_SboxInst_15_L2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1547) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[0]), .B(Key_s0[0]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[0]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1260), .B(Key_s1[0]), .S(rst), .Z(
        new_AGEMA_signal_1262) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[1]), .B(Key_s0[1]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[1]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1263), .B(Key_s1[1]), .S(rst), .Z(
        new_AGEMA_signal_1265) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[2]), .B(Key_s0[2]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[2]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1266), .B(Key_s1[2]), .S(rst), .Z(
        new_AGEMA_signal_1268) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[3]), .B(Key_s0[3]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[3]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1269), .B(Key_s1[3]), .S(rst), .Z(
        new_AGEMA_signal_1271) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[4]), .B(Key_s0[4]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[4]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1272), .B(Key_s1[4]), .S(rst), .Z(
        new_AGEMA_signal_1274) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[5]), .B(Key_s0[5]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[5]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1275), .B(Key_s1[5]), .S(rst), .Z(
        new_AGEMA_signal_1277) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[6]), .B(Key_s0[6]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[6]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1278), .B(Key_s1[6]), .S(rst), .Z(
        new_AGEMA_signal_1280) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[7]), .B(Key_s0[7]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[7]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1281), .B(Key_s1[7]), .S(rst), .Z(
        new_AGEMA_signal_1283) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[8]), .B(Key_s0[8]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[8]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1284), .B(Key_s1[8]), .S(rst), .Z(
        new_AGEMA_signal_1286) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[9]), .B(Key_s0[9]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[9]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1287), .B(Key_s1[9]), .S(rst), .Z(
        new_AGEMA_signal_1289) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[10]), .B(Key_s0[10]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[10]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1290), .B(Key_s1[10]), .S(rst), .Z(
        new_AGEMA_signal_1292) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[11]), .B(Key_s0[11]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[11]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1293), .B(Key_s1[11]), .S(rst), .Z(
        new_AGEMA_signal_1295) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[12]), .B(Key_s0[12]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[12]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1296), .B(Key_s1[12]), .S(rst), .Z(
        new_AGEMA_signal_1298) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[13]), .B(Key_s0[13]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[13]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1299), .B(Key_s1[13]), .S(rst), .Z(
        new_AGEMA_signal_1301) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[14]), .B(Key_s0[14]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[14]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1302), .B(Key_s1[14]), .S(rst), .Z(
        new_AGEMA_signal_1304) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[15]), .B(Key_s0[15]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[15]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1305), .B(Key_s1[15]), .S(rst), .Z(
        new_AGEMA_signal_1307) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[16]), .B(Key_s0[16]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[16]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1308), .B(Key_s1[16]), .S(rst), .Z(
        new_AGEMA_signal_1310) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[17]), .B(Key_s0[17]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[17]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1311), .B(Key_s1[17]), .S(rst), .Z(
        new_AGEMA_signal_1313) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[18]), .B(Key_s0[18]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[18]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1314), .B(Key_s1[18]), .S(rst), .Z(
        new_AGEMA_signal_1316) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[19]), .B(Key_s0[19]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[19]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1317), .B(Key_s1[19]), .S(rst), .Z(
        new_AGEMA_signal_1319) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[20]), .B(Key_s0[20]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[20]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1320), .B(Key_s1[20]), .S(rst), .Z(
        new_AGEMA_signal_1322) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[21]), .B(Key_s0[21]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[21]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1323), .B(Key_s1[21]), .S(rst), .Z(
        new_AGEMA_signal_1325) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[22]), .B(Key_s0[22]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[22]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1326), .B(Key_s1[22]), .S(rst), .Z(
        new_AGEMA_signal_1328) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[23]), .B(Key_s0[23]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[23]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1329), .B(Key_s1[23]), .S(rst), .Z(
        new_AGEMA_signal_1331) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[24]), .B(Key_s0[24]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[24]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1332), .B(Key_s1[24]), .S(rst), .Z(
        new_AGEMA_signal_1334) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[25]), .B(Key_s0[25]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[25]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1335), .B(Key_s1[25]), .S(rst), .Z(
        new_AGEMA_signal_1337) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[26]), .B(Key_s0[26]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[26]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1338), .B(Key_s1[26]), .S(rst), .Z(
        new_AGEMA_signal_1340) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[27]), .B(Key_s0[27]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[27]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1341), .B(Key_s1[27]), .S(rst), .Z(
        new_AGEMA_signal_1343) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[28]), .B(Key_s0[28]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[28]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1344), .B(Key_s1[28]), .S(rst), .Z(
        new_AGEMA_signal_1346) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[29]), .B(Key_s0[29]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[29]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1347), .B(Key_s1[29]), .S(rst), .Z(
        new_AGEMA_signal_1349) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[30]), .B(Key_s0[30]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[30]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1350), .B(Key_s1[30]), .S(rst), .Z(
        new_AGEMA_signal_1352) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[31]), .B(Key_s0[31]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[31]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1353), .B(Key_s1[31]), .S(rst), .Z(
        new_AGEMA_signal_1355) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[32]), .B(Key_s0[32]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[32]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1356), .B(Key_s1[32]), .S(rst), .Z(
        new_AGEMA_signal_1358) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[33]), .B(Key_s0[33]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[33]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1359), .B(Key_s1[33]), .S(rst), .Z(
        new_AGEMA_signal_1361) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[34]), .B(Key_s0[34]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[34]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1362), .B(Key_s1[34]), .S(rst), .Z(
        new_AGEMA_signal_1364) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[35]), .B(Key_s0[35]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[35]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1365), .B(Key_s1[35]), .S(rst), .Z(
        new_AGEMA_signal_1367) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[36]), .B(Key_s0[36]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[36]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1368), .B(Key_s1[36]), .S(rst), .Z(
        new_AGEMA_signal_1370) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[37]), .B(Key_s0[37]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[37]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1371), .B(Key_s1[37]), .S(rst), .Z(
        new_AGEMA_signal_1373) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[38]), .B(Key_s0[38]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[38]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1374), .B(Key_s1[38]), .S(rst), .Z(
        new_AGEMA_signal_1376) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[39]), .B(Key_s0[39]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[39]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1377), .B(Key_s1[39]), .S(rst), .Z(
        new_AGEMA_signal_1379) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[40]), .B(Key_s0[40]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[40]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1380), .B(Key_s1[40]), .S(rst), .Z(
        new_AGEMA_signal_1382) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[41]), .B(Key_s0[41]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[41]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1383), .B(Key_s1[41]), .S(rst), .Z(
        new_AGEMA_signal_1385) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[42]), .B(Key_s0[42]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[42]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1386), .B(Key_s1[42]), .S(rst), .Z(
        new_AGEMA_signal_1388) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[43]), .B(Key_s0[43]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[43]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1389), .B(Key_s1[43]), .S(rst), .Z(
        new_AGEMA_signal_1391) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[44]), .B(Key_s0[44]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[44]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1392), .B(Key_s1[44]), .S(rst), .Z(
        new_AGEMA_signal_1394) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[45]), .B(Key_s0[45]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[45]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1395), .B(Key_s1[45]), .S(rst), .Z(
        new_AGEMA_signal_1397) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[46]), .B(Key_s0[46]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[46]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1398), .B(Key_s1[46]), .S(rst), .Z(
        new_AGEMA_signal_1400) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[47]), .B(Key_s0[47]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[47]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1401), .B(Key_s1[47]), .S(rst), .Z(
        new_AGEMA_signal_1403) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[48]), .B(Key_s0[48]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[48]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1404), .B(Key_s1[48]), .S(rst), .Z(
        new_AGEMA_signal_1406) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[49]), .B(Key_s0[49]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[49]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1407), .B(Key_s1[49]), .S(rst), .Z(
        new_AGEMA_signal_1409) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[50]), .B(Key_s0[50]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[50]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1410), .B(Key_s1[50]), .S(rst), .Z(
        new_AGEMA_signal_1412) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[51]), .B(Key_s0[51]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[51]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1413), .B(Key_s1[51]), .S(rst), .Z(
        new_AGEMA_signal_1415) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[52]), .B(Key_s0[52]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[52]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1416), .B(Key_s1[52]), .S(rst), .Z(
        new_AGEMA_signal_1418) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[53]), .B(Key_s0[53]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[53]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1419), .B(Key_s1[53]), .S(rst), .Z(
        new_AGEMA_signal_1421) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[54]), .B(Key_s0[54]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[54]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1422), .B(Key_s1[54]), .S(rst), .Z(
        new_AGEMA_signal_1424) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[55]), .B(Key_s0[55]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[55]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1425), .B(Key_s1[55]), .S(rst), .Z(
        new_AGEMA_signal_1427) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[56]), .B(Key_s0[56]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[56]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1428), .B(Key_s1[56]), .S(rst), .Z(
        new_AGEMA_signal_1430) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[57]), .B(Key_s0[57]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[57]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1431), .B(Key_s1[57]), .S(rst), .Z(
        new_AGEMA_signal_1433) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[58]), .B(Key_s0[58]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[58]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1434), .B(Key_s1[58]), .S(rst), .Z(
        new_AGEMA_signal_1436) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[59]), .B(Key_s0[59]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[59]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1437), .B(Key_s1[59]), .S(rst), .Z(
        new_AGEMA_signal_1439) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[60]), .B(Key_s0[60]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[60]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1440), .B(Key_s1[60]), .S(rst), .Z(
        new_AGEMA_signal_1442) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[61]), .B(Key_s0[61]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[61]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1443), .B(Key_s1[61]), .S(rst), .Z(
        new_AGEMA_signal_1445) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[62]), .B(Key_s0[62]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[62]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1446), .B(Key_s1[62]), .S(rst), .Z(
        new_AGEMA_signal_1448) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[63]), .B(Key_s0[63]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[63]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1449), .B(Key_s1[63]), .S(rst), .Z(
        new_AGEMA_signal_1451) );
  DFF_X1 new_AGEMA_reg_buffer_1000_s_current_state_reg ( .D(rst), .CK(clk), 
        .Q(new_AGEMA_signal_2189), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1002_s_current_state_reg ( .D(Plaintext_s0[2]), 
        .CK(clk), .Q(new_AGEMA_signal_2191), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1004_s_current_state_reg ( .D(Plaintext_s1[2]), 
        .CK(clk), .Q(new_AGEMA_signal_2193), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1006_s_current_state_reg ( .D(Plaintext_s0[3]), 
        .CK(clk), .Q(new_AGEMA_signal_2195), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1008_s_current_state_reg ( .D(Plaintext_s1[3]), 
        .CK(clk), .Q(new_AGEMA_signal_2197), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1010_s_current_state_reg ( .D(Plaintext_s0[6]), 
        .CK(clk), .Q(new_AGEMA_signal_2199), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1012_s_current_state_reg ( .D(Plaintext_s1[6]), 
        .CK(clk), .Q(new_AGEMA_signal_2201), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1014_s_current_state_reg ( .D(Plaintext_s0[7]), 
        .CK(clk), .Q(new_AGEMA_signal_2203), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1016_s_current_state_reg ( .D(Plaintext_s1[7]), 
        .CK(clk), .Q(new_AGEMA_signal_2205), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1018_s_current_state_reg ( .D(Plaintext_s0[10]), 
        .CK(clk), .Q(new_AGEMA_signal_2207), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1020_s_current_state_reg ( .D(Plaintext_s1[10]), 
        .CK(clk), .Q(new_AGEMA_signal_2209), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1022_s_current_state_reg ( .D(Plaintext_s0[11]), 
        .CK(clk), .Q(new_AGEMA_signal_2211), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1024_s_current_state_reg ( .D(Plaintext_s1[11]), 
        .CK(clk), .Q(new_AGEMA_signal_2213), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1026_s_current_state_reg ( .D(Plaintext_s0[14]), 
        .CK(clk), .Q(new_AGEMA_signal_2215), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1028_s_current_state_reg ( .D(Plaintext_s1[14]), 
        .CK(clk), .Q(new_AGEMA_signal_2217), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1030_s_current_state_reg ( .D(Plaintext_s0[15]), 
        .CK(clk), .Q(new_AGEMA_signal_2219), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1032_s_current_state_reg ( .D(Plaintext_s1[15]), 
        .CK(clk), .Q(new_AGEMA_signal_2221), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1034_s_current_state_reg ( .D(Plaintext_s0[18]), 
        .CK(clk), .Q(new_AGEMA_signal_2223), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1036_s_current_state_reg ( .D(Plaintext_s1[18]), 
        .CK(clk), .Q(new_AGEMA_signal_2225), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1038_s_current_state_reg ( .D(Plaintext_s0[19]), 
        .CK(clk), .Q(new_AGEMA_signal_2227), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1040_s_current_state_reg ( .D(Plaintext_s1[19]), 
        .CK(clk), .Q(new_AGEMA_signal_2229), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1042_s_current_state_reg ( .D(Plaintext_s0[22]), 
        .CK(clk), .Q(new_AGEMA_signal_2231), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1044_s_current_state_reg ( .D(Plaintext_s1[22]), 
        .CK(clk), .Q(new_AGEMA_signal_2233), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1046_s_current_state_reg ( .D(Plaintext_s0[23]), 
        .CK(clk), .Q(new_AGEMA_signal_2235), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1048_s_current_state_reg ( .D(Plaintext_s1[23]), 
        .CK(clk), .Q(new_AGEMA_signal_2237), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1050_s_current_state_reg ( .D(Plaintext_s0[26]), 
        .CK(clk), .Q(new_AGEMA_signal_2239), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1052_s_current_state_reg ( .D(Plaintext_s1[26]), 
        .CK(clk), .Q(new_AGEMA_signal_2241), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1054_s_current_state_reg ( .D(Plaintext_s0[27]), 
        .CK(clk), .Q(new_AGEMA_signal_2243), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1056_s_current_state_reg ( .D(Plaintext_s1[27]), 
        .CK(clk), .Q(new_AGEMA_signal_2245), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1058_s_current_state_reg ( .D(Plaintext_s0[30]), 
        .CK(clk), .Q(new_AGEMA_signal_2247), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1060_s_current_state_reg ( .D(Plaintext_s1[30]), 
        .CK(clk), .Q(new_AGEMA_signal_2249), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1062_s_current_state_reg ( .D(Plaintext_s0[31]), 
        .CK(clk), .Q(new_AGEMA_signal_2251), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1064_s_current_state_reg ( .D(Plaintext_s1[31]), 
        .CK(clk), .Q(new_AGEMA_signal_2253), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1066_s_current_state_reg ( .D(Plaintext_s0[34]), 
        .CK(clk), .Q(new_AGEMA_signal_2255), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1068_s_current_state_reg ( .D(Plaintext_s1[34]), 
        .CK(clk), .Q(new_AGEMA_signal_2257), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1070_s_current_state_reg ( .D(Plaintext_s0[35]), 
        .CK(clk), .Q(new_AGEMA_signal_2259), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1072_s_current_state_reg ( .D(Plaintext_s1[35]), 
        .CK(clk), .Q(new_AGEMA_signal_2261), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1074_s_current_state_reg ( .D(Plaintext_s0[38]), 
        .CK(clk), .Q(new_AGEMA_signal_2263), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1076_s_current_state_reg ( .D(Plaintext_s1[38]), 
        .CK(clk), .Q(new_AGEMA_signal_2265), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1078_s_current_state_reg ( .D(Plaintext_s0[39]), 
        .CK(clk), .Q(new_AGEMA_signal_2267), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1080_s_current_state_reg ( .D(Plaintext_s1[39]), 
        .CK(clk), .Q(new_AGEMA_signal_2269), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1082_s_current_state_reg ( .D(Plaintext_s0[42]), 
        .CK(clk), .Q(new_AGEMA_signal_2271), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1084_s_current_state_reg ( .D(Plaintext_s1[42]), 
        .CK(clk), .Q(new_AGEMA_signal_2273), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1086_s_current_state_reg ( .D(Plaintext_s0[43]), 
        .CK(clk), .Q(new_AGEMA_signal_2275), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1088_s_current_state_reg ( .D(Plaintext_s1[43]), 
        .CK(clk), .Q(new_AGEMA_signal_2277), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1090_s_current_state_reg ( .D(Plaintext_s0[46]), 
        .CK(clk), .Q(new_AGEMA_signal_2279), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1092_s_current_state_reg ( .D(Plaintext_s1[46]), 
        .CK(clk), .Q(new_AGEMA_signal_2281), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1094_s_current_state_reg ( .D(Plaintext_s0[47]), 
        .CK(clk), .Q(new_AGEMA_signal_2283), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1096_s_current_state_reg ( .D(Plaintext_s1[47]), 
        .CK(clk), .Q(new_AGEMA_signal_2285), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1098_s_current_state_reg ( .D(Plaintext_s0[50]), 
        .CK(clk), .Q(new_AGEMA_signal_2287), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1100_s_current_state_reg ( .D(Plaintext_s1[50]), 
        .CK(clk), .Q(new_AGEMA_signal_2289), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1102_s_current_state_reg ( .D(Plaintext_s0[51]), 
        .CK(clk), .Q(new_AGEMA_signal_2291), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1104_s_current_state_reg ( .D(Plaintext_s1[51]), 
        .CK(clk), .Q(new_AGEMA_signal_2293), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1106_s_current_state_reg ( .D(Plaintext_s0[54]), 
        .CK(clk), .Q(new_AGEMA_signal_2295), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1108_s_current_state_reg ( .D(Plaintext_s1[54]), 
        .CK(clk), .Q(new_AGEMA_signal_2297), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1110_s_current_state_reg ( .D(Plaintext_s0[55]), 
        .CK(clk), .Q(new_AGEMA_signal_2299), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1112_s_current_state_reg ( .D(Plaintext_s1[55]), 
        .CK(clk), .Q(new_AGEMA_signal_2301), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1114_s_current_state_reg ( .D(Plaintext_s0[58]), 
        .CK(clk), .Q(new_AGEMA_signal_2303), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1116_s_current_state_reg ( .D(Plaintext_s1[58]), 
        .CK(clk), .Q(new_AGEMA_signal_2305), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1118_s_current_state_reg ( .D(Plaintext_s0[59]), 
        .CK(clk), .Q(new_AGEMA_signal_2307), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1120_s_current_state_reg ( .D(Plaintext_s1[59]), 
        .CK(clk), .Q(new_AGEMA_signal_2309), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1122_s_current_state_reg ( .D(Plaintext_s0[62]), 
        .CK(clk), .Q(new_AGEMA_signal_2311), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1124_s_current_state_reg ( .D(Plaintext_s1[62]), 
        .CK(clk), .Q(new_AGEMA_signal_2313), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1126_s_current_state_reg ( .D(Plaintext_s0[63]), 
        .CK(clk), .Q(new_AGEMA_signal_2315), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1128_s_current_state_reg ( .D(Plaintext_s1[63]), 
        .CK(clk), .Q(new_AGEMA_signal_2317), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1130_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_Q0), .CK(clk), .Q(new_AGEMA_signal_2319), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1132_s_current_state_reg ( .D(
        new_AGEMA_signal_1453), .CK(clk), .Q(new_AGEMA_signal_2321), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1134_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_L1), .CK(clk), .Q(new_AGEMA_signal_2323), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1136_s_current_state_reg ( .D(
        new_AGEMA_signal_1550), .CK(clk), .Q(new_AGEMA_signal_2325), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1138_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2327), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1140_s_current_state_reg ( .D(
        new_AGEMA_signal_1169), .CK(clk), .Q(new_AGEMA_signal_2329), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1142_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2331), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1144_s_current_state_reg ( .D(
        new_AGEMA_signal_1167), .CK(clk), .Q(new_AGEMA_signal_2333), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1146_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_Q0), .CK(clk), .Q(new_AGEMA_signal_2335), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1148_s_current_state_reg ( .D(
        new_AGEMA_signal_1459), .CK(clk), .Q(new_AGEMA_signal_2337), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1150_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_L1), .CK(clk), .Q(new_AGEMA_signal_2339), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1152_s_current_state_reg ( .D(
        new_AGEMA_signal_1553), .CK(clk), .Q(new_AGEMA_signal_2341), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1154_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2343), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1156_s_current_state_reg ( .D(
        new_AGEMA_signal_1175), .CK(clk), .Q(new_AGEMA_signal_2345), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1158_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2347), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1160_s_current_state_reg ( .D(
        new_AGEMA_signal_1173), .CK(clk), .Q(new_AGEMA_signal_2349), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1162_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_Q0), .CK(clk), .Q(new_AGEMA_signal_2351), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1164_s_current_state_reg ( .D(
        new_AGEMA_signal_1465), .CK(clk), .Q(new_AGEMA_signal_2353), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1166_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_L1), .CK(clk), .Q(new_AGEMA_signal_2355), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1168_s_current_state_reg ( .D(
        new_AGEMA_signal_1556), .CK(clk), .Q(new_AGEMA_signal_2357), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1170_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2359), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1172_s_current_state_reg ( .D(
        new_AGEMA_signal_1181), .CK(clk), .Q(new_AGEMA_signal_2361), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1174_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2363), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1176_s_current_state_reg ( .D(
        new_AGEMA_signal_1179), .CK(clk), .Q(new_AGEMA_signal_2365), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1178_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_Q0), .CK(clk), .Q(new_AGEMA_signal_2367), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1180_s_current_state_reg ( .D(
        new_AGEMA_signal_1471), .CK(clk), .Q(new_AGEMA_signal_2369), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1182_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_L1), .CK(clk), .Q(new_AGEMA_signal_2371), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1184_s_current_state_reg ( .D(
        new_AGEMA_signal_1559), .CK(clk), .Q(new_AGEMA_signal_2373), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1186_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2375), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1188_s_current_state_reg ( .D(
        new_AGEMA_signal_1187), .CK(clk), .Q(new_AGEMA_signal_2377), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1190_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2379), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1192_s_current_state_reg ( .D(
        new_AGEMA_signal_1185), .CK(clk), .Q(new_AGEMA_signal_2381), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1194_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_Q0), .CK(clk), .Q(new_AGEMA_signal_2383), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1196_s_current_state_reg ( .D(
        new_AGEMA_signal_1477), .CK(clk), .Q(new_AGEMA_signal_2385), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1198_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_L1), .CK(clk), .Q(new_AGEMA_signal_2387), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1200_s_current_state_reg ( .D(
        new_AGEMA_signal_1562), .CK(clk), .Q(new_AGEMA_signal_2389), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1202_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2391), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1204_s_current_state_reg ( .D(
        new_AGEMA_signal_1193), .CK(clk), .Q(new_AGEMA_signal_2393), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1206_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2395), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1208_s_current_state_reg ( .D(
        new_AGEMA_signal_1191), .CK(clk), .Q(new_AGEMA_signal_2397), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1210_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_Q0), .CK(clk), .Q(new_AGEMA_signal_2399), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1212_s_current_state_reg ( .D(
        new_AGEMA_signal_1483), .CK(clk), .Q(new_AGEMA_signal_2401), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1214_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_L1), .CK(clk), .Q(new_AGEMA_signal_2403), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1216_s_current_state_reg ( .D(
        new_AGEMA_signal_1565), .CK(clk), .Q(new_AGEMA_signal_2405), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1218_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2407), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1220_s_current_state_reg ( .D(
        new_AGEMA_signal_1199), .CK(clk), .Q(new_AGEMA_signal_2409), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1222_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2411), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1224_s_current_state_reg ( .D(
        new_AGEMA_signal_1197), .CK(clk), .Q(new_AGEMA_signal_2413), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1226_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_Q0), .CK(clk), .Q(new_AGEMA_signal_2415), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1228_s_current_state_reg ( .D(
        new_AGEMA_signal_1489), .CK(clk), .Q(new_AGEMA_signal_2417), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1230_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_L1), .CK(clk), .Q(new_AGEMA_signal_2419), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1232_s_current_state_reg ( .D(
        new_AGEMA_signal_1568), .CK(clk), .Q(new_AGEMA_signal_2421), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1234_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2423), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1236_s_current_state_reg ( .D(
        new_AGEMA_signal_1205), .CK(clk), .Q(new_AGEMA_signal_2425), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1238_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2427), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1240_s_current_state_reg ( .D(
        new_AGEMA_signal_1203), .CK(clk), .Q(new_AGEMA_signal_2429), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1242_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_Q0), .CK(clk), .Q(new_AGEMA_signal_2431), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1244_s_current_state_reg ( .D(
        new_AGEMA_signal_1495), .CK(clk), .Q(new_AGEMA_signal_2433), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1246_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_L1), .CK(clk), .Q(new_AGEMA_signal_2435), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1248_s_current_state_reg ( .D(
        new_AGEMA_signal_1571), .CK(clk), .Q(new_AGEMA_signal_2437), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1250_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2439), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1252_s_current_state_reg ( .D(
        new_AGEMA_signal_1211), .CK(clk), .Q(new_AGEMA_signal_2441), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1254_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2443), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1256_s_current_state_reg ( .D(
        new_AGEMA_signal_1209), .CK(clk), .Q(new_AGEMA_signal_2445), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1258_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_Q0), .CK(clk), .Q(new_AGEMA_signal_2447), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1260_s_current_state_reg ( .D(
        new_AGEMA_signal_1501), .CK(clk), .Q(new_AGEMA_signal_2449), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1262_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_L1), .CK(clk), .Q(new_AGEMA_signal_2451), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1264_s_current_state_reg ( .D(
        new_AGEMA_signal_1574), .CK(clk), .Q(new_AGEMA_signal_2453), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1266_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2455), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1268_s_current_state_reg ( .D(
        new_AGEMA_signal_1217), .CK(clk), .Q(new_AGEMA_signal_2457), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1270_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2459), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1272_s_current_state_reg ( .D(
        new_AGEMA_signal_1215), .CK(clk), .Q(new_AGEMA_signal_2461), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1274_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_Q0), .CK(clk), .Q(new_AGEMA_signal_2463), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1276_s_current_state_reg ( .D(
        new_AGEMA_signal_1507), .CK(clk), .Q(new_AGEMA_signal_2465), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1278_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_L1), .CK(clk), .Q(new_AGEMA_signal_2467), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1280_s_current_state_reg ( .D(
        new_AGEMA_signal_1577), .CK(clk), .Q(new_AGEMA_signal_2469), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1282_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2471), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1284_s_current_state_reg ( .D(
        new_AGEMA_signal_1223), .CK(clk), .Q(new_AGEMA_signal_2473), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1286_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2475), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1288_s_current_state_reg ( .D(
        new_AGEMA_signal_1221), .CK(clk), .Q(new_AGEMA_signal_2477), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1290_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_Q0), .CK(clk), .Q(new_AGEMA_signal_2479), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1292_s_current_state_reg ( .D(
        new_AGEMA_signal_1513), .CK(clk), .Q(new_AGEMA_signal_2481), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1294_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_L1), .CK(clk), .Q(new_AGEMA_signal_2483), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1296_s_current_state_reg ( .D(
        new_AGEMA_signal_1580), .CK(clk), .Q(new_AGEMA_signal_2485), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1298_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2487), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1300_s_current_state_reg ( .D(
        new_AGEMA_signal_1229), .CK(clk), .Q(new_AGEMA_signal_2489), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1302_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2491), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1304_s_current_state_reg ( .D(
        new_AGEMA_signal_1227), .CK(clk), .Q(new_AGEMA_signal_2493), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1306_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_Q0), .CK(clk), .Q(new_AGEMA_signal_2495), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1308_s_current_state_reg ( .D(
        new_AGEMA_signal_1519), .CK(clk), .Q(new_AGEMA_signal_2497), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1310_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_L1), .CK(clk), .Q(new_AGEMA_signal_2499), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1312_s_current_state_reg ( .D(
        new_AGEMA_signal_1583), .CK(clk), .Q(new_AGEMA_signal_2501), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1314_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2503), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1316_s_current_state_reg ( .D(
        new_AGEMA_signal_1235), .CK(clk), .Q(new_AGEMA_signal_2505), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1318_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2507), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1320_s_current_state_reg ( .D(
        new_AGEMA_signal_1233), .CK(clk), .Q(new_AGEMA_signal_2509), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1322_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_Q0), .CK(clk), .Q(new_AGEMA_signal_2511), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1324_s_current_state_reg ( .D(
        new_AGEMA_signal_1525), .CK(clk), .Q(new_AGEMA_signal_2513), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1326_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_L1), .CK(clk), .Q(new_AGEMA_signal_2515), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1328_s_current_state_reg ( .D(
        new_AGEMA_signal_1586), .CK(clk), .Q(new_AGEMA_signal_2517), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1330_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2519), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1332_s_current_state_reg ( .D(
        new_AGEMA_signal_1241), .CK(clk), .Q(new_AGEMA_signal_2521), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1334_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2523), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1336_s_current_state_reg ( .D(
        new_AGEMA_signal_1239), .CK(clk), .Q(new_AGEMA_signal_2525), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1338_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_Q0), .CK(clk), .Q(new_AGEMA_signal_2527), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1340_s_current_state_reg ( .D(
        new_AGEMA_signal_1531), .CK(clk), .Q(new_AGEMA_signal_2529), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1342_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_L1), .CK(clk), .Q(new_AGEMA_signal_2531), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1344_s_current_state_reg ( .D(
        new_AGEMA_signal_1589), .CK(clk), .Q(new_AGEMA_signal_2533), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1346_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2535), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1348_s_current_state_reg ( .D(
        new_AGEMA_signal_1247), .CK(clk), .Q(new_AGEMA_signal_2537), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1350_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2539), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1352_s_current_state_reg ( .D(
        new_AGEMA_signal_1245), .CK(clk), .Q(new_AGEMA_signal_2541), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1354_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_Q0), .CK(clk), .Q(new_AGEMA_signal_2543), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1356_s_current_state_reg ( .D(
        new_AGEMA_signal_1537), .CK(clk), .Q(new_AGEMA_signal_2545), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1358_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_L1), .CK(clk), .Q(new_AGEMA_signal_2547), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1360_s_current_state_reg ( .D(
        new_AGEMA_signal_1592), .CK(clk), .Q(new_AGEMA_signal_2549), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1362_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2551), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1364_s_current_state_reg ( .D(
        new_AGEMA_signal_1253), .CK(clk), .Q(new_AGEMA_signal_2553), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1366_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2555), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1368_s_current_state_reg ( .D(
        new_AGEMA_signal_1251), .CK(clk), .Q(new_AGEMA_signal_2557), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1370_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_Q0), .CK(clk), .Q(new_AGEMA_signal_2559), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1372_s_current_state_reg ( .D(
        new_AGEMA_signal_1543), .CK(clk), .Q(new_AGEMA_signal_2561), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1374_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_L1), .CK(clk), .Q(new_AGEMA_signal_2563), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1376_s_current_state_reg ( .D(
        new_AGEMA_signal_1595), .CK(clk), .Q(new_AGEMA_signal_2565), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1378_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_XX_2_), .CK(clk), .Q(new_AGEMA_signal_2567), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1380_s_current_state_reg ( .D(
        new_AGEMA_signal_1259), .CK(clk), .Q(new_AGEMA_signal_2569), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1382_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_XX_1_), .CK(clk), .Q(new_AGEMA_signal_2571), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1384_s_current_state_reg ( .D(
        new_AGEMA_signal_1257), .CK(clk), .Q(new_AGEMA_signal_2573), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1386_s_current_state_reg ( .D(FSMUpdate[3]), 
        .CK(clk), .Q(new_AGEMA_signal_2575), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1388_s_current_state_reg ( .D(FSMUpdate[4]), 
        .CK(clk), .Q(new_AGEMA_signal_2577), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1390_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[2]), .CK(clk), .Q(new_AGEMA_signal_2579), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1392_s_current_state_reg ( .D(
        new_AGEMA_signal_1266), .CK(clk), .Q(new_AGEMA_signal_2581), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1394_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[3]), .CK(clk), .Q(new_AGEMA_signal_2583), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1396_s_current_state_reg ( .D(
        new_AGEMA_signal_1269), .CK(clk), .Q(new_AGEMA_signal_2585), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1398_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[6]), .CK(clk), .Q(new_AGEMA_signal_2587), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1400_s_current_state_reg ( .D(
        new_AGEMA_signal_1278), .CK(clk), .Q(new_AGEMA_signal_2589), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1402_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[7]), .CK(clk), .Q(new_AGEMA_signal_2591), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1404_s_current_state_reg ( .D(
        new_AGEMA_signal_1281), .CK(clk), .Q(new_AGEMA_signal_2593), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1406_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[10]), .CK(clk), .Q(
        new_AGEMA_signal_2595), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1408_s_current_state_reg ( .D(
        new_AGEMA_signal_1290), .CK(clk), .Q(new_AGEMA_signal_2597), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1410_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[11]), .CK(clk), .Q(
        new_AGEMA_signal_2599), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1412_s_current_state_reg ( .D(
        new_AGEMA_signal_1293), .CK(clk), .Q(new_AGEMA_signal_2601), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1414_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[14]), .CK(clk), .Q(
        new_AGEMA_signal_2603), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1416_s_current_state_reg ( .D(
        new_AGEMA_signal_1302), .CK(clk), .Q(new_AGEMA_signal_2605), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1418_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[15]), .CK(clk), .Q(
        new_AGEMA_signal_2607), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1420_s_current_state_reg ( .D(
        new_AGEMA_signal_1305), .CK(clk), .Q(new_AGEMA_signal_2609), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1422_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[18]), .CK(clk), .Q(
        new_AGEMA_signal_2611), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1424_s_current_state_reg ( .D(
        new_AGEMA_signal_1314), .CK(clk), .Q(new_AGEMA_signal_2613), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1426_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[19]), .CK(clk), .Q(
        new_AGEMA_signal_2615), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1428_s_current_state_reg ( .D(
        new_AGEMA_signal_1317), .CK(clk), .Q(new_AGEMA_signal_2617), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1430_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[22]), .CK(clk), .Q(
        new_AGEMA_signal_2619), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1432_s_current_state_reg ( .D(
        new_AGEMA_signal_1326), .CK(clk), .Q(new_AGEMA_signal_2621), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1434_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[23]), .CK(clk), .Q(
        new_AGEMA_signal_2623), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1436_s_current_state_reg ( .D(
        new_AGEMA_signal_1329), .CK(clk), .Q(new_AGEMA_signal_2625), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1438_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[26]), .CK(clk), .Q(
        new_AGEMA_signal_2627), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1440_s_current_state_reg ( .D(
        new_AGEMA_signal_1338), .CK(clk), .Q(new_AGEMA_signal_2629), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1442_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[27]), .CK(clk), .Q(
        new_AGEMA_signal_2631), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1444_s_current_state_reg ( .D(
        new_AGEMA_signal_1341), .CK(clk), .Q(new_AGEMA_signal_2633), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1446_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[30]), .CK(clk), .Q(
        new_AGEMA_signal_2635), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1448_s_current_state_reg ( .D(
        new_AGEMA_signal_1350), .CK(clk), .Q(new_AGEMA_signal_2637), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1450_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[31]), .CK(clk), .Q(
        new_AGEMA_signal_2639), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1452_s_current_state_reg ( .D(
        new_AGEMA_signal_1353), .CK(clk), .Q(new_AGEMA_signal_2641), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1456_s_current_state_reg ( .D(Plaintext_s0[0]), 
        .CK(clk), .Q(new_AGEMA_signal_2645), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1460_s_current_state_reg ( .D(Plaintext_s1[0]), 
        .CK(clk), .Q(new_AGEMA_signal_2649), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1464_s_current_state_reg ( .D(Plaintext_s0[1]), 
        .CK(clk), .Q(new_AGEMA_signal_2653), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1468_s_current_state_reg ( .D(Plaintext_s1[1]), 
        .CK(clk), .Q(new_AGEMA_signal_2657), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1472_s_current_state_reg ( .D(Plaintext_s0[4]), 
        .CK(clk), .Q(new_AGEMA_signal_2661), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1476_s_current_state_reg ( .D(Plaintext_s1[4]), 
        .CK(clk), .Q(new_AGEMA_signal_2665), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1480_s_current_state_reg ( .D(Plaintext_s0[5]), 
        .CK(clk), .Q(new_AGEMA_signal_2669), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1484_s_current_state_reg ( .D(Plaintext_s1[5]), 
        .CK(clk), .Q(new_AGEMA_signal_2673), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1488_s_current_state_reg ( .D(Plaintext_s0[8]), 
        .CK(clk), .Q(new_AGEMA_signal_2677), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1492_s_current_state_reg ( .D(Plaintext_s1[8]), 
        .CK(clk), .Q(new_AGEMA_signal_2681), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1496_s_current_state_reg ( .D(Plaintext_s0[9]), 
        .CK(clk), .Q(new_AGEMA_signal_2685), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1500_s_current_state_reg ( .D(Plaintext_s1[9]), 
        .CK(clk), .Q(new_AGEMA_signal_2689), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1504_s_current_state_reg ( .D(Plaintext_s0[12]), 
        .CK(clk), .Q(new_AGEMA_signal_2693), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1508_s_current_state_reg ( .D(Plaintext_s1[12]), 
        .CK(clk), .Q(new_AGEMA_signal_2697), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1512_s_current_state_reg ( .D(Plaintext_s0[13]), 
        .CK(clk), .Q(new_AGEMA_signal_2701), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1516_s_current_state_reg ( .D(Plaintext_s1[13]), 
        .CK(clk), .Q(new_AGEMA_signal_2705), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1520_s_current_state_reg ( .D(Plaintext_s0[16]), 
        .CK(clk), .Q(new_AGEMA_signal_2709), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1524_s_current_state_reg ( .D(Plaintext_s1[16]), 
        .CK(clk), .Q(new_AGEMA_signal_2713), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1528_s_current_state_reg ( .D(Plaintext_s0[17]), 
        .CK(clk), .Q(new_AGEMA_signal_2717), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1532_s_current_state_reg ( .D(Plaintext_s1[17]), 
        .CK(clk), .Q(new_AGEMA_signal_2721), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1536_s_current_state_reg ( .D(Plaintext_s0[20]), 
        .CK(clk), .Q(new_AGEMA_signal_2725), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1540_s_current_state_reg ( .D(Plaintext_s1[20]), 
        .CK(clk), .Q(new_AGEMA_signal_2729), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1544_s_current_state_reg ( .D(Plaintext_s0[21]), 
        .CK(clk), .Q(new_AGEMA_signal_2733), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1548_s_current_state_reg ( .D(Plaintext_s1[21]), 
        .CK(clk), .Q(new_AGEMA_signal_2737), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1552_s_current_state_reg ( .D(Plaintext_s0[24]), 
        .CK(clk), .Q(new_AGEMA_signal_2741), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1556_s_current_state_reg ( .D(Plaintext_s1[24]), 
        .CK(clk), .Q(new_AGEMA_signal_2745), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1560_s_current_state_reg ( .D(Plaintext_s0[25]), 
        .CK(clk), .Q(new_AGEMA_signal_2749), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1564_s_current_state_reg ( .D(Plaintext_s1[25]), 
        .CK(clk), .Q(new_AGEMA_signal_2753), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1568_s_current_state_reg ( .D(Plaintext_s0[28]), 
        .CK(clk), .Q(new_AGEMA_signal_2757), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1572_s_current_state_reg ( .D(Plaintext_s1[28]), 
        .CK(clk), .Q(new_AGEMA_signal_2761), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1576_s_current_state_reg ( .D(Plaintext_s0[29]), 
        .CK(clk), .Q(new_AGEMA_signal_2765), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1580_s_current_state_reg ( .D(Plaintext_s1[29]), 
        .CK(clk), .Q(new_AGEMA_signal_2769), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1584_s_current_state_reg ( .D(Plaintext_s0[32]), 
        .CK(clk), .Q(new_AGEMA_signal_2773), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1588_s_current_state_reg ( .D(Plaintext_s1[32]), 
        .CK(clk), .Q(new_AGEMA_signal_2777), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1592_s_current_state_reg ( .D(Plaintext_s0[33]), 
        .CK(clk), .Q(new_AGEMA_signal_2781), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1596_s_current_state_reg ( .D(Plaintext_s1[33]), 
        .CK(clk), .Q(new_AGEMA_signal_2785), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1600_s_current_state_reg ( .D(Plaintext_s0[36]), 
        .CK(clk), .Q(new_AGEMA_signal_2789), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1604_s_current_state_reg ( .D(Plaintext_s1[36]), 
        .CK(clk), .Q(new_AGEMA_signal_2793), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1608_s_current_state_reg ( .D(Plaintext_s0[37]), 
        .CK(clk), .Q(new_AGEMA_signal_2797), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1612_s_current_state_reg ( .D(Plaintext_s1[37]), 
        .CK(clk), .Q(new_AGEMA_signal_2801), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1616_s_current_state_reg ( .D(Plaintext_s0[40]), 
        .CK(clk), .Q(new_AGEMA_signal_2805), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1620_s_current_state_reg ( .D(Plaintext_s1[40]), 
        .CK(clk), .Q(new_AGEMA_signal_2809), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1624_s_current_state_reg ( .D(Plaintext_s0[41]), 
        .CK(clk), .Q(new_AGEMA_signal_2813), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1628_s_current_state_reg ( .D(Plaintext_s1[41]), 
        .CK(clk), .Q(new_AGEMA_signal_2817), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1632_s_current_state_reg ( .D(Plaintext_s0[44]), 
        .CK(clk), .Q(new_AGEMA_signal_2821), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1636_s_current_state_reg ( .D(Plaintext_s1[44]), 
        .CK(clk), .Q(new_AGEMA_signal_2825), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1640_s_current_state_reg ( .D(Plaintext_s0[45]), 
        .CK(clk), .Q(new_AGEMA_signal_2829), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1644_s_current_state_reg ( .D(Plaintext_s1[45]), 
        .CK(clk), .Q(new_AGEMA_signal_2833), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1648_s_current_state_reg ( .D(Plaintext_s0[48]), 
        .CK(clk), .Q(new_AGEMA_signal_2837), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1652_s_current_state_reg ( .D(Plaintext_s1[48]), 
        .CK(clk), .Q(new_AGEMA_signal_2841), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1656_s_current_state_reg ( .D(Plaintext_s0[49]), 
        .CK(clk), .Q(new_AGEMA_signal_2845), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1660_s_current_state_reg ( .D(Plaintext_s1[49]), 
        .CK(clk), .Q(new_AGEMA_signal_2849), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1664_s_current_state_reg ( .D(Plaintext_s0[52]), 
        .CK(clk), .Q(new_AGEMA_signal_2853), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1668_s_current_state_reg ( .D(Plaintext_s1[52]), 
        .CK(clk), .Q(new_AGEMA_signal_2857), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1672_s_current_state_reg ( .D(Plaintext_s0[53]), 
        .CK(clk), .Q(new_AGEMA_signal_2861), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1676_s_current_state_reg ( .D(Plaintext_s1[53]), 
        .CK(clk), .Q(new_AGEMA_signal_2865), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1680_s_current_state_reg ( .D(Plaintext_s0[56]), 
        .CK(clk), .Q(new_AGEMA_signal_2869), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1684_s_current_state_reg ( .D(Plaintext_s1[56]), 
        .CK(clk), .Q(new_AGEMA_signal_2873), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1688_s_current_state_reg ( .D(Plaintext_s0[57]), 
        .CK(clk), .Q(new_AGEMA_signal_2877), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1692_s_current_state_reg ( .D(Plaintext_s1[57]), 
        .CK(clk), .Q(new_AGEMA_signal_2881), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1696_s_current_state_reg ( .D(Plaintext_s0[60]), 
        .CK(clk), .Q(new_AGEMA_signal_2885), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1700_s_current_state_reg ( .D(Plaintext_s1[60]), 
        .CK(clk), .Q(new_AGEMA_signal_2889), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1704_s_current_state_reg ( .D(Plaintext_s0[61]), 
        .CK(clk), .Q(new_AGEMA_signal_2893), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1708_s_current_state_reg ( .D(Plaintext_s1[61]), 
        .CK(clk), .Q(new_AGEMA_signal_2897), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1712_s_current_state_reg ( .D(Ciphertext_s0[1]), 
        .CK(clk), .Q(new_AGEMA_signal_2901), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1714_s_current_state_reg ( .D(Ciphertext_s1[1]), 
        .CK(clk), .Q(new_AGEMA_signal_2903), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1720_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_Q6), .CK(clk), .Q(new_AGEMA_signal_2909), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1722_s_current_state_reg ( .D(
        new_AGEMA_signal_1456), .CK(clk), .Q(new_AGEMA_signal_2911), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1724_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_L2), .CK(clk), .Q(new_AGEMA_signal_2913), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1728_s_current_state_reg ( .D(
        new_AGEMA_signal_1457), .CK(clk), .Q(new_AGEMA_signal_2917), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1736_s_current_state_reg ( .D(Ciphertext_s0[5]), 
        .CK(clk), .Q(new_AGEMA_signal_2925), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1738_s_current_state_reg ( .D(Ciphertext_s1[5]), 
        .CK(clk), .Q(new_AGEMA_signal_2927), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1744_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_Q6), .CK(clk), .Q(new_AGEMA_signal_2933), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1746_s_current_state_reg ( .D(
        new_AGEMA_signal_1462), .CK(clk), .Q(new_AGEMA_signal_2935), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1748_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_L2), .CK(clk), .Q(new_AGEMA_signal_2937), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1752_s_current_state_reg ( .D(
        new_AGEMA_signal_1463), .CK(clk), .Q(new_AGEMA_signal_2941), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1760_s_current_state_reg ( .D(Ciphertext_s0[9]), 
        .CK(clk), .Q(new_AGEMA_signal_2949), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1762_s_current_state_reg ( .D(Ciphertext_s1[9]), 
        .CK(clk), .Q(new_AGEMA_signal_2951), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1768_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_Q6), .CK(clk), .Q(new_AGEMA_signal_2957), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1770_s_current_state_reg ( .D(
        new_AGEMA_signal_1468), .CK(clk), .Q(new_AGEMA_signal_2959), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1772_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_L2), .CK(clk), .Q(new_AGEMA_signal_2961), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1776_s_current_state_reg ( .D(
        new_AGEMA_signal_1469), .CK(clk), .Q(new_AGEMA_signal_2965), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1784_s_current_state_reg ( .D(Ciphertext_s0[13]), 
        .CK(clk), .Q(new_AGEMA_signal_2973), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1786_s_current_state_reg ( .D(Ciphertext_s1[13]), 
        .CK(clk), .Q(new_AGEMA_signal_2975), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1792_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_Q6), .CK(clk), .Q(new_AGEMA_signal_2981), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1794_s_current_state_reg ( .D(
        new_AGEMA_signal_1474), .CK(clk), .Q(new_AGEMA_signal_2983), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1796_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_L2), .CK(clk), .Q(new_AGEMA_signal_2985), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1800_s_current_state_reg ( .D(
        new_AGEMA_signal_1475), .CK(clk), .Q(new_AGEMA_signal_2989), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1808_s_current_state_reg ( .D(Ciphertext_s0[17]), 
        .CK(clk), .Q(new_AGEMA_signal_2997), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1810_s_current_state_reg ( .D(Ciphertext_s1[17]), 
        .CK(clk), .Q(new_AGEMA_signal_2999), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1816_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_Q6), .CK(clk), .Q(new_AGEMA_signal_3005), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1818_s_current_state_reg ( .D(
        new_AGEMA_signal_1480), .CK(clk), .Q(new_AGEMA_signal_3007), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1820_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_L2), .CK(clk), .Q(new_AGEMA_signal_3009), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1824_s_current_state_reg ( .D(
        new_AGEMA_signal_1481), .CK(clk), .Q(new_AGEMA_signal_3013), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1832_s_current_state_reg ( .D(Ciphertext_s0[21]), 
        .CK(clk), .Q(new_AGEMA_signal_3021), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1834_s_current_state_reg ( .D(Ciphertext_s1[21]), 
        .CK(clk), .Q(new_AGEMA_signal_3023), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1840_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_Q6), .CK(clk), .Q(new_AGEMA_signal_3029), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1842_s_current_state_reg ( .D(
        new_AGEMA_signal_1486), .CK(clk), .Q(new_AGEMA_signal_3031), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1844_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_L2), .CK(clk), .Q(new_AGEMA_signal_3033), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1848_s_current_state_reg ( .D(
        new_AGEMA_signal_1487), .CK(clk), .Q(new_AGEMA_signal_3037), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1856_s_current_state_reg ( .D(Ciphertext_s0[25]), 
        .CK(clk), .Q(new_AGEMA_signal_3045), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1858_s_current_state_reg ( .D(Ciphertext_s1[25]), 
        .CK(clk), .Q(new_AGEMA_signal_3047), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1864_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_Q6), .CK(clk), .Q(new_AGEMA_signal_3053), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1866_s_current_state_reg ( .D(
        new_AGEMA_signal_1492), .CK(clk), .Q(new_AGEMA_signal_3055), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1868_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_L2), .CK(clk), .Q(new_AGEMA_signal_3057), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1872_s_current_state_reg ( .D(
        new_AGEMA_signal_1493), .CK(clk), .Q(new_AGEMA_signal_3061), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1880_s_current_state_reg ( .D(Ciphertext_s0[29]), 
        .CK(clk), .Q(new_AGEMA_signal_3069), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1882_s_current_state_reg ( .D(Ciphertext_s1[29]), 
        .CK(clk), .Q(new_AGEMA_signal_3071), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1888_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_Q6), .CK(clk), .Q(new_AGEMA_signal_3077), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1890_s_current_state_reg ( .D(
        new_AGEMA_signal_1498), .CK(clk), .Q(new_AGEMA_signal_3079), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1892_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_L2), .CK(clk), .Q(new_AGEMA_signal_3081), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1896_s_current_state_reg ( .D(
        new_AGEMA_signal_1499), .CK(clk), .Q(new_AGEMA_signal_3085), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1904_s_current_state_reg ( .D(Ciphertext_s0[33]), 
        .CK(clk), .Q(new_AGEMA_signal_3093), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1906_s_current_state_reg ( .D(Ciphertext_s1[33]), 
        .CK(clk), .Q(new_AGEMA_signal_3095), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1912_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_Q6), .CK(clk), .Q(new_AGEMA_signal_3101), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1914_s_current_state_reg ( .D(
        new_AGEMA_signal_1504), .CK(clk), .Q(new_AGEMA_signal_3103), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1916_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_L2), .CK(clk), .Q(new_AGEMA_signal_3105), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1920_s_current_state_reg ( .D(
        new_AGEMA_signal_1505), .CK(clk), .Q(new_AGEMA_signal_3109), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1928_s_current_state_reg ( .D(Ciphertext_s0[37]), 
        .CK(clk), .Q(new_AGEMA_signal_3117), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1930_s_current_state_reg ( .D(Ciphertext_s1[37]), 
        .CK(clk), .Q(new_AGEMA_signal_3119), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1936_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_Q6), .CK(clk), .Q(new_AGEMA_signal_3125), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1938_s_current_state_reg ( .D(
        new_AGEMA_signal_1510), .CK(clk), .Q(new_AGEMA_signal_3127), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1940_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_L2), .CK(clk), .Q(new_AGEMA_signal_3129), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1944_s_current_state_reg ( .D(
        new_AGEMA_signal_1511), .CK(clk), .Q(new_AGEMA_signal_3133), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1952_s_current_state_reg ( .D(Ciphertext_s0[41]), 
        .CK(clk), .Q(new_AGEMA_signal_3141), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1954_s_current_state_reg ( .D(Ciphertext_s1[41]), 
        .CK(clk), .Q(new_AGEMA_signal_3143), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1960_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_Q6), .CK(clk), .Q(new_AGEMA_signal_3149), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1962_s_current_state_reg ( .D(
        new_AGEMA_signal_1516), .CK(clk), .Q(new_AGEMA_signal_3151), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1964_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_L2), .CK(clk), .Q(new_AGEMA_signal_3153), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1968_s_current_state_reg ( .D(
        new_AGEMA_signal_1517), .CK(clk), .Q(new_AGEMA_signal_3157), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1976_s_current_state_reg ( .D(Ciphertext_s0[45]), 
        .CK(clk), .Q(new_AGEMA_signal_3165), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1978_s_current_state_reg ( .D(Ciphertext_s1[45]), 
        .CK(clk), .Q(new_AGEMA_signal_3167), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1984_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_Q6), .CK(clk), .Q(new_AGEMA_signal_3173), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1986_s_current_state_reg ( .D(
        new_AGEMA_signal_1522), .CK(clk), .Q(new_AGEMA_signal_3175), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1988_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_L2), .CK(clk), .Q(new_AGEMA_signal_3177), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1992_s_current_state_reg ( .D(
        new_AGEMA_signal_1523), .CK(clk), .Q(new_AGEMA_signal_3181), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2000_s_current_state_reg ( .D(Ciphertext_s0[49]), 
        .CK(clk), .Q(new_AGEMA_signal_3189), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2002_s_current_state_reg ( .D(Ciphertext_s1[49]), 
        .CK(clk), .Q(new_AGEMA_signal_3191), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2008_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_Q6), .CK(clk), .Q(new_AGEMA_signal_3197), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2010_s_current_state_reg ( .D(
        new_AGEMA_signal_1528), .CK(clk), .Q(new_AGEMA_signal_3199), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2012_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_L2), .CK(clk), .Q(new_AGEMA_signal_3201), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2016_s_current_state_reg ( .D(
        new_AGEMA_signal_1529), .CK(clk), .Q(new_AGEMA_signal_3205), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2024_s_current_state_reg ( .D(Ciphertext_s0[53]), 
        .CK(clk), .Q(new_AGEMA_signal_3213), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2026_s_current_state_reg ( .D(Ciphertext_s1[53]), 
        .CK(clk), .Q(new_AGEMA_signal_3215), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2032_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_Q6), .CK(clk), .Q(new_AGEMA_signal_3221), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2034_s_current_state_reg ( .D(
        new_AGEMA_signal_1534), .CK(clk), .Q(new_AGEMA_signal_3223), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2036_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_L2), .CK(clk), .Q(new_AGEMA_signal_3225), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2040_s_current_state_reg ( .D(
        new_AGEMA_signal_1535), .CK(clk), .Q(new_AGEMA_signal_3229), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2048_s_current_state_reg ( .D(Ciphertext_s0[57]), 
        .CK(clk), .Q(new_AGEMA_signal_3237), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2050_s_current_state_reg ( .D(Ciphertext_s1[57]), 
        .CK(clk), .Q(new_AGEMA_signal_3239), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2056_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_Q6), .CK(clk), .Q(new_AGEMA_signal_3245), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2058_s_current_state_reg ( .D(
        new_AGEMA_signal_1540), .CK(clk), .Q(new_AGEMA_signal_3247), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2060_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_L2), .CK(clk), .Q(new_AGEMA_signal_3249), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2064_s_current_state_reg ( .D(
        new_AGEMA_signal_1541), .CK(clk), .Q(new_AGEMA_signal_3253), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2072_s_current_state_reg ( .D(Ciphertext_s0[61]), 
        .CK(clk), .Q(new_AGEMA_signal_3261), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2074_s_current_state_reg ( .D(Ciphertext_s1[61]), 
        .CK(clk), .Q(new_AGEMA_signal_3263), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2080_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_Q6), .CK(clk), .Q(new_AGEMA_signal_3269), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2082_s_current_state_reg ( .D(
        new_AGEMA_signal_1546), .CK(clk), .Q(new_AGEMA_signal_3271), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2084_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_L2), .CK(clk), .Q(new_AGEMA_signal_3273), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2088_s_current_state_reg ( .D(
        new_AGEMA_signal_1547), .CK(clk), .Q(new_AGEMA_signal_3277), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2096_s_current_state_reg ( .D(FSMUpdate[1]), 
        .CK(clk), .Q(new_AGEMA_signal_3285), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2100_s_current_state_reg ( .D(FSM_1), .CK(clk), 
        .Q(new_AGEMA_signal_3289), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2104_s_current_state_reg ( .D(FSM[4]), .CK(clk), 
        .Q(new_AGEMA_signal_3293), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2108_s_current_state_reg ( .D(FSM[5]), .CK(clk), 
        .Q(new_AGEMA_signal_3297), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2112_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[0]), .CK(clk), .Q(new_AGEMA_signal_3301), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2116_s_current_state_reg ( .D(
        new_AGEMA_signal_1260), .CK(clk), .Q(new_AGEMA_signal_3305), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2120_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[1]), .CK(clk), .Q(new_AGEMA_signal_3309), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2124_s_current_state_reg ( .D(
        new_AGEMA_signal_1263), .CK(clk), .Q(new_AGEMA_signal_3313), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2128_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[4]), .CK(clk), .Q(new_AGEMA_signal_3317), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2132_s_current_state_reg ( .D(
        new_AGEMA_signal_1272), .CK(clk), .Q(new_AGEMA_signal_3321), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2136_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[5]), .CK(clk), .Q(new_AGEMA_signal_3325), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2140_s_current_state_reg ( .D(
        new_AGEMA_signal_1275), .CK(clk), .Q(new_AGEMA_signal_3329), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2144_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[8]), .CK(clk), .Q(new_AGEMA_signal_3333), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2148_s_current_state_reg ( .D(
        new_AGEMA_signal_1284), .CK(clk), .Q(new_AGEMA_signal_3337), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2152_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[9]), .CK(clk), .Q(new_AGEMA_signal_3341), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2156_s_current_state_reg ( .D(
        new_AGEMA_signal_1287), .CK(clk), .Q(new_AGEMA_signal_3345), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2160_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[12]), .CK(clk), .Q(
        new_AGEMA_signal_3349), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2164_s_current_state_reg ( .D(
        new_AGEMA_signal_1296), .CK(clk), .Q(new_AGEMA_signal_3353), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2168_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[13]), .CK(clk), .Q(
        new_AGEMA_signal_3357), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2172_s_current_state_reg ( .D(
        new_AGEMA_signal_1299), .CK(clk), .Q(new_AGEMA_signal_3361), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2176_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[16]), .CK(clk), .Q(
        new_AGEMA_signal_3365), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2180_s_current_state_reg ( .D(
        new_AGEMA_signal_1308), .CK(clk), .Q(new_AGEMA_signal_3369), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2184_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[17]), .CK(clk), .Q(
        new_AGEMA_signal_3373), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2188_s_current_state_reg ( .D(
        new_AGEMA_signal_1311), .CK(clk), .Q(new_AGEMA_signal_3377), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2192_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[20]), .CK(clk), .Q(
        new_AGEMA_signal_3381), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2196_s_current_state_reg ( .D(
        new_AGEMA_signal_1320), .CK(clk), .Q(new_AGEMA_signal_3385), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2200_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[21]), .CK(clk), .Q(
        new_AGEMA_signal_3389), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2204_s_current_state_reg ( .D(
        new_AGEMA_signal_1323), .CK(clk), .Q(new_AGEMA_signal_3393), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2208_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[24]), .CK(clk), .Q(
        new_AGEMA_signal_3397), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2212_s_current_state_reg ( .D(
        new_AGEMA_signal_1332), .CK(clk), .Q(new_AGEMA_signal_3401), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2216_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[25]), .CK(clk), .Q(
        new_AGEMA_signal_3405), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2220_s_current_state_reg ( .D(
        new_AGEMA_signal_1335), .CK(clk), .Q(new_AGEMA_signal_3409), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2224_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[28]), .CK(clk), .Q(
        new_AGEMA_signal_3413), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2228_s_current_state_reg ( .D(
        new_AGEMA_signal_1344), .CK(clk), .Q(new_AGEMA_signal_3417), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2232_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[29]), .CK(clk), .Q(
        new_AGEMA_signal_3421), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2236_s_current_state_reg ( .D(
        new_AGEMA_signal_1347), .CK(clk), .Q(new_AGEMA_signal_3425), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2368_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[63]), .CK(clk), .Q(
        new_AGEMA_signal_3557), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2372_s_current_state_reg ( .D(
        new_AGEMA_signal_1451), .CK(clk), .Q(new_AGEMA_signal_3561), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2376_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[62]), .CK(clk), .Q(
        new_AGEMA_signal_3565), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2380_s_current_state_reg ( .D(
        new_AGEMA_signal_1448), .CK(clk), .Q(new_AGEMA_signal_3569), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2384_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[61]), .CK(clk), .Q(
        new_AGEMA_signal_3573), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2388_s_current_state_reg ( .D(
        new_AGEMA_signal_1445), .CK(clk), .Q(new_AGEMA_signal_3577), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2392_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[60]), .CK(clk), .Q(
        new_AGEMA_signal_3581), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2396_s_current_state_reg ( .D(
        new_AGEMA_signal_1442), .CK(clk), .Q(new_AGEMA_signal_3585), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2400_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[59]), .CK(clk), .Q(
        new_AGEMA_signal_3589), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2404_s_current_state_reg ( .D(
        new_AGEMA_signal_1439), .CK(clk), .Q(new_AGEMA_signal_3593), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2408_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[58]), .CK(clk), .Q(
        new_AGEMA_signal_3597), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2412_s_current_state_reg ( .D(
        new_AGEMA_signal_1436), .CK(clk), .Q(new_AGEMA_signal_3601), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2416_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[57]), .CK(clk), .Q(
        new_AGEMA_signal_3605), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2420_s_current_state_reg ( .D(
        new_AGEMA_signal_1433), .CK(clk), .Q(new_AGEMA_signal_3609), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2424_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[56]), .CK(clk), .Q(
        new_AGEMA_signal_3613), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2428_s_current_state_reg ( .D(
        new_AGEMA_signal_1430), .CK(clk), .Q(new_AGEMA_signal_3617), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2432_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[55]), .CK(clk), .Q(
        new_AGEMA_signal_3621), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2436_s_current_state_reg ( .D(
        new_AGEMA_signal_1427), .CK(clk), .Q(new_AGEMA_signal_3625), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2440_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[54]), .CK(clk), .Q(
        new_AGEMA_signal_3629), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2444_s_current_state_reg ( .D(
        new_AGEMA_signal_1424), .CK(clk), .Q(new_AGEMA_signal_3633), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2448_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[53]), .CK(clk), .Q(
        new_AGEMA_signal_3637), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2452_s_current_state_reg ( .D(
        new_AGEMA_signal_1421), .CK(clk), .Q(new_AGEMA_signal_3641), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2456_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[52]), .CK(clk), .Q(
        new_AGEMA_signal_3645), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2460_s_current_state_reg ( .D(
        new_AGEMA_signal_1418), .CK(clk), .Q(new_AGEMA_signal_3649), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2464_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[51]), .CK(clk), .Q(
        new_AGEMA_signal_3653), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2468_s_current_state_reg ( .D(
        new_AGEMA_signal_1415), .CK(clk), .Q(new_AGEMA_signal_3657), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2472_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[50]), .CK(clk), .Q(
        new_AGEMA_signal_3661), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2476_s_current_state_reg ( .D(
        new_AGEMA_signal_1412), .CK(clk), .Q(new_AGEMA_signal_3665), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2480_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[49]), .CK(clk), .Q(
        new_AGEMA_signal_3669), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2484_s_current_state_reg ( .D(
        new_AGEMA_signal_1409), .CK(clk), .Q(new_AGEMA_signal_3673), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2488_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[48]), .CK(clk), .Q(
        new_AGEMA_signal_3677), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2492_s_current_state_reg ( .D(
        new_AGEMA_signal_1406), .CK(clk), .Q(new_AGEMA_signal_3681), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2496_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[47]), .CK(clk), .Q(
        new_AGEMA_signal_3685), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2500_s_current_state_reg ( .D(
        new_AGEMA_signal_1403), .CK(clk), .Q(new_AGEMA_signal_3689), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2504_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[46]), .CK(clk), .Q(
        new_AGEMA_signal_3693), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2508_s_current_state_reg ( .D(
        new_AGEMA_signal_1400), .CK(clk), .Q(new_AGEMA_signal_3697), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2512_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[45]), .CK(clk), .Q(
        new_AGEMA_signal_3701), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2516_s_current_state_reg ( .D(
        new_AGEMA_signal_1397), .CK(clk), .Q(new_AGEMA_signal_3705), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2520_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[44]), .CK(clk), .Q(
        new_AGEMA_signal_3709), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2524_s_current_state_reg ( .D(
        new_AGEMA_signal_1394), .CK(clk), .Q(new_AGEMA_signal_3713), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2528_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[43]), .CK(clk), .Q(
        new_AGEMA_signal_3717), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2532_s_current_state_reg ( .D(
        new_AGEMA_signal_1391), .CK(clk), .Q(new_AGEMA_signal_3721), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2536_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[42]), .CK(clk), .Q(
        new_AGEMA_signal_3725), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2540_s_current_state_reg ( .D(
        new_AGEMA_signal_1388), .CK(clk), .Q(new_AGEMA_signal_3729), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2544_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[41]), .CK(clk), .Q(
        new_AGEMA_signal_3733), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2548_s_current_state_reg ( .D(
        new_AGEMA_signal_1385), .CK(clk), .Q(new_AGEMA_signal_3737), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2552_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[40]), .CK(clk), .Q(
        new_AGEMA_signal_3741), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2556_s_current_state_reg ( .D(
        new_AGEMA_signal_1382), .CK(clk), .Q(new_AGEMA_signal_3745), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2560_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[39]), .CK(clk), .Q(
        new_AGEMA_signal_3749), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2564_s_current_state_reg ( .D(
        new_AGEMA_signal_1379), .CK(clk), .Q(new_AGEMA_signal_3753), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2568_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[38]), .CK(clk), .Q(
        new_AGEMA_signal_3757), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2572_s_current_state_reg ( .D(
        new_AGEMA_signal_1376), .CK(clk), .Q(new_AGEMA_signal_3761), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2576_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[37]), .CK(clk), .Q(
        new_AGEMA_signal_3765), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2580_s_current_state_reg ( .D(
        new_AGEMA_signal_1373), .CK(clk), .Q(new_AGEMA_signal_3769), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2584_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[36]), .CK(clk), .Q(
        new_AGEMA_signal_3773), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2588_s_current_state_reg ( .D(
        new_AGEMA_signal_1370), .CK(clk), .Q(new_AGEMA_signal_3777), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2592_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[35]), .CK(clk), .Q(
        new_AGEMA_signal_3781), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2596_s_current_state_reg ( .D(
        new_AGEMA_signal_1367), .CK(clk), .Q(new_AGEMA_signal_3785), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2600_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[34]), .CK(clk), .Q(
        new_AGEMA_signal_3789), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2604_s_current_state_reg ( .D(
        new_AGEMA_signal_1364), .CK(clk), .Q(new_AGEMA_signal_3793), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2608_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[33]), .CK(clk), .Q(
        new_AGEMA_signal_3797), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2612_s_current_state_reg ( .D(
        new_AGEMA_signal_1361), .CK(clk), .Q(new_AGEMA_signal_3801), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2616_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[32]), .CK(clk), .Q(
        new_AGEMA_signal_3805), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2620_s_current_state_reg ( .D(
        new_AGEMA_signal_1358), .CK(clk), .Q(new_AGEMA_signal_3809), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2624_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[31]), .CK(clk), .Q(
        new_AGEMA_signal_3813), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2628_s_current_state_reg ( .D(
        new_AGEMA_signal_1355), .CK(clk), .Q(new_AGEMA_signal_3817), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2632_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[30]), .CK(clk), .Q(
        new_AGEMA_signal_3821), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2636_s_current_state_reg ( .D(
        new_AGEMA_signal_1352), .CK(clk), .Q(new_AGEMA_signal_3825), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2640_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[29]), .CK(clk), .Q(
        new_AGEMA_signal_3829), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2644_s_current_state_reg ( .D(
        new_AGEMA_signal_1349), .CK(clk), .Q(new_AGEMA_signal_3833), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2648_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[28]), .CK(clk), .Q(
        new_AGEMA_signal_3837), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2652_s_current_state_reg ( .D(
        new_AGEMA_signal_1346), .CK(clk), .Q(new_AGEMA_signal_3841), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2656_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[27]), .CK(clk), .Q(
        new_AGEMA_signal_3845), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2660_s_current_state_reg ( .D(
        new_AGEMA_signal_1343), .CK(clk), .Q(new_AGEMA_signal_3849), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2664_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[26]), .CK(clk), .Q(
        new_AGEMA_signal_3853), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2668_s_current_state_reg ( .D(
        new_AGEMA_signal_1340), .CK(clk), .Q(new_AGEMA_signal_3857), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2672_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[25]), .CK(clk), .Q(
        new_AGEMA_signal_3861), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2676_s_current_state_reg ( .D(
        new_AGEMA_signal_1337), .CK(clk), .Q(new_AGEMA_signal_3865), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2680_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[24]), .CK(clk), .Q(
        new_AGEMA_signal_3869), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2684_s_current_state_reg ( .D(
        new_AGEMA_signal_1334), .CK(clk), .Q(new_AGEMA_signal_3873), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2688_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[23]), .CK(clk), .Q(
        new_AGEMA_signal_3877), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2692_s_current_state_reg ( .D(
        new_AGEMA_signal_1331), .CK(clk), .Q(new_AGEMA_signal_3881), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2696_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[22]), .CK(clk), .Q(
        new_AGEMA_signal_3885), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2700_s_current_state_reg ( .D(
        new_AGEMA_signal_1328), .CK(clk), .Q(new_AGEMA_signal_3889), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2704_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[21]), .CK(clk), .Q(
        new_AGEMA_signal_3893), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2708_s_current_state_reg ( .D(
        new_AGEMA_signal_1325), .CK(clk), .Q(new_AGEMA_signal_3897), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2712_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[20]), .CK(clk), .Q(
        new_AGEMA_signal_3901), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2716_s_current_state_reg ( .D(
        new_AGEMA_signal_1322), .CK(clk), .Q(new_AGEMA_signal_3905), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2720_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[19]), .CK(clk), .Q(
        new_AGEMA_signal_3909), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2724_s_current_state_reg ( .D(
        new_AGEMA_signal_1319), .CK(clk), .Q(new_AGEMA_signal_3913), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2728_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[18]), .CK(clk), .Q(
        new_AGEMA_signal_3917), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2732_s_current_state_reg ( .D(
        new_AGEMA_signal_1316), .CK(clk), .Q(new_AGEMA_signal_3921), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2736_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[17]), .CK(clk), .Q(
        new_AGEMA_signal_3925), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2740_s_current_state_reg ( .D(
        new_AGEMA_signal_1313), .CK(clk), .Q(new_AGEMA_signal_3929), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2744_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[16]), .CK(clk), .Q(
        new_AGEMA_signal_3933), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2748_s_current_state_reg ( .D(
        new_AGEMA_signal_1310), .CK(clk), .Q(new_AGEMA_signal_3937), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2752_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[15]), .CK(clk), .Q(
        new_AGEMA_signal_3941), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2756_s_current_state_reg ( .D(
        new_AGEMA_signal_1307), .CK(clk), .Q(new_AGEMA_signal_3945), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2760_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[14]), .CK(clk), .Q(
        new_AGEMA_signal_3949), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2764_s_current_state_reg ( .D(
        new_AGEMA_signal_1304), .CK(clk), .Q(new_AGEMA_signal_3953), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2768_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[13]), .CK(clk), .Q(
        new_AGEMA_signal_3957), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2772_s_current_state_reg ( .D(
        new_AGEMA_signal_1301), .CK(clk), .Q(new_AGEMA_signal_3961), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2776_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[12]), .CK(clk), .Q(
        new_AGEMA_signal_3965), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2780_s_current_state_reg ( .D(
        new_AGEMA_signal_1298), .CK(clk), .Q(new_AGEMA_signal_3969), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2784_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[11]), .CK(clk), .Q(
        new_AGEMA_signal_3973), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2788_s_current_state_reg ( .D(
        new_AGEMA_signal_1295), .CK(clk), .Q(new_AGEMA_signal_3977), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2792_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[10]), .CK(clk), .Q(
        new_AGEMA_signal_3981), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2796_s_current_state_reg ( .D(
        new_AGEMA_signal_1292), .CK(clk), .Q(new_AGEMA_signal_3985), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2800_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[9]), .CK(clk), .Q(
        new_AGEMA_signal_3989), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2804_s_current_state_reg ( .D(
        new_AGEMA_signal_1289), .CK(clk), .Q(new_AGEMA_signal_3993), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2808_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[8]), .CK(clk), .Q(
        new_AGEMA_signal_3997), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2812_s_current_state_reg ( .D(
        new_AGEMA_signal_1286), .CK(clk), .Q(new_AGEMA_signal_4001), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2816_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[7]), .CK(clk), .Q(
        new_AGEMA_signal_4005), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2820_s_current_state_reg ( .D(
        new_AGEMA_signal_1283), .CK(clk), .Q(new_AGEMA_signal_4009), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2824_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[6]), .CK(clk), .Q(
        new_AGEMA_signal_4013), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2828_s_current_state_reg ( .D(
        new_AGEMA_signal_1280), .CK(clk), .Q(new_AGEMA_signal_4017), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2832_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[5]), .CK(clk), .Q(
        new_AGEMA_signal_4021), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2836_s_current_state_reg ( .D(
        new_AGEMA_signal_1277), .CK(clk), .Q(new_AGEMA_signal_4025), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2840_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[4]), .CK(clk), .Q(
        new_AGEMA_signal_4029), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2844_s_current_state_reg ( .D(
        new_AGEMA_signal_1274), .CK(clk), .Q(new_AGEMA_signal_4033), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2848_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[3]), .CK(clk), .Q(
        new_AGEMA_signal_4037), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2852_s_current_state_reg ( .D(
        new_AGEMA_signal_1271), .CK(clk), .Q(new_AGEMA_signal_4041), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2856_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[2]), .CK(clk), .Q(
        new_AGEMA_signal_4045), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2860_s_current_state_reg ( .D(
        new_AGEMA_signal_1268), .CK(clk), .Q(new_AGEMA_signal_4049), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2864_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[1]), .CK(clk), .Q(
        new_AGEMA_signal_4053), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2868_s_current_state_reg ( .D(
        new_AGEMA_signal_1265), .CK(clk), .Q(new_AGEMA_signal_4057), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2872_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[0]), .CK(clk), .Q(
        new_AGEMA_signal_4061), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2876_s_current_state_reg ( .D(
        new_AGEMA_signal_1262), .CK(clk), .Q(new_AGEMA_signal_4065), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2880_s_current_state_reg ( .D(FSMSelected[5]), 
        .CK(clk), .Q(new_AGEMA_signal_4069), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2884_s_current_state_reg ( .D(FSMSelected[4]), 
        .CK(clk), .Q(new_AGEMA_signal_4073), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2888_s_current_state_reg ( .D(FSMSelected[3]), 
        .CK(clk), .Q(new_AGEMA_signal_4077), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2892_s_current_state_reg ( .D(FSMSelected[2]), 
        .CK(clk), .Q(new_AGEMA_signal_4081), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2896_s_current_state_reg ( .D(FSMSelected[1]), 
        .CK(clk), .Q(new_AGEMA_signal_4085), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2900_s_current_state_reg ( .D(FSMSelected[0]), 
        .CK(clk), .Q(new_AGEMA_signal_4089), .QN() );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_0_U1 ( .A(MCOutput[2]), .B(
        new_AGEMA_signal_2192), .S(new_AGEMA_signal_2190), .Z(StateRegInput[2]) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1915), .B(
        new_AGEMA_signal_2194), .S(new_AGEMA_signal_2190), .Z(
        new_AGEMA_signal_1922) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_0_U1 ( .A(MCOutput[3]), .B(
        new_AGEMA_signal_2196), .S(new_AGEMA_signal_2190), .Z(StateRegInput[3]) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1975), .B(
        new_AGEMA_signal_2198), .S(new_AGEMA_signal_2190), .Z(
        new_AGEMA_signal_1982) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_0_U1 ( .A(MCOutput[6]), .B(
        new_AGEMA_signal_2200), .S(new_AGEMA_signal_2190), .Z(StateRegInput[6]) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1917), .B(
        new_AGEMA_signal_2202), .S(new_AGEMA_signal_2190), .Z(
        new_AGEMA_signal_1924) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_0_U1 ( .A(MCOutput[7]), .B(
        new_AGEMA_signal_2204), .S(new_AGEMA_signal_2190), .Z(StateRegInput[7]) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1977), .B(
        new_AGEMA_signal_2206), .S(new_AGEMA_signal_2190), .Z(
        new_AGEMA_signal_1984) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_0_U1 ( .A(MCOutput[10]), .B(
        new_AGEMA_signal_2208), .S(n39), .Z(StateRegInput[10]) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1919), .B(
        new_AGEMA_signal_2210), .S(n39), .Z(new_AGEMA_signal_1926) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_0_U1 ( .A(MCOutput[11]), .B(
        new_AGEMA_signal_2212), .S(n39), .Z(StateRegInput[11]) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1979), .B(
        new_AGEMA_signal_2214), .S(n39), .Z(new_AGEMA_signal_1986) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_0_U1 ( .A(MCOutput[14]), .B(
        new_AGEMA_signal_2216), .S(n39), .Z(StateRegInput[14]) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2033), .B(
        new_AGEMA_signal_2218), .S(n39), .Z(new_AGEMA_signal_2042) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_0_U1 ( .A(MCOutput[15]), .B(
        new_AGEMA_signal_2220), .S(n39), .Z(StateRegInput[15]) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2077), .B(
        new_AGEMA_signal_2222), .S(n39), .Z(new_AGEMA_signal_2085) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_0_U1 ( .A(MCOutput[18]), .B(
        new_AGEMA_signal_2224), .S(n39), .Z(StateRegInput[18]) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1909), .B(
        new_AGEMA_signal_2226), .S(n39), .Z(new_AGEMA_signal_1928) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_0_U1 ( .A(MCOutput[19]), .B(
        new_AGEMA_signal_2228), .S(n39), .Z(StateRegInput[19]) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1968), .B(
        new_AGEMA_signal_2230), .S(n39), .Z(new_AGEMA_signal_1988) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_0_U1 ( .A(MCOutput[22]), .B(
        new_AGEMA_signal_2232), .S(n39), .Z(StateRegInput[22]) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1911), .B(
        new_AGEMA_signal_2234), .S(n39), .Z(new_AGEMA_signal_1930) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_0_U1 ( .A(MCOutput[23]), .B(
        new_AGEMA_signal_2236), .S(n38), .Z(StateRegInput[23]) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1970), .B(
        new_AGEMA_signal_2238), .S(n38), .Z(new_AGEMA_signal_1990) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_0_U1 ( .A(MCOutput[26]), .B(
        new_AGEMA_signal_2240), .S(n38), .Z(StateRegInput[26]) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2023), .B(
        new_AGEMA_signal_2242), .S(n38), .Z(new_AGEMA_signal_2048) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_0_U1 ( .A(MCOutput[27]), .B(
        new_AGEMA_signal_2244), .S(n38), .Z(StateRegInput[27]) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2071), .B(
        new_AGEMA_signal_2246), .S(n38), .Z(new_AGEMA_signal_2091) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_0_U1 ( .A(MCOutput[30]), .B(
        new_AGEMA_signal_2248), .S(n38), .Z(StateRegInput[30]) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1913), .B(
        new_AGEMA_signal_2250), .S(n38), .Z(new_AGEMA_signal_1932) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_0_U1 ( .A(MCOutput[31]), .B(
        new_AGEMA_signal_2252), .S(n38), .Z(StateRegInput[31]) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1973), .B(
        new_AGEMA_signal_2254), .S(n38), .Z(new_AGEMA_signal_1992) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_0_U1 ( .A(MCOutput[34]), .B(
        new_AGEMA_signal_2256), .S(n38), .Z(StateRegInput[34]) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1810), .B(
        new_AGEMA_signal_2258), .S(n38), .Z(new_AGEMA_signal_1821) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_0_U1 ( .A(MCOutput[35]), .B(
        new_AGEMA_signal_2260), .S(n38), .Z(StateRegInput[35]) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1854), .B(
        new_AGEMA_signal_2262), .S(n38), .Z(new_AGEMA_signal_1874) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_0_U1 ( .A(MCOutput[38]), .B(
        new_AGEMA_signal_2264), .S(n37), .Z(StateRegInput[38]) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1812), .B(
        new_AGEMA_signal_2266), .S(n37), .Z(new_AGEMA_signal_1823) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_0_U1 ( .A(MCOutput[39]), .B(
        new_AGEMA_signal_2268), .S(n37), .Z(StateRegInput[39]) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1856), .B(
        new_AGEMA_signal_2270), .S(n37), .Z(new_AGEMA_signal_1876) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_0_U1 ( .A(MCOutput[42]), .B(
        new_AGEMA_signal_2272), .S(n37), .Z(StateRegInput[42]) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1814), .B(
        new_AGEMA_signal_2274), .S(n37), .Z(new_AGEMA_signal_1825) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_0_U1 ( .A(MCOutput[43]), .B(
        new_AGEMA_signal_2276), .S(n37), .Z(StateRegInput[43]) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1858), .B(
        new_AGEMA_signal_2278), .S(n37), .Z(new_AGEMA_signal_1878) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_0_U1 ( .A(MCOutput[46]), .B(
        new_AGEMA_signal_2280), .S(n37), .Z(StateRegInput[46]) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1898), .B(
        new_AGEMA_signal_2282), .S(n37), .Z(new_AGEMA_signal_1940) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_0_U1 ( .A(MCOutput[47]), .B(
        new_AGEMA_signal_2284), .S(n37), .Z(StateRegInput[47]) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1958), .B(
        new_AGEMA_signal_2286), .S(n37), .Z(new_AGEMA_signal_2000) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_0_U1 ( .A(MCOutput[50]), .B(
        new_AGEMA_signal_2288), .S(n37), .Z(StateRegInput[50]) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1901), .B(
        new_AGEMA_signal_2290), .S(n37), .Z(new_AGEMA_signal_1942) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_0_U1 ( .A(MCOutput[51]), .B(
        new_AGEMA_signal_2292), .S(new_AGEMA_signal_2190), .Z(
        StateRegInput[51]) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1960), .B(
        new_AGEMA_signal_2294), .S(new_AGEMA_signal_2190), .Z(
        new_AGEMA_signal_2002) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_0_U1 ( .A(MCOutput[54]), .B(
        new_AGEMA_signal_2296), .S(new_AGEMA_signal_2190), .Z(
        StateRegInput[54]) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1903), .B(
        new_AGEMA_signal_2298), .S(new_AGEMA_signal_2190), .Z(
        new_AGEMA_signal_1944) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_0_U1 ( .A(MCOutput[55]), .B(
        new_AGEMA_signal_2300), .S(new_AGEMA_signal_2190), .Z(
        StateRegInput[55]) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1963), .B(
        new_AGEMA_signal_2302), .S(new_AGEMA_signal_2190), .Z(
        new_AGEMA_signal_2004) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_0_U1 ( .A(MCOutput[58]), .B(
        new_AGEMA_signal_2304), .S(new_AGEMA_signal_2190), .Z(
        StateRegInput[58]) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1906), .B(
        new_AGEMA_signal_2306), .S(new_AGEMA_signal_2190), .Z(
        new_AGEMA_signal_1946) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_0_U1 ( .A(MCOutput[59]), .B(
        new_AGEMA_signal_2308), .S(n39), .Z(StateRegInput[59]) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1965), .B(
        new_AGEMA_signal_2310), .S(n39), .Z(new_AGEMA_signal_2006) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_0_U1 ( .A(MCOutput[62]), .B(
        new_AGEMA_signal_2312), .S(n38), .Z(StateRegInput[62]) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2017), .B(
        new_AGEMA_signal_2314), .S(n38), .Z(new_AGEMA_signal_2060) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_0_U1 ( .A(MCOutput[63]), .B(
        new_AGEMA_signal_2316), .S(n37), .Z(StateRegInput[63]) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2067), .B(
        new_AGEMA_signal_2318), .S(n37), .Z(new_AGEMA_signal_2103) );
  INV_X1 SubCellInst_SboxInst_0_U3_U1 ( .A(SubCellInst_SboxInst_0_YY_1_), .ZN(
        ShiftRowsOutput[7]) );
  INV_X1 SubCellInst_SboxInst_0_U2_U1 ( .A(SubCellInst_SboxInst_0_YY_0_), .ZN(
        ShiftRowsOutput[6]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U14 ( .A(Fresh[0]), .B(
        SubCellInst_SboxInst_0_Q1), .Z(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U13 ( .A(Fresh[0]), .B(
        new_AGEMA_signal_1454), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U10 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U8 ( .A(Fresh[0]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U7 ( .A1(new_AGEMA_signal_1454), .A2(
        Ciphertext_s1[2]), .ZN(SubCellInst_SboxInst_0_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_0_Q1), 
        .A2(SubCellInst_SboxInst_0_n3), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n8), .B(
        SubCellInst_SboxInst_0_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1548) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n7), .B(
        SubCellInst_SboxInst_0_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_0_T0) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2320), 
        .B(SubCellInst_SboxInst_0_T0), .Z(SubCellInst_SboxInst_0_Q2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2322), 
        .B(new_AGEMA_signal_1548), .Z(new_AGEMA_signal_1596) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U14 ( .A(Fresh[1]), .B(
        SubCellInst_SboxInst_0_Q4), .Z(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U13 ( .A(Fresh[1]), .B(
        new_AGEMA_signal_1455), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U10 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U8 ( .A(Fresh[1]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U7 ( .A1(new_AGEMA_signal_1455), .A2(
        Ciphertext_s1[2]), .ZN(SubCellInst_SboxInst_0_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_0_Q4), 
        .A2(SubCellInst_SboxInst_0_n3), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n8), .B(
        SubCellInst_SboxInst_0_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1549) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n7), .B(
        SubCellInst_SboxInst_0_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_0_T2) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2324), 
        .B(SubCellInst_SboxInst_0_T2), .Z(SubCellInst_SboxInst_0_Q7) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2326), 
        .B(new_AGEMA_signal_1549), .Z(new_AGEMA_signal_1597) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2328), 
        .B(SubCellInst_SboxInst_0_T0), .Z(SubCellInst_SboxInst_0_L3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2330), 
        .B(new_AGEMA_signal_1548), .Z(new_AGEMA_signal_1598) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L3), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1598), 
        .B(new_AGEMA_signal_1549), .Z(new_AGEMA_signal_1724) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2332), 
        .B(SubCellInst_SboxInst_0_T2), .Z(SubCellInst_SboxInst_0_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2334), 
        .B(new_AGEMA_signal_1549), .Z(new_AGEMA_signal_1660) );
  INV_X1 SubCellInst_SboxInst_1_U3_U1 ( .A(SubCellInst_SboxInst_1_YY_1_), .ZN(
        ShiftRowsOutput[11]) );
  INV_X1 SubCellInst_SboxInst_1_U2_U1 ( .A(SubCellInst_SboxInst_1_YY_0_), .ZN(
        ShiftRowsOutput[10]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U14 ( .A(Fresh[2]), .B(
        SubCellInst_SboxInst_1_Q1), .Z(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U13 ( .A(Fresh[2]), .B(
        new_AGEMA_signal_1460), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U10 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U8 ( .A(Fresh[2]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U7 ( .A1(new_AGEMA_signal_1460), .A2(
        Ciphertext_s1[6]), .ZN(SubCellInst_SboxInst_1_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_1_Q1), 
        .A2(SubCellInst_SboxInst_1_n3), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n8), .B(
        SubCellInst_SboxInst_1_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1551) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n7), .B(
        SubCellInst_SboxInst_1_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_1_T0) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2336), 
        .B(SubCellInst_SboxInst_1_T0), .Z(SubCellInst_SboxInst_1_Q2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2338), 
        .B(new_AGEMA_signal_1551), .Z(new_AGEMA_signal_1600) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U14 ( .A(Fresh[3]), .B(
        SubCellInst_SboxInst_1_Q4), .Z(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U13 ( .A(Fresh[3]), .B(
        new_AGEMA_signal_1461), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U10 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U8 ( .A(Fresh[3]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U7 ( .A1(new_AGEMA_signal_1461), .A2(
        Ciphertext_s1[6]), .ZN(SubCellInst_SboxInst_1_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_1_Q4), 
        .A2(SubCellInst_SboxInst_1_n3), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n8), .B(
        SubCellInst_SboxInst_1_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1552) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n7), .B(
        SubCellInst_SboxInst_1_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_1_T2) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2340), 
        .B(SubCellInst_SboxInst_1_T2), .Z(SubCellInst_SboxInst_1_Q7) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2342), 
        .B(new_AGEMA_signal_1552), .Z(new_AGEMA_signal_1601) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2344), 
        .B(SubCellInst_SboxInst_1_T0), .Z(SubCellInst_SboxInst_1_L3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2346), 
        .B(new_AGEMA_signal_1551), .Z(new_AGEMA_signal_1602) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L3), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1602), 
        .B(new_AGEMA_signal_1552), .Z(new_AGEMA_signal_1726) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2348), 
        .B(SubCellInst_SboxInst_1_T2), .Z(SubCellInst_SboxInst_1_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2350), 
        .B(new_AGEMA_signal_1552), .Z(new_AGEMA_signal_1664) );
  INV_X1 SubCellInst_SboxInst_2_U3_U1 ( .A(SubCellInst_SboxInst_2_YY_1_), .ZN(
        ShiftRowsOutput[15]) );
  INV_X1 SubCellInst_SboxInst_2_U2_U1 ( .A(SubCellInst_SboxInst_2_YY_0_), .ZN(
        ShiftRowsOutput[14]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U14 ( .A(Fresh[4]), .B(
        SubCellInst_SboxInst_2_Q1), .Z(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U13 ( .A(Fresh[4]), .B(
        new_AGEMA_signal_1466), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U10 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U8 ( .A(Fresh[4]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U7 ( .A1(new_AGEMA_signal_1466), .A2(
        Ciphertext_s1[10]), .ZN(SubCellInst_SboxInst_2_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_2_Q1), 
        .A2(SubCellInst_SboxInst_2_n3), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n8), .B(
        SubCellInst_SboxInst_2_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1554) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n7), .B(
        SubCellInst_SboxInst_2_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_2_T0) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2352), 
        .B(SubCellInst_SboxInst_2_T0), .Z(SubCellInst_SboxInst_2_Q2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2354), 
        .B(new_AGEMA_signal_1554), .Z(new_AGEMA_signal_1604) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U14 ( .A(Fresh[5]), .B(
        SubCellInst_SboxInst_2_Q4), .Z(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U13 ( .A(Fresh[5]), .B(
        new_AGEMA_signal_1467), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U10 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U8 ( .A(Fresh[5]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U7 ( .A1(new_AGEMA_signal_1467), .A2(
        Ciphertext_s1[10]), .ZN(SubCellInst_SboxInst_2_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_2_Q4), 
        .A2(SubCellInst_SboxInst_2_n3), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n8), .B(
        SubCellInst_SboxInst_2_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1555) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n7), .B(
        SubCellInst_SboxInst_2_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_2_T2) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2356), 
        .B(SubCellInst_SboxInst_2_T2), .Z(SubCellInst_SboxInst_2_Q7) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2358), 
        .B(new_AGEMA_signal_1555), .Z(new_AGEMA_signal_1605) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2360), 
        .B(SubCellInst_SboxInst_2_T0), .Z(SubCellInst_SboxInst_2_L3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2362), 
        .B(new_AGEMA_signal_1554), .Z(new_AGEMA_signal_1606) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L3), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1606), 
        .B(new_AGEMA_signal_1555), .Z(new_AGEMA_signal_1728) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2364), 
        .B(SubCellInst_SboxInst_2_T2), .Z(SubCellInst_SboxInst_2_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2366), 
        .B(new_AGEMA_signal_1555), .Z(new_AGEMA_signal_1668) );
  INV_X1 SubCellInst_SboxInst_3_U3_U1 ( .A(SubCellInst_SboxInst_3_YY_1_), .ZN(
        ShiftRowsOutput[3]) );
  INV_X1 SubCellInst_SboxInst_3_U2_U1 ( .A(SubCellInst_SboxInst_3_YY_0_), .ZN(
        ShiftRowsOutput[2]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U14 ( .A(Fresh[6]), .B(
        SubCellInst_SboxInst_3_Q1), .Z(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U13 ( .A(Fresh[6]), .B(
        new_AGEMA_signal_1472), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U10 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U8 ( .A(Fresh[6]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U7 ( .A1(new_AGEMA_signal_1472), .A2(
        Ciphertext_s1[14]), .ZN(SubCellInst_SboxInst_3_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_3_Q1), 
        .A2(SubCellInst_SboxInst_3_n3), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n8), .B(
        SubCellInst_SboxInst_3_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1557) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n7), .B(
        SubCellInst_SboxInst_3_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_3_T0) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2368), 
        .B(SubCellInst_SboxInst_3_T0), .Z(SubCellInst_SboxInst_3_Q2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2370), 
        .B(new_AGEMA_signal_1557), .Z(new_AGEMA_signal_1608) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U14 ( .A(Fresh[7]), .B(
        SubCellInst_SboxInst_3_Q4), .Z(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U13 ( .A(Fresh[7]), .B(
        new_AGEMA_signal_1473), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U10 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U8 ( .A(Fresh[7]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U7 ( .A1(new_AGEMA_signal_1473), .A2(
        Ciphertext_s1[14]), .ZN(SubCellInst_SboxInst_3_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_3_Q4), 
        .A2(SubCellInst_SboxInst_3_n3), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n8), .B(
        SubCellInst_SboxInst_3_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1558) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n7), .B(
        SubCellInst_SboxInst_3_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_3_T2) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2372), 
        .B(SubCellInst_SboxInst_3_T2), .Z(SubCellInst_SboxInst_3_Q7) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2374), 
        .B(new_AGEMA_signal_1558), .Z(new_AGEMA_signal_1609) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2376), 
        .B(SubCellInst_SboxInst_3_T0), .Z(SubCellInst_SboxInst_3_L3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2378), 
        .B(new_AGEMA_signal_1557), .Z(new_AGEMA_signal_1610) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L3), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1610), 
        .B(new_AGEMA_signal_1558), .Z(new_AGEMA_signal_1730) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2380), 
        .B(SubCellInst_SboxInst_3_T2), .Z(SubCellInst_SboxInst_3_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2382), 
        .B(new_AGEMA_signal_1558), .Z(new_AGEMA_signal_1672) );
  INV_X1 SubCellInst_SboxInst_4_U3_U1 ( .A(SubCellInst_SboxInst_4_YY_1_), .ZN(
        ShiftRowsOutput[27]) );
  INV_X1 SubCellInst_SboxInst_4_U2_U1 ( .A(SubCellInst_SboxInst_4_YY_0_), .ZN(
        ShiftRowsOutput[26]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U14 ( .A(Fresh[8]), .B(
        SubCellInst_SboxInst_4_Q1), .Z(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U13 ( .A(Fresh[8]), .B(
        new_AGEMA_signal_1478), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U10 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U8 ( .A(Fresh[8]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U7 ( .A1(new_AGEMA_signal_1478), .A2(
        Ciphertext_s1[18]), .ZN(SubCellInst_SboxInst_4_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_4_Q1), 
        .A2(SubCellInst_SboxInst_4_n3), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n8), .B(
        SubCellInst_SboxInst_4_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1560) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n7), .B(
        SubCellInst_SboxInst_4_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_4_T0) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2384), 
        .B(SubCellInst_SboxInst_4_T0), .Z(SubCellInst_SboxInst_4_Q2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2386), 
        .B(new_AGEMA_signal_1560), .Z(new_AGEMA_signal_1612) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U14 ( .A(Fresh[9]), .B(
        SubCellInst_SboxInst_4_Q4), .Z(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U13 ( .A(Fresh[9]), .B(
        new_AGEMA_signal_1479), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U10 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U8 ( .A(Fresh[9]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U7 ( .A1(new_AGEMA_signal_1479), .A2(
        Ciphertext_s1[18]), .ZN(SubCellInst_SboxInst_4_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_4_Q4), 
        .A2(SubCellInst_SboxInst_4_n3), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n8), .B(
        SubCellInst_SboxInst_4_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1561) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n7), .B(
        SubCellInst_SboxInst_4_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_4_T2) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2388), 
        .B(SubCellInst_SboxInst_4_T2), .Z(SubCellInst_SboxInst_4_Q7) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2390), 
        .B(new_AGEMA_signal_1561), .Z(new_AGEMA_signal_1613) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2392), 
        .B(SubCellInst_SboxInst_4_T0), .Z(SubCellInst_SboxInst_4_L3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2394), 
        .B(new_AGEMA_signal_1560), .Z(new_AGEMA_signal_1614) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L3), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1614), 
        .B(new_AGEMA_signal_1561), .Z(new_AGEMA_signal_1732) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2396), 
        .B(SubCellInst_SboxInst_4_T2), .Z(SubCellInst_SboxInst_4_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2398), 
        .B(new_AGEMA_signal_1561), .Z(new_AGEMA_signal_1676) );
  INV_X1 SubCellInst_SboxInst_5_U3_U1 ( .A(SubCellInst_SboxInst_5_YY_1_), .ZN(
        ShiftRowsOutput[31]) );
  INV_X1 SubCellInst_SboxInst_5_U2_U1 ( .A(SubCellInst_SboxInst_5_YY_0_), .ZN(
        ShiftRowsOutput[30]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U14 ( .A(Fresh[10]), .B(
        SubCellInst_SboxInst_5_Q1), .Z(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U13 ( .A(Fresh[10]), .B(
        new_AGEMA_signal_1484), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U10 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U8 ( .A(Fresh[10]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U7 ( .A1(new_AGEMA_signal_1484), .A2(
        Ciphertext_s1[22]), .ZN(SubCellInst_SboxInst_5_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_5_Q1), 
        .A2(SubCellInst_SboxInst_5_n3), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n8), .B(
        SubCellInst_SboxInst_5_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1563) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n7), .B(
        SubCellInst_SboxInst_5_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_5_T0) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2400), 
        .B(SubCellInst_SboxInst_5_T0), .Z(SubCellInst_SboxInst_5_Q2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2402), 
        .B(new_AGEMA_signal_1563), .Z(new_AGEMA_signal_1616) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U14 ( .A(Fresh[11]), .B(
        SubCellInst_SboxInst_5_Q4), .Z(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U13 ( .A(Fresh[11]), .B(
        new_AGEMA_signal_1485), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U10 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U8 ( .A(Fresh[11]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U7 ( .A1(new_AGEMA_signal_1485), .A2(
        Ciphertext_s1[22]), .ZN(SubCellInst_SboxInst_5_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_5_Q4), 
        .A2(SubCellInst_SboxInst_5_n3), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n8), .B(
        SubCellInst_SboxInst_5_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1564) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n7), .B(
        SubCellInst_SboxInst_5_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_5_T2) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2404), 
        .B(SubCellInst_SboxInst_5_T2), .Z(SubCellInst_SboxInst_5_Q7) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2406), 
        .B(new_AGEMA_signal_1564), .Z(new_AGEMA_signal_1617) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2408), 
        .B(SubCellInst_SboxInst_5_T0), .Z(SubCellInst_SboxInst_5_L3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2410), 
        .B(new_AGEMA_signal_1563), .Z(new_AGEMA_signal_1618) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L3), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1618), 
        .B(new_AGEMA_signal_1564), .Z(new_AGEMA_signal_1734) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2412), 
        .B(SubCellInst_SboxInst_5_T2), .Z(SubCellInst_SboxInst_5_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2414), 
        .B(new_AGEMA_signal_1564), .Z(new_AGEMA_signal_1680) );
  INV_X1 SubCellInst_SboxInst_6_U3_U1 ( .A(SubCellInst_SboxInst_6_YY_1_), .ZN(
        ShiftRowsOutput[19]) );
  INV_X1 SubCellInst_SboxInst_6_U2_U1 ( .A(SubCellInst_SboxInst_6_YY_0_), .ZN(
        ShiftRowsOutput[18]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U14 ( .A(Fresh[12]), .B(
        SubCellInst_SboxInst_6_Q1), .Z(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U13 ( .A(Fresh[12]), .B(
        new_AGEMA_signal_1490), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U10 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U8 ( .A(Fresh[12]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U7 ( .A1(new_AGEMA_signal_1490), .A2(
        Ciphertext_s1[26]), .ZN(SubCellInst_SboxInst_6_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_6_Q1), 
        .A2(SubCellInst_SboxInst_6_n3), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n8), .B(
        SubCellInst_SboxInst_6_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1566) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n7), .B(
        SubCellInst_SboxInst_6_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_6_T0) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2416), 
        .B(SubCellInst_SboxInst_6_T0), .Z(SubCellInst_SboxInst_6_Q2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2418), 
        .B(new_AGEMA_signal_1566), .Z(new_AGEMA_signal_1620) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U14 ( .A(Fresh[13]), .B(
        SubCellInst_SboxInst_6_Q4), .Z(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U13 ( .A(Fresh[13]), .B(
        new_AGEMA_signal_1491), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U10 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U8 ( .A(Fresh[13]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U7 ( .A1(new_AGEMA_signal_1491), .A2(
        Ciphertext_s1[26]), .ZN(SubCellInst_SboxInst_6_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_6_Q4), 
        .A2(SubCellInst_SboxInst_6_n3), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n8), .B(
        SubCellInst_SboxInst_6_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1567) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n7), .B(
        SubCellInst_SboxInst_6_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_6_T2) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2420), 
        .B(SubCellInst_SboxInst_6_T2), .Z(SubCellInst_SboxInst_6_Q7) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2422), 
        .B(new_AGEMA_signal_1567), .Z(new_AGEMA_signal_1621) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2424), 
        .B(SubCellInst_SboxInst_6_T0), .Z(SubCellInst_SboxInst_6_L3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2426), 
        .B(new_AGEMA_signal_1566), .Z(new_AGEMA_signal_1622) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L3), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1622), 
        .B(new_AGEMA_signal_1567), .Z(new_AGEMA_signal_1736) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2428), 
        .B(SubCellInst_SboxInst_6_T2), .Z(SubCellInst_SboxInst_6_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2430), 
        .B(new_AGEMA_signal_1567), .Z(new_AGEMA_signal_1684) );
  INV_X1 SubCellInst_SboxInst_7_U3_U1 ( .A(SubCellInst_SboxInst_7_YY_1_), .ZN(
        ShiftRowsOutput[23]) );
  INV_X1 SubCellInst_SboxInst_7_U2_U1 ( .A(SubCellInst_SboxInst_7_YY_0_), .ZN(
        ShiftRowsOutput[22]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U14 ( .A(Fresh[14]), .B(
        SubCellInst_SboxInst_7_Q1), .Z(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U13 ( .A(Fresh[14]), .B(
        new_AGEMA_signal_1496), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U10 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U8 ( .A(Fresh[14]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U7 ( .A1(new_AGEMA_signal_1496), .A2(
        Ciphertext_s1[30]), .ZN(SubCellInst_SboxInst_7_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_7_Q1), 
        .A2(SubCellInst_SboxInst_7_n3), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n8), .B(
        SubCellInst_SboxInst_7_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1569) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n7), .B(
        SubCellInst_SboxInst_7_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_7_T0) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2432), 
        .B(SubCellInst_SboxInst_7_T0), .Z(SubCellInst_SboxInst_7_Q2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2434), 
        .B(new_AGEMA_signal_1569), .Z(new_AGEMA_signal_1624) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U14 ( .A(Fresh[15]), .B(
        SubCellInst_SboxInst_7_Q4), .Z(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U13 ( .A(Fresh[15]), .B(
        new_AGEMA_signal_1497), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U10 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U8 ( .A(Fresh[15]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U7 ( .A1(new_AGEMA_signal_1497), .A2(
        Ciphertext_s1[30]), .ZN(SubCellInst_SboxInst_7_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_7_Q4), 
        .A2(SubCellInst_SboxInst_7_n3), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n8), .B(
        SubCellInst_SboxInst_7_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1570) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n7), .B(
        SubCellInst_SboxInst_7_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_7_T2) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2436), 
        .B(SubCellInst_SboxInst_7_T2), .Z(SubCellInst_SboxInst_7_Q7) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2438), 
        .B(new_AGEMA_signal_1570), .Z(new_AGEMA_signal_1625) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2440), 
        .B(SubCellInst_SboxInst_7_T0), .Z(SubCellInst_SboxInst_7_L3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2442), 
        .B(new_AGEMA_signal_1569), .Z(new_AGEMA_signal_1626) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L3), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1626), 
        .B(new_AGEMA_signal_1570), .Z(new_AGEMA_signal_1738) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2444), 
        .B(SubCellInst_SboxInst_7_T2), .Z(SubCellInst_SboxInst_7_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2446), 
        .B(new_AGEMA_signal_1570), .Z(new_AGEMA_signal_1688) );
  INV_X1 SubCellInst_SboxInst_8_U3_U1 ( .A(SubCellInst_SboxInst_8_YY_1_), .ZN(
        AddRoundConstantOutput[35]) );
  INV_X1 SubCellInst_SboxInst_8_U2_U1 ( .A(SubCellInst_SboxInst_8_YY_0_), .ZN(
        AddRoundConstantOutput[34]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U14 ( .A(Fresh[16]), .B(
        SubCellInst_SboxInst_8_Q1), .Z(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U13 ( .A(Fresh[16]), .B(
        new_AGEMA_signal_1502), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U10 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U8 ( .A(Fresh[16]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U7 ( .A1(new_AGEMA_signal_1502), .A2(
        Ciphertext_s1[34]), .ZN(SubCellInst_SboxInst_8_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_8_Q1), 
        .A2(SubCellInst_SboxInst_8_n3), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n8), .B(
        SubCellInst_SboxInst_8_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1572) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n7), .B(
        SubCellInst_SboxInst_8_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_8_T0) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2448), 
        .B(SubCellInst_SboxInst_8_T0), .Z(SubCellInst_SboxInst_8_Q2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2450), 
        .B(new_AGEMA_signal_1572), .Z(new_AGEMA_signal_1628) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U14 ( .A(Fresh[17]), .B(
        SubCellInst_SboxInst_8_Q4), .Z(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U13 ( .A(Fresh[17]), .B(
        new_AGEMA_signal_1503), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U10 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U8 ( .A(Fresh[17]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U7 ( .A1(new_AGEMA_signal_1503), .A2(
        Ciphertext_s1[34]), .ZN(SubCellInst_SboxInst_8_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_8_Q4), 
        .A2(SubCellInst_SboxInst_8_n3), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n8), .B(
        SubCellInst_SboxInst_8_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1573) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n7), .B(
        SubCellInst_SboxInst_8_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_8_T2) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2452), 
        .B(SubCellInst_SboxInst_8_T2), .Z(SubCellInst_SboxInst_8_Q7) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2454), 
        .B(new_AGEMA_signal_1573), .Z(new_AGEMA_signal_1629) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2456), 
        .B(SubCellInst_SboxInst_8_T0), .Z(SubCellInst_SboxInst_8_L3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2458), 
        .B(new_AGEMA_signal_1572), .Z(new_AGEMA_signal_1630) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L3), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1630), 
        .B(new_AGEMA_signal_1573), .Z(new_AGEMA_signal_1740) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2460), 
        .B(SubCellInst_SboxInst_8_T2), .Z(SubCellInst_SboxInst_8_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2462), 
        .B(new_AGEMA_signal_1573), .Z(new_AGEMA_signal_1692) );
  INV_X1 SubCellInst_SboxInst_9_U3_U1 ( .A(SubCellInst_SboxInst_9_YY_1_), .ZN(
        AddRoundConstantOutput[39]) );
  INV_X1 SubCellInst_SboxInst_9_U2_U1 ( .A(SubCellInst_SboxInst_9_YY_0_), .ZN(
        AddRoundConstantOutput[38]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U14 ( .A(Fresh[18]), .B(
        SubCellInst_SboxInst_9_Q1), .Z(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U13 ( .A(Fresh[18]), .B(
        new_AGEMA_signal_1508), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U10 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U8 ( .A(Fresh[18]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U7 ( .A1(new_AGEMA_signal_1508), .A2(
        Ciphertext_s1[38]), .ZN(SubCellInst_SboxInst_9_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_9_Q1), 
        .A2(SubCellInst_SboxInst_9_n3), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n8), .B(
        SubCellInst_SboxInst_9_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1575) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n7), .B(
        SubCellInst_SboxInst_9_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_9_T0) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2464), 
        .B(SubCellInst_SboxInst_9_T0), .Z(SubCellInst_SboxInst_9_Q2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2466), 
        .B(new_AGEMA_signal_1575), .Z(new_AGEMA_signal_1632) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U14 ( .A(Fresh[19]), .B(
        SubCellInst_SboxInst_9_Q4), .Z(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U13 ( .A(Fresh[19]), .B(
        new_AGEMA_signal_1509), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U10 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U8 ( .A(Fresh[19]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U7 ( .A1(new_AGEMA_signal_1509), .A2(
        Ciphertext_s1[38]), .ZN(SubCellInst_SboxInst_9_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_9_Q4), 
        .A2(SubCellInst_SboxInst_9_n3), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n8), .B(
        SubCellInst_SboxInst_9_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1576) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n7), .B(
        SubCellInst_SboxInst_9_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_9_T2) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2468), 
        .B(SubCellInst_SboxInst_9_T2), .Z(SubCellInst_SboxInst_9_Q7) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2470), 
        .B(new_AGEMA_signal_1576), .Z(new_AGEMA_signal_1633) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2472), 
        .B(SubCellInst_SboxInst_9_T0), .Z(SubCellInst_SboxInst_9_L3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2474), 
        .B(new_AGEMA_signal_1575), .Z(new_AGEMA_signal_1634) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L3), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1634), 
        .B(new_AGEMA_signal_1576), .Z(new_AGEMA_signal_1742) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2476), 
        .B(SubCellInst_SboxInst_9_T2), .Z(SubCellInst_SboxInst_9_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2478), 
        .B(new_AGEMA_signal_1576), .Z(new_AGEMA_signal_1696) );
  INV_X1 SubCellInst_SboxInst_10_U3_U1 ( .A(SubCellInst_SboxInst_10_YY_1_), 
        .ZN(AddRoundConstantOutput[43]) );
  INV_X1 SubCellInst_SboxInst_10_U2_U1 ( .A(SubCellInst_SboxInst_10_YY_0_), 
        .ZN(AddRoundConstantOutput[42]) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U14 ( .A(Fresh[20]), .B(
        SubCellInst_SboxInst_10_Q1), .Z(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U13 ( .A(Fresh[20]), .B(
        new_AGEMA_signal_1514), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U10 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_10_n3), 
        .A2(SubCellInst_SboxInst_10_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U8 ( .A(Fresh[20]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U7 ( .A1(new_AGEMA_signal_1514), 
        .A2(Ciphertext_s1[42]), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_10_Q1), 
        .A2(SubCellInst_SboxInst_10_n3), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n8), .B(
        SubCellInst_SboxInst_10_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1578)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n7), .B(
        SubCellInst_SboxInst_10_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_10_T0) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2480), 
        .B(SubCellInst_SboxInst_10_T0), .Z(SubCellInst_SboxInst_10_Q2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2482), 
        .B(new_AGEMA_signal_1578), .Z(new_AGEMA_signal_1636) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U14 ( .A(Fresh[21]), .B(
        SubCellInst_SboxInst_10_Q4), .Z(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U13 ( .A(Fresh[21]), .B(
        new_AGEMA_signal_1515), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U10 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_10_n3), 
        .A2(SubCellInst_SboxInst_10_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U8 ( .A(Fresh[21]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U7 ( .A1(new_AGEMA_signal_1515), 
        .A2(Ciphertext_s1[42]), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_10_Q4), 
        .A2(SubCellInst_SboxInst_10_n3), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n8), .B(
        SubCellInst_SboxInst_10_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1579)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n7), .B(
        SubCellInst_SboxInst_10_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_10_T2) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2484), 
        .B(SubCellInst_SboxInst_10_T2), .Z(SubCellInst_SboxInst_10_Q7) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2486), 
        .B(new_AGEMA_signal_1579), .Z(new_AGEMA_signal_1637) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2488), .B(SubCellInst_SboxInst_10_T0), .Z(SubCellInst_SboxInst_10_L3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2490), .B(new_AGEMA_signal_1578), .Z(new_AGEMA_signal_1638) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L3), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1638), .B(new_AGEMA_signal_1579), .Z(new_AGEMA_signal_1744) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2492), .B(SubCellInst_SboxInst_10_T2), .Z(SubCellInst_SboxInst_10_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2494), .B(new_AGEMA_signal_1579), .Z(new_AGEMA_signal_1700) );
  INV_X1 SubCellInst_SboxInst_11_U3_U1 ( .A(SubCellInst_SboxInst_11_YY_1_), 
        .ZN(SubCellOutput_47) );
  INV_X1 SubCellInst_SboxInst_11_U2_U1 ( .A(SubCellInst_SboxInst_11_YY_0_), 
        .ZN(SubCellOutput_46) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U14 ( .A(Fresh[22]), .B(
        SubCellInst_SboxInst_11_Q1), .Z(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U13 ( .A(Fresh[22]), .B(
        new_AGEMA_signal_1520), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U10 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_11_n3), 
        .A2(SubCellInst_SboxInst_11_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U8 ( .A(Fresh[22]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U7 ( .A1(new_AGEMA_signal_1520), 
        .A2(Ciphertext_s1[46]), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_11_Q1), 
        .A2(SubCellInst_SboxInst_11_n3), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n8), .B(
        SubCellInst_SboxInst_11_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1581)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n7), .B(
        SubCellInst_SboxInst_11_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_11_T0) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2496), 
        .B(SubCellInst_SboxInst_11_T0), .Z(SubCellInst_SboxInst_11_Q2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2498), 
        .B(new_AGEMA_signal_1581), .Z(new_AGEMA_signal_1640) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U14 ( .A(Fresh[23]), .B(
        SubCellInst_SboxInst_11_Q4), .Z(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U13 ( .A(Fresh[23]), .B(
        new_AGEMA_signal_1521), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U10 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_11_n3), 
        .A2(SubCellInst_SboxInst_11_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U8 ( .A(Fresh[23]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U7 ( .A1(new_AGEMA_signal_1521), 
        .A2(Ciphertext_s1[46]), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_11_Q4), 
        .A2(SubCellInst_SboxInst_11_n3), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n8), .B(
        SubCellInst_SboxInst_11_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1582)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n7), .B(
        SubCellInst_SboxInst_11_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_11_T2) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2500), 
        .B(SubCellInst_SboxInst_11_T2), .Z(SubCellInst_SboxInst_11_Q7) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2502), 
        .B(new_AGEMA_signal_1582), .Z(new_AGEMA_signal_1641) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2504), .B(SubCellInst_SboxInst_11_T0), .Z(SubCellInst_SboxInst_11_L3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2506), .B(new_AGEMA_signal_1581), .Z(new_AGEMA_signal_1642) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L3), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1642), .B(new_AGEMA_signal_1582), .Z(new_AGEMA_signal_1746) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2508), .B(SubCellInst_SboxInst_11_T2), .Z(SubCellInst_SboxInst_11_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2510), .B(new_AGEMA_signal_1582), .Z(new_AGEMA_signal_1704) );
  INV_X1 SubCellInst_SboxInst_12_U3_U1 ( .A(SubCellInst_SboxInst_12_YY_1_), 
        .ZN(AddRoundConstantOutput[51]) );
  INV_X1 SubCellInst_SboxInst_12_U2_U1 ( .A(SubCellInst_SboxInst_12_YY_0_), 
        .ZN(AddRoundConstantOutput[50]) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U14 ( .A(Fresh[24]), .B(
        SubCellInst_SboxInst_12_Q1), .Z(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U13 ( .A(Fresh[24]), .B(
        new_AGEMA_signal_1526), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U10 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_12_n3), 
        .A2(SubCellInst_SboxInst_12_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U8 ( .A(Fresh[24]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U7 ( .A1(new_AGEMA_signal_1526), 
        .A2(Ciphertext_s1[50]), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_12_Q1), 
        .A2(SubCellInst_SboxInst_12_n3), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n8), .B(
        SubCellInst_SboxInst_12_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1584)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n7), .B(
        SubCellInst_SboxInst_12_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_12_T0) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2512), 
        .B(SubCellInst_SboxInst_12_T0), .Z(SubCellInst_SboxInst_12_Q2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2514), 
        .B(new_AGEMA_signal_1584), .Z(new_AGEMA_signal_1644) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U14 ( .A(Fresh[25]), .B(
        SubCellInst_SboxInst_12_Q4), .Z(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U13 ( .A(Fresh[25]), .B(
        new_AGEMA_signal_1527), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U10 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_12_n3), 
        .A2(SubCellInst_SboxInst_12_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U8 ( .A(Fresh[25]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U7 ( .A1(new_AGEMA_signal_1527), 
        .A2(Ciphertext_s1[50]), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_12_Q4), 
        .A2(SubCellInst_SboxInst_12_n3), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n8), .B(
        SubCellInst_SboxInst_12_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1585)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n7), .B(
        SubCellInst_SboxInst_12_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_12_T2) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2516), 
        .B(SubCellInst_SboxInst_12_T2), .Z(SubCellInst_SboxInst_12_Q7) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2518), 
        .B(new_AGEMA_signal_1585), .Z(new_AGEMA_signal_1645) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2520), .B(SubCellInst_SboxInst_12_T0), .Z(SubCellInst_SboxInst_12_L3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2522), .B(new_AGEMA_signal_1584), .Z(new_AGEMA_signal_1646) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L3), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1646), .B(new_AGEMA_signal_1585), .Z(new_AGEMA_signal_1748) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2524), .B(SubCellInst_SboxInst_12_T2), .Z(SubCellInst_SboxInst_12_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2526), .B(new_AGEMA_signal_1585), .Z(new_AGEMA_signal_1708) );
  INV_X1 SubCellInst_SboxInst_13_U3_U1 ( .A(SubCellInst_SboxInst_13_YY_1_), 
        .ZN(AddRoundConstantOutput[55]) );
  INV_X1 SubCellInst_SboxInst_13_U2_U1 ( .A(SubCellInst_SboxInst_13_YY_0_), 
        .ZN(AddRoundConstantOutput[54]) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U14 ( .A(Fresh[26]), .B(
        SubCellInst_SboxInst_13_Q1), .Z(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U13 ( .A(Fresh[26]), .B(
        new_AGEMA_signal_1532), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U10 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_13_n3), 
        .A2(SubCellInst_SboxInst_13_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U8 ( .A(Fresh[26]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U7 ( .A1(new_AGEMA_signal_1532), 
        .A2(Ciphertext_s1[54]), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_13_Q1), 
        .A2(SubCellInst_SboxInst_13_n3), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n8), .B(
        SubCellInst_SboxInst_13_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1587)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n7), .B(
        SubCellInst_SboxInst_13_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_13_T0) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2528), 
        .B(SubCellInst_SboxInst_13_T0), .Z(SubCellInst_SboxInst_13_Q2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2530), 
        .B(new_AGEMA_signal_1587), .Z(new_AGEMA_signal_1648) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U14 ( .A(Fresh[27]), .B(
        SubCellInst_SboxInst_13_Q4), .Z(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U13 ( .A(Fresh[27]), .B(
        new_AGEMA_signal_1533), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U10 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_13_n3), 
        .A2(SubCellInst_SboxInst_13_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U8 ( .A(Fresh[27]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U7 ( .A1(new_AGEMA_signal_1533), 
        .A2(Ciphertext_s1[54]), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_13_Q4), 
        .A2(SubCellInst_SboxInst_13_n3), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n8), .B(
        SubCellInst_SboxInst_13_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1588)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n7), .B(
        SubCellInst_SboxInst_13_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_13_T2) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2532), 
        .B(SubCellInst_SboxInst_13_T2), .Z(SubCellInst_SboxInst_13_Q7) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2534), 
        .B(new_AGEMA_signal_1588), .Z(new_AGEMA_signal_1649) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2536), .B(SubCellInst_SboxInst_13_T0), .Z(SubCellInst_SboxInst_13_L3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2538), .B(new_AGEMA_signal_1587), .Z(new_AGEMA_signal_1650) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L3), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1650), .B(new_AGEMA_signal_1588), .Z(new_AGEMA_signal_1750) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2540), .B(SubCellInst_SboxInst_13_T2), .Z(SubCellInst_SboxInst_13_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2542), .B(new_AGEMA_signal_1588), .Z(new_AGEMA_signal_1712) );
  INV_X1 SubCellInst_SboxInst_14_U3_U1 ( .A(SubCellInst_SboxInst_14_YY_1_), 
        .ZN(AddRoundConstantOutput[59]) );
  INV_X1 SubCellInst_SboxInst_14_U2_U1 ( .A(SubCellInst_SboxInst_14_YY_0_), 
        .ZN(AddRoundConstantOutput[58]) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U14 ( .A(Fresh[28]), .B(
        SubCellInst_SboxInst_14_Q1), .Z(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U13 ( .A(Fresh[28]), .B(
        new_AGEMA_signal_1538), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U10 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_14_n3), 
        .A2(SubCellInst_SboxInst_14_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U8 ( .A(Fresh[28]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U7 ( .A1(new_AGEMA_signal_1538), 
        .A2(Ciphertext_s1[58]), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_14_Q1), 
        .A2(SubCellInst_SboxInst_14_n3), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n8), .B(
        SubCellInst_SboxInst_14_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1590)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n7), .B(
        SubCellInst_SboxInst_14_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_14_T0) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2544), 
        .B(SubCellInst_SboxInst_14_T0), .Z(SubCellInst_SboxInst_14_Q2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2546), 
        .B(new_AGEMA_signal_1590), .Z(new_AGEMA_signal_1652) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U14 ( .A(Fresh[29]), .B(
        SubCellInst_SboxInst_14_Q4), .Z(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U13 ( .A(Fresh[29]), .B(
        new_AGEMA_signal_1539), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U10 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_14_n3), 
        .A2(SubCellInst_SboxInst_14_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U8 ( .A(Fresh[29]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U7 ( .A1(new_AGEMA_signal_1539), 
        .A2(Ciphertext_s1[58]), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_14_Q4), 
        .A2(SubCellInst_SboxInst_14_n3), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n8), .B(
        SubCellInst_SboxInst_14_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1591)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n7), .B(
        SubCellInst_SboxInst_14_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_14_T2) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2548), 
        .B(SubCellInst_SboxInst_14_T2), .Z(SubCellInst_SboxInst_14_Q7) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2550), 
        .B(new_AGEMA_signal_1591), .Z(new_AGEMA_signal_1653) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2552), .B(SubCellInst_SboxInst_14_T0), .Z(SubCellInst_SboxInst_14_L3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2554), .B(new_AGEMA_signal_1590), .Z(new_AGEMA_signal_1654) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L3), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1654), .B(new_AGEMA_signal_1591), .Z(new_AGEMA_signal_1752) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2556), .B(SubCellInst_SboxInst_14_T2), .Z(SubCellInst_SboxInst_14_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2558), .B(new_AGEMA_signal_1591), .Z(new_AGEMA_signal_1716) );
  INV_X1 SubCellInst_SboxInst_15_U3_U1 ( .A(SubCellInst_SboxInst_15_YY_1_), 
        .ZN(SubCellOutput[63]) );
  INV_X1 SubCellInst_SboxInst_15_U2_U1 ( .A(SubCellInst_SboxInst_15_YY_0_), 
        .ZN(SubCellOutput[62]) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U14 ( .A(Fresh[30]), .B(
        SubCellInst_SboxInst_15_Q1), .Z(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U13 ( .A(Fresh[30]), .B(
        new_AGEMA_signal_1544), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U10 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_15_n3), 
        .A2(SubCellInst_SboxInst_15_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U8 ( .A(Fresh[30]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U7 ( .A1(new_AGEMA_signal_1544), 
        .A2(Ciphertext_s1[62]), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_15_Q1), 
        .A2(SubCellInst_SboxInst_15_n3), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n8), .B(
        SubCellInst_SboxInst_15_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1593)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n7), .B(
        SubCellInst_SboxInst_15_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_15_T0) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2560), 
        .B(SubCellInst_SboxInst_15_T0), .Z(SubCellInst_SboxInst_15_Q2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2562), 
        .B(new_AGEMA_signal_1593), .Z(new_AGEMA_signal_1656) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U14 ( .A(Fresh[31]), .B(
        SubCellInst_SboxInst_15_Q4), .Z(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U13 ( .A(Fresh[31]), .B(
        new_AGEMA_signal_1545), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U10 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_15_n3), 
        .A2(SubCellInst_SboxInst_15_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U8 ( .A(Fresh[31]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U7 ( .A1(new_AGEMA_signal_1545), 
        .A2(Ciphertext_s1[62]), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_15_Q4), 
        .A2(SubCellInst_SboxInst_15_n3), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n8), .B(
        SubCellInst_SboxInst_15_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1594)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n7), .B(
        SubCellInst_SboxInst_15_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_15_T2) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2564), 
        .B(SubCellInst_SboxInst_15_T2), .Z(SubCellInst_SboxInst_15_Q7) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2566), 
        .B(new_AGEMA_signal_1594), .Z(new_AGEMA_signal_1657) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2568), .B(SubCellInst_SboxInst_15_T0), .Z(SubCellInst_SboxInst_15_L3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2570), .B(new_AGEMA_signal_1593), .Z(new_AGEMA_signal_1658) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L3), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1658), .B(new_AGEMA_signal_1594), .Z(new_AGEMA_signal_1754) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_2572), .B(SubCellInst_SboxInst_15_T2), .Z(SubCellInst_SboxInst_15_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2574), .B(new_AGEMA_signal_1594), .Z(new_AGEMA_signal_1720) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_2_n1), .B(new_AGEMA_signal_2576), 
        .ZN(AddRoundConstantOutput[62]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1756), .B(1'b0), .Z(new_AGEMA_signal_1800) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[62]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_2_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1720), .Z(new_AGEMA_signal_1756) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_3_n1), .B(new_AGEMA_signal_2578), 
        .ZN(AddRoundConstantOutput[63]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1801), .B(1'b0), .Z(new_AGEMA_signal_1843) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[63]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_3_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1754), .Z(new_AGEMA_signal_1801) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_2_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[46]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1757), .B(1'b0), .Z(new_AGEMA_signal_1802) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_46), .ZN(AddConstXOR_AddConstXOR_XORInst_1_2_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1704), .Z(new_AGEMA_signal_1757) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_3_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[47]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1803), .B(1'b0), .Z(new_AGEMA_signal_1845) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_47), .ZN(AddConstXOR_AddConstXOR_XORInst_1_3_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1746), .Z(new_AGEMA_signal_1803) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_2_n1), .B(new_AGEMA_signal_2580), .ZN(
        ShiftRowsOutput[46]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1758), .B(new_AGEMA_signal_2582), .Z(
        new_AGEMA_signal_1804) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[34]), .ZN(AddRoundTweakeyXOR_XORInst_0_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1692), .Z(new_AGEMA_signal_1758) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_3_n1), .B(new_AGEMA_signal_2584), .ZN(
        ShiftRowsOutput[47]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1805), .B(new_AGEMA_signal_2586), .Z(
        new_AGEMA_signal_1847) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[35]), .ZN(AddRoundTweakeyXOR_XORInst_0_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1740), .Z(new_AGEMA_signal_1805) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_2_n1), .B(new_AGEMA_signal_2588), .ZN(
        ShiftRowsOutput[34]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1759), .B(new_AGEMA_signal_2590), .Z(
        new_AGEMA_signal_1806) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[38]), .ZN(AddRoundTweakeyXOR_XORInst_1_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1696), .Z(new_AGEMA_signal_1759) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_3_n1), .B(new_AGEMA_signal_2592), .ZN(
        ShiftRowsOutput[35]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1807), .B(new_AGEMA_signal_2594), .Z(
        new_AGEMA_signal_1849) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[39]), .ZN(AddRoundTweakeyXOR_XORInst_1_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1742), .Z(new_AGEMA_signal_1807) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_2_n1), .B(new_AGEMA_signal_2596), .ZN(
        ShiftRowsOutput[38]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1760), .B(new_AGEMA_signal_2598), .Z(
        new_AGEMA_signal_1808) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[42]), .ZN(AddRoundTweakeyXOR_XORInst_2_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1700), .Z(new_AGEMA_signal_1760) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_3_n1), .B(new_AGEMA_signal_2600), .ZN(
        ShiftRowsOutput[39]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1809), .B(new_AGEMA_signal_2602), .Z(
        new_AGEMA_signal_1851) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[43]), .ZN(AddRoundTweakeyXOR_XORInst_2_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1744), .Z(new_AGEMA_signal_1809) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_2_n1), .B(new_AGEMA_signal_2604), .ZN(
        ShiftRowsOutput[42]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1852), .B(new_AGEMA_signal_2606), .Z(
        new_AGEMA_signal_1890) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[46]), .ZN(AddRoundTweakeyXOR_XORInst_3_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1802), .Z(new_AGEMA_signal_1852) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_3_n1), .B(new_AGEMA_signal_2608), .ZN(
        ShiftRowsOutput[43]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1891), .B(new_AGEMA_signal_2610), .Z(
        new_AGEMA_signal_1953) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[47]), .ZN(AddRoundTweakeyXOR_XORInst_3_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1845), .Z(new_AGEMA_signal_1891) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_2_n1), .B(new_AGEMA_signal_2612), .ZN(
        MCOutput[34]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1761), .B(new_AGEMA_signal_2614), .Z(
        new_AGEMA_signal_1810) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[50]), .ZN(AddRoundTweakeyXOR_XORInst_4_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1708), .Z(new_AGEMA_signal_1761) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_3_n1), .B(new_AGEMA_signal_2616), .ZN(
        MCOutput[35]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1811), .B(new_AGEMA_signal_2618), .Z(
        new_AGEMA_signal_1854) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[51]), .ZN(AddRoundTweakeyXOR_XORInst_4_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1748), .Z(new_AGEMA_signal_1811) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_2_n1), .B(new_AGEMA_signal_2620), .ZN(
        MCOutput[38]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1762), .B(new_AGEMA_signal_2622), .Z(
        new_AGEMA_signal_1812) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[54]), .ZN(AddRoundTweakeyXOR_XORInst_5_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1712), .Z(new_AGEMA_signal_1762) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_3_n1), .B(new_AGEMA_signal_2624), .ZN(
        MCOutput[39]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1813), .B(new_AGEMA_signal_2626), .Z(
        new_AGEMA_signal_1856) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[55]), .ZN(AddRoundTweakeyXOR_XORInst_5_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1750), .Z(new_AGEMA_signal_1813) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_2_n1), .B(new_AGEMA_signal_2628), .ZN(
        MCOutput[42]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1763), .B(new_AGEMA_signal_2630), .Z(
        new_AGEMA_signal_1814) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[58]), .ZN(AddRoundTweakeyXOR_XORInst_6_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1716), .Z(new_AGEMA_signal_1763) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_3_n1), .B(new_AGEMA_signal_2632), .ZN(
        MCOutput[43]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1815), .B(new_AGEMA_signal_2634), .Z(
        new_AGEMA_signal_1858) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[59]), .ZN(AddRoundTweakeyXOR_XORInst_6_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1752), .Z(new_AGEMA_signal_1815) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_2_n1), .B(new_AGEMA_signal_2636), .ZN(
        MCOutput[46]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1859), .B(new_AGEMA_signal_2638), .Z(
        new_AGEMA_signal_1898) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[62]), .ZN(AddRoundTweakeyXOR_XORInst_7_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1800), .Z(new_AGEMA_signal_1859) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_3_n1), .B(new_AGEMA_signal_2640), .ZN(
        MCOutput[47]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1899), .B(new_AGEMA_signal_2642), .Z(
        new_AGEMA_signal_1958) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[63]), .ZN(AddRoundTweakeyXOR_XORInst_7_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1843), .Z(new_AGEMA_signal_1899) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_2_n2), 
        .B(MCInst_MCR0_XORInst_0_2_n1), .ZN(MCOutput[50]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1861), .B(
        new_AGEMA_signal_1764), .Z(new_AGEMA_signal_1901) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[18]), .B(
        ShiftRowsOutput[2]), .ZN(MCInst_MCR0_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1684), .B(
        new_AGEMA_signal_1672), .Z(new_AGEMA_signal_1764) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[34]), 
        .Z(MCInst_MCR0_XORInst_0_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1810), .Z(new_AGEMA_signal_1861) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_3_n2), 
        .B(MCInst_MCR0_XORInst_0_3_n1), .ZN(MCOutput[51]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1902), .B(
        new_AGEMA_signal_1816), .Z(new_AGEMA_signal_1960) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[19]), .B(
        ShiftRowsOutput[3]), .ZN(MCInst_MCR0_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1736), .B(
        new_AGEMA_signal_1730), .Z(new_AGEMA_signal_1816) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[35]), 
        .Z(MCInst_MCR0_XORInst_0_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1854), .Z(new_AGEMA_signal_1902) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_2_n2), 
        .B(MCInst_MCR0_XORInst_1_2_n1), .ZN(MCOutput[54]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1863), .B(
        new_AGEMA_signal_1765), .Z(new_AGEMA_signal_1903) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[22]), .B(
        ShiftRowsOutput[6]), .ZN(MCInst_MCR0_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1688), .B(
        new_AGEMA_signal_1660), .Z(new_AGEMA_signal_1765) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[38]), 
        .Z(MCInst_MCR0_XORInst_1_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1812), .Z(new_AGEMA_signal_1863) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_3_n2), 
        .B(MCInst_MCR0_XORInst_1_3_n1), .ZN(MCOutput[55]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1904), .B(
        new_AGEMA_signal_1817), .Z(new_AGEMA_signal_1963) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[23]), .B(
        ShiftRowsOutput[7]), .ZN(MCInst_MCR0_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1738), .B(
        new_AGEMA_signal_1724), .Z(new_AGEMA_signal_1817) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[39]), 
        .Z(MCInst_MCR0_XORInst_1_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1856), .Z(new_AGEMA_signal_1904) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_2_n2), 
        .B(MCInst_MCR0_XORInst_2_2_n1), .ZN(MCOutput[58]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1865), .B(
        new_AGEMA_signal_1766), .Z(new_AGEMA_signal_1906) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[26]), .B(
        ShiftRowsOutput[10]), .ZN(MCInst_MCR0_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1676), .B(
        new_AGEMA_signal_1664), .Z(new_AGEMA_signal_1766) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[42]), 
        .Z(MCInst_MCR0_XORInst_2_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1814), .Z(new_AGEMA_signal_1865) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_3_n2), 
        .B(MCInst_MCR0_XORInst_2_3_n1), .ZN(MCOutput[59]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1907), .B(
        new_AGEMA_signal_1818), .Z(new_AGEMA_signal_1965) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[27]), .B(
        ShiftRowsOutput[11]), .ZN(MCInst_MCR0_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1732), .B(
        new_AGEMA_signal_1726), .Z(new_AGEMA_signal_1818) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[43]), 
        .Z(MCInst_MCR0_XORInst_2_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1858), .Z(new_AGEMA_signal_1907) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_2_n2), 
        .B(MCInst_MCR0_XORInst_3_2_n1), .ZN(MCOutput[62]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1966), .B(
        new_AGEMA_signal_1767), .Z(new_AGEMA_signal_2017) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[30]), .B(
        ShiftRowsOutput[14]), .ZN(MCInst_MCR0_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1680), .B(
        new_AGEMA_signal_1668), .Z(new_AGEMA_signal_1767) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[46]), 
        .Z(MCInst_MCR0_XORInst_3_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1898), .Z(new_AGEMA_signal_1966) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_3_n2), 
        .B(MCInst_MCR0_XORInst_3_3_n1), .ZN(MCOutput[63]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2018), .B(
        new_AGEMA_signal_1819), .Z(new_AGEMA_signal_2067) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[31]), .B(
        ShiftRowsOutput[15]), .ZN(MCInst_MCR0_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1734), .B(
        new_AGEMA_signal_1728), .Z(new_AGEMA_signal_1819) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[47]), 
        .Z(MCInst_MCR0_XORInst_3_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2018) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_2_n1), 
        .B(ShiftRowsOutput[18]), .ZN(MCOutput[18]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1867), .B(
        new_AGEMA_signal_1684), .Z(new_AGEMA_signal_1909) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[34]), .ZN(MCInst_MCR2_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1806), .Z(new_AGEMA_signal_1867) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_3_n1), 
        .B(ShiftRowsOutput[19]), .ZN(MCOutput[19]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1910), .B(
        new_AGEMA_signal_1736), .Z(new_AGEMA_signal_1968) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[35]), .ZN(MCInst_MCR2_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1849), .Z(new_AGEMA_signal_1910) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_2_n1), 
        .B(ShiftRowsOutput[22]), .ZN(MCOutput[22]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1868), .B(
        new_AGEMA_signal_1688), .Z(new_AGEMA_signal_1911) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[38]), .ZN(MCInst_MCR2_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1808), .Z(new_AGEMA_signal_1868) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_3_n1), 
        .B(ShiftRowsOutput[23]), .ZN(MCOutput[23]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1912), .B(
        new_AGEMA_signal_1738), .Z(new_AGEMA_signal_1970) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[39]), .ZN(MCInst_MCR2_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1851), .Z(new_AGEMA_signal_1912) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_2_n1), 
        .B(ShiftRowsOutput[26]), .ZN(MCOutput[26]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1971), .B(
        new_AGEMA_signal_1676), .Z(new_AGEMA_signal_2023) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[42]), .ZN(MCInst_MCR2_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1890), .Z(new_AGEMA_signal_1971) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_3_n1), 
        .B(ShiftRowsOutput[27]), .ZN(MCOutput[27]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2024), .B(
        new_AGEMA_signal_1732), .Z(new_AGEMA_signal_2071) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[43]), .ZN(MCInst_MCR2_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1953), .Z(new_AGEMA_signal_2024) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_2_n1), 
        .B(ShiftRowsOutput[30]), .ZN(MCOutput[30]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1869), .B(
        new_AGEMA_signal_1680), .Z(new_AGEMA_signal_1913) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[46]), .ZN(MCInst_MCR2_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1804), .Z(new_AGEMA_signal_1869) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_3_n1), 
        .B(ShiftRowsOutput[31]), .ZN(MCOutput[31]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1914), .B(
        new_AGEMA_signal_1734), .Z(new_AGEMA_signal_1973) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[47]), .ZN(MCInst_MCR2_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1847), .Z(new_AGEMA_signal_1914) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_2_n1), 
        .B(ShiftRowsOutput[18]), .ZN(MCOutput[2]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1870), .B(
        new_AGEMA_signal_1684), .Z(new_AGEMA_signal_1915) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[34]), 
        .ZN(MCInst_MCR3_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1810), .Z(new_AGEMA_signal_1870) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_3_n1), 
        .B(ShiftRowsOutput[19]), .ZN(MCOutput[3]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1916), .B(
        new_AGEMA_signal_1736), .Z(new_AGEMA_signal_1975) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[35]), 
        .ZN(MCInst_MCR3_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1854), .Z(new_AGEMA_signal_1916) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_2_n1), 
        .B(ShiftRowsOutput[22]), .ZN(MCOutput[6]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1871), .B(
        new_AGEMA_signal_1688), .Z(new_AGEMA_signal_1917) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[38]), 
        .ZN(MCInst_MCR3_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1812), .Z(new_AGEMA_signal_1871) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_3_n1), 
        .B(ShiftRowsOutput[23]), .ZN(MCOutput[7]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1918), .B(
        new_AGEMA_signal_1738), .Z(new_AGEMA_signal_1977) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[39]), 
        .ZN(MCInst_MCR3_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1856), .Z(new_AGEMA_signal_1918) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_2_n1), 
        .B(ShiftRowsOutput[26]), .ZN(MCOutput[10]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1872), .B(
        new_AGEMA_signal_1676), .Z(new_AGEMA_signal_1919) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[42]), 
        .ZN(MCInst_MCR3_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1814), .Z(new_AGEMA_signal_1872) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_3_n1), 
        .B(ShiftRowsOutput[27]), .ZN(MCOutput[11]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1920), .B(
        new_AGEMA_signal_1732), .Z(new_AGEMA_signal_1979) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[43]), 
        .ZN(MCInst_MCR3_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1858), .Z(new_AGEMA_signal_1920) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_2_n1), 
        .B(ShiftRowsOutput[30]), .ZN(MCOutput[14]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1980), .B(
        new_AGEMA_signal_1680), .Z(new_AGEMA_signal_2033) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[46]), 
        .ZN(MCInst_MCR3_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1898), .Z(new_AGEMA_signal_1980) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_3_n1), 
        .B(ShiftRowsOutput[31]), .ZN(MCOutput[15]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2034), .B(
        new_AGEMA_signal_1734), .Z(new_AGEMA_signal_2077) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[47]), 
        .ZN(MCInst_MCR3_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2034) );
  DFF_X1 new_AGEMA_reg_buffer_1001_s_current_state_reg ( .D(
        new_AGEMA_signal_2189), .CK(clk), .Q(new_AGEMA_signal_2190), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1003_s_current_state_reg ( .D(
        new_AGEMA_signal_2191), .CK(clk), .Q(new_AGEMA_signal_2192), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1005_s_current_state_reg ( .D(
        new_AGEMA_signal_2193), .CK(clk), .Q(new_AGEMA_signal_2194), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1007_s_current_state_reg ( .D(
        new_AGEMA_signal_2195), .CK(clk), .Q(new_AGEMA_signal_2196), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1009_s_current_state_reg ( .D(
        new_AGEMA_signal_2197), .CK(clk), .Q(new_AGEMA_signal_2198), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1011_s_current_state_reg ( .D(
        new_AGEMA_signal_2199), .CK(clk), .Q(new_AGEMA_signal_2200), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1013_s_current_state_reg ( .D(
        new_AGEMA_signal_2201), .CK(clk), .Q(new_AGEMA_signal_2202), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1015_s_current_state_reg ( .D(
        new_AGEMA_signal_2203), .CK(clk), .Q(new_AGEMA_signal_2204), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1017_s_current_state_reg ( .D(
        new_AGEMA_signal_2205), .CK(clk), .Q(new_AGEMA_signal_2206), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1019_s_current_state_reg ( .D(
        new_AGEMA_signal_2207), .CK(clk), .Q(new_AGEMA_signal_2208), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1021_s_current_state_reg ( .D(
        new_AGEMA_signal_2209), .CK(clk), .Q(new_AGEMA_signal_2210), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1023_s_current_state_reg ( .D(
        new_AGEMA_signal_2211), .CK(clk), .Q(new_AGEMA_signal_2212), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1025_s_current_state_reg ( .D(
        new_AGEMA_signal_2213), .CK(clk), .Q(new_AGEMA_signal_2214), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1027_s_current_state_reg ( .D(
        new_AGEMA_signal_2215), .CK(clk), .Q(new_AGEMA_signal_2216), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1029_s_current_state_reg ( .D(
        new_AGEMA_signal_2217), .CK(clk), .Q(new_AGEMA_signal_2218), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1031_s_current_state_reg ( .D(
        new_AGEMA_signal_2219), .CK(clk), .Q(new_AGEMA_signal_2220), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1033_s_current_state_reg ( .D(
        new_AGEMA_signal_2221), .CK(clk), .Q(new_AGEMA_signal_2222), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1035_s_current_state_reg ( .D(
        new_AGEMA_signal_2223), .CK(clk), .Q(new_AGEMA_signal_2224), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1037_s_current_state_reg ( .D(
        new_AGEMA_signal_2225), .CK(clk), .Q(new_AGEMA_signal_2226), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1039_s_current_state_reg ( .D(
        new_AGEMA_signal_2227), .CK(clk), .Q(new_AGEMA_signal_2228), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1041_s_current_state_reg ( .D(
        new_AGEMA_signal_2229), .CK(clk), .Q(new_AGEMA_signal_2230), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1043_s_current_state_reg ( .D(
        new_AGEMA_signal_2231), .CK(clk), .Q(new_AGEMA_signal_2232), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1045_s_current_state_reg ( .D(
        new_AGEMA_signal_2233), .CK(clk), .Q(new_AGEMA_signal_2234), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1047_s_current_state_reg ( .D(
        new_AGEMA_signal_2235), .CK(clk), .Q(new_AGEMA_signal_2236), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1049_s_current_state_reg ( .D(
        new_AGEMA_signal_2237), .CK(clk), .Q(new_AGEMA_signal_2238), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1051_s_current_state_reg ( .D(
        new_AGEMA_signal_2239), .CK(clk), .Q(new_AGEMA_signal_2240), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1053_s_current_state_reg ( .D(
        new_AGEMA_signal_2241), .CK(clk), .Q(new_AGEMA_signal_2242), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1055_s_current_state_reg ( .D(
        new_AGEMA_signal_2243), .CK(clk), .Q(new_AGEMA_signal_2244), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1057_s_current_state_reg ( .D(
        new_AGEMA_signal_2245), .CK(clk), .Q(new_AGEMA_signal_2246), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1059_s_current_state_reg ( .D(
        new_AGEMA_signal_2247), .CK(clk), .Q(new_AGEMA_signal_2248), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1061_s_current_state_reg ( .D(
        new_AGEMA_signal_2249), .CK(clk), .Q(new_AGEMA_signal_2250), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1063_s_current_state_reg ( .D(
        new_AGEMA_signal_2251), .CK(clk), .Q(new_AGEMA_signal_2252), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1065_s_current_state_reg ( .D(
        new_AGEMA_signal_2253), .CK(clk), .Q(new_AGEMA_signal_2254), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1067_s_current_state_reg ( .D(
        new_AGEMA_signal_2255), .CK(clk), .Q(new_AGEMA_signal_2256), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1069_s_current_state_reg ( .D(
        new_AGEMA_signal_2257), .CK(clk), .Q(new_AGEMA_signal_2258), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1071_s_current_state_reg ( .D(
        new_AGEMA_signal_2259), .CK(clk), .Q(new_AGEMA_signal_2260), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1073_s_current_state_reg ( .D(
        new_AGEMA_signal_2261), .CK(clk), .Q(new_AGEMA_signal_2262), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1075_s_current_state_reg ( .D(
        new_AGEMA_signal_2263), .CK(clk), .Q(new_AGEMA_signal_2264), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1077_s_current_state_reg ( .D(
        new_AGEMA_signal_2265), .CK(clk), .Q(new_AGEMA_signal_2266), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1079_s_current_state_reg ( .D(
        new_AGEMA_signal_2267), .CK(clk), .Q(new_AGEMA_signal_2268), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1081_s_current_state_reg ( .D(
        new_AGEMA_signal_2269), .CK(clk), .Q(new_AGEMA_signal_2270), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1083_s_current_state_reg ( .D(
        new_AGEMA_signal_2271), .CK(clk), .Q(new_AGEMA_signal_2272), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1085_s_current_state_reg ( .D(
        new_AGEMA_signal_2273), .CK(clk), .Q(new_AGEMA_signal_2274), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1087_s_current_state_reg ( .D(
        new_AGEMA_signal_2275), .CK(clk), .Q(new_AGEMA_signal_2276), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1089_s_current_state_reg ( .D(
        new_AGEMA_signal_2277), .CK(clk), .Q(new_AGEMA_signal_2278), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1091_s_current_state_reg ( .D(
        new_AGEMA_signal_2279), .CK(clk), .Q(new_AGEMA_signal_2280), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1093_s_current_state_reg ( .D(
        new_AGEMA_signal_2281), .CK(clk), .Q(new_AGEMA_signal_2282), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1095_s_current_state_reg ( .D(
        new_AGEMA_signal_2283), .CK(clk), .Q(new_AGEMA_signal_2284), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1097_s_current_state_reg ( .D(
        new_AGEMA_signal_2285), .CK(clk), .Q(new_AGEMA_signal_2286), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1099_s_current_state_reg ( .D(
        new_AGEMA_signal_2287), .CK(clk), .Q(new_AGEMA_signal_2288), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1101_s_current_state_reg ( .D(
        new_AGEMA_signal_2289), .CK(clk), .Q(new_AGEMA_signal_2290), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1103_s_current_state_reg ( .D(
        new_AGEMA_signal_2291), .CK(clk), .Q(new_AGEMA_signal_2292), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1105_s_current_state_reg ( .D(
        new_AGEMA_signal_2293), .CK(clk), .Q(new_AGEMA_signal_2294), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1107_s_current_state_reg ( .D(
        new_AGEMA_signal_2295), .CK(clk), .Q(new_AGEMA_signal_2296), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1109_s_current_state_reg ( .D(
        new_AGEMA_signal_2297), .CK(clk), .Q(new_AGEMA_signal_2298), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1111_s_current_state_reg ( .D(
        new_AGEMA_signal_2299), .CK(clk), .Q(new_AGEMA_signal_2300), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1113_s_current_state_reg ( .D(
        new_AGEMA_signal_2301), .CK(clk), .Q(new_AGEMA_signal_2302), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1115_s_current_state_reg ( .D(
        new_AGEMA_signal_2303), .CK(clk), .Q(new_AGEMA_signal_2304), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1117_s_current_state_reg ( .D(
        new_AGEMA_signal_2305), .CK(clk), .Q(new_AGEMA_signal_2306), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1119_s_current_state_reg ( .D(
        new_AGEMA_signal_2307), .CK(clk), .Q(new_AGEMA_signal_2308), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1121_s_current_state_reg ( .D(
        new_AGEMA_signal_2309), .CK(clk), .Q(new_AGEMA_signal_2310), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1123_s_current_state_reg ( .D(
        new_AGEMA_signal_2311), .CK(clk), .Q(new_AGEMA_signal_2312), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1125_s_current_state_reg ( .D(
        new_AGEMA_signal_2313), .CK(clk), .Q(new_AGEMA_signal_2314), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1127_s_current_state_reg ( .D(
        new_AGEMA_signal_2315), .CK(clk), .Q(new_AGEMA_signal_2316), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1129_s_current_state_reg ( .D(
        new_AGEMA_signal_2317), .CK(clk), .Q(new_AGEMA_signal_2318), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1131_s_current_state_reg ( .D(
        new_AGEMA_signal_2319), .CK(clk), .Q(new_AGEMA_signal_2320), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1133_s_current_state_reg ( .D(
        new_AGEMA_signal_2321), .CK(clk), .Q(new_AGEMA_signal_2322), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1135_s_current_state_reg ( .D(
        new_AGEMA_signal_2323), .CK(clk), .Q(new_AGEMA_signal_2324), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1137_s_current_state_reg ( .D(
        new_AGEMA_signal_2325), .CK(clk), .Q(new_AGEMA_signal_2326), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1139_s_current_state_reg ( .D(
        new_AGEMA_signal_2327), .CK(clk), .Q(new_AGEMA_signal_2328), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1141_s_current_state_reg ( .D(
        new_AGEMA_signal_2329), .CK(clk), .Q(new_AGEMA_signal_2330), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1143_s_current_state_reg ( .D(
        new_AGEMA_signal_2331), .CK(clk), .Q(new_AGEMA_signal_2332), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1145_s_current_state_reg ( .D(
        new_AGEMA_signal_2333), .CK(clk), .Q(new_AGEMA_signal_2334), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1147_s_current_state_reg ( .D(
        new_AGEMA_signal_2335), .CK(clk), .Q(new_AGEMA_signal_2336), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1149_s_current_state_reg ( .D(
        new_AGEMA_signal_2337), .CK(clk), .Q(new_AGEMA_signal_2338), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1151_s_current_state_reg ( .D(
        new_AGEMA_signal_2339), .CK(clk), .Q(new_AGEMA_signal_2340), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1153_s_current_state_reg ( .D(
        new_AGEMA_signal_2341), .CK(clk), .Q(new_AGEMA_signal_2342), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1155_s_current_state_reg ( .D(
        new_AGEMA_signal_2343), .CK(clk), .Q(new_AGEMA_signal_2344), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1157_s_current_state_reg ( .D(
        new_AGEMA_signal_2345), .CK(clk), .Q(new_AGEMA_signal_2346), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1159_s_current_state_reg ( .D(
        new_AGEMA_signal_2347), .CK(clk), .Q(new_AGEMA_signal_2348), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1161_s_current_state_reg ( .D(
        new_AGEMA_signal_2349), .CK(clk), .Q(new_AGEMA_signal_2350), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1163_s_current_state_reg ( .D(
        new_AGEMA_signal_2351), .CK(clk), .Q(new_AGEMA_signal_2352), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1165_s_current_state_reg ( .D(
        new_AGEMA_signal_2353), .CK(clk), .Q(new_AGEMA_signal_2354), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1167_s_current_state_reg ( .D(
        new_AGEMA_signal_2355), .CK(clk), .Q(new_AGEMA_signal_2356), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1169_s_current_state_reg ( .D(
        new_AGEMA_signal_2357), .CK(clk), .Q(new_AGEMA_signal_2358), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1171_s_current_state_reg ( .D(
        new_AGEMA_signal_2359), .CK(clk), .Q(new_AGEMA_signal_2360), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1173_s_current_state_reg ( .D(
        new_AGEMA_signal_2361), .CK(clk), .Q(new_AGEMA_signal_2362), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1175_s_current_state_reg ( .D(
        new_AGEMA_signal_2363), .CK(clk), .Q(new_AGEMA_signal_2364), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1177_s_current_state_reg ( .D(
        new_AGEMA_signal_2365), .CK(clk), .Q(new_AGEMA_signal_2366), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1179_s_current_state_reg ( .D(
        new_AGEMA_signal_2367), .CK(clk), .Q(new_AGEMA_signal_2368), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1181_s_current_state_reg ( .D(
        new_AGEMA_signal_2369), .CK(clk), .Q(new_AGEMA_signal_2370), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1183_s_current_state_reg ( .D(
        new_AGEMA_signal_2371), .CK(clk), .Q(new_AGEMA_signal_2372), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1185_s_current_state_reg ( .D(
        new_AGEMA_signal_2373), .CK(clk), .Q(new_AGEMA_signal_2374), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1187_s_current_state_reg ( .D(
        new_AGEMA_signal_2375), .CK(clk), .Q(new_AGEMA_signal_2376), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1189_s_current_state_reg ( .D(
        new_AGEMA_signal_2377), .CK(clk), .Q(new_AGEMA_signal_2378), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1191_s_current_state_reg ( .D(
        new_AGEMA_signal_2379), .CK(clk), .Q(new_AGEMA_signal_2380), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1193_s_current_state_reg ( .D(
        new_AGEMA_signal_2381), .CK(clk), .Q(new_AGEMA_signal_2382), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1195_s_current_state_reg ( .D(
        new_AGEMA_signal_2383), .CK(clk), .Q(new_AGEMA_signal_2384), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1197_s_current_state_reg ( .D(
        new_AGEMA_signal_2385), .CK(clk), .Q(new_AGEMA_signal_2386), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1199_s_current_state_reg ( .D(
        new_AGEMA_signal_2387), .CK(clk), .Q(new_AGEMA_signal_2388), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1201_s_current_state_reg ( .D(
        new_AGEMA_signal_2389), .CK(clk), .Q(new_AGEMA_signal_2390), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1203_s_current_state_reg ( .D(
        new_AGEMA_signal_2391), .CK(clk), .Q(new_AGEMA_signal_2392), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1205_s_current_state_reg ( .D(
        new_AGEMA_signal_2393), .CK(clk), .Q(new_AGEMA_signal_2394), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1207_s_current_state_reg ( .D(
        new_AGEMA_signal_2395), .CK(clk), .Q(new_AGEMA_signal_2396), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1209_s_current_state_reg ( .D(
        new_AGEMA_signal_2397), .CK(clk), .Q(new_AGEMA_signal_2398), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1211_s_current_state_reg ( .D(
        new_AGEMA_signal_2399), .CK(clk), .Q(new_AGEMA_signal_2400), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1213_s_current_state_reg ( .D(
        new_AGEMA_signal_2401), .CK(clk), .Q(new_AGEMA_signal_2402), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1215_s_current_state_reg ( .D(
        new_AGEMA_signal_2403), .CK(clk), .Q(new_AGEMA_signal_2404), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1217_s_current_state_reg ( .D(
        new_AGEMA_signal_2405), .CK(clk), .Q(new_AGEMA_signal_2406), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1219_s_current_state_reg ( .D(
        new_AGEMA_signal_2407), .CK(clk), .Q(new_AGEMA_signal_2408), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1221_s_current_state_reg ( .D(
        new_AGEMA_signal_2409), .CK(clk), .Q(new_AGEMA_signal_2410), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1223_s_current_state_reg ( .D(
        new_AGEMA_signal_2411), .CK(clk), .Q(new_AGEMA_signal_2412), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1225_s_current_state_reg ( .D(
        new_AGEMA_signal_2413), .CK(clk), .Q(new_AGEMA_signal_2414), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1227_s_current_state_reg ( .D(
        new_AGEMA_signal_2415), .CK(clk), .Q(new_AGEMA_signal_2416), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1229_s_current_state_reg ( .D(
        new_AGEMA_signal_2417), .CK(clk), .Q(new_AGEMA_signal_2418), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1231_s_current_state_reg ( .D(
        new_AGEMA_signal_2419), .CK(clk), .Q(new_AGEMA_signal_2420), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1233_s_current_state_reg ( .D(
        new_AGEMA_signal_2421), .CK(clk), .Q(new_AGEMA_signal_2422), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1235_s_current_state_reg ( .D(
        new_AGEMA_signal_2423), .CK(clk), .Q(new_AGEMA_signal_2424), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1237_s_current_state_reg ( .D(
        new_AGEMA_signal_2425), .CK(clk), .Q(new_AGEMA_signal_2426), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1239_s_current_state_reg ( .D(
        new_AGEMA_signal_2427), .CK(clk), .Q(new_AGEMA_signal_2428), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1241_s_current_state_reg ( .D(
        new_AGEMA_signal_2429), .CK(clk), .Q(new_AGEMA_signal_2430), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1243_s_current_state_reg ( .D(
        new_AGEMA_signal_2431), .CK(clk), .Q(new_AGEMA_signal_2432), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1245_s_current_state_reg ( .D(
        new_AGEMA_signal_2433), .CK(clk), .Q(new_AGEMA_signal_2434), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1247_s_current_state_reg ( .D(
        new_AGEMA_signal_2435), .CK(clk), .Q(new_AGEMA_signal_2436), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1249_s_current_state_reg ( .D(
        new_AGEMA_signal_2437), .CK(clk), .Q(new_AGEMA_signal_2438), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1251_s_current_state_reg ( .D(
        new_AGEMA_signal_2439), .CK(clk), .Q(new_AGEMA_signal_2440), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1253_s_current_state_reg ( .D(
        new_AGEMA_signal_2441), .CK(clk), .Q(new_AGEMA_signal_2442), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1255_s_current_state_reg ( .D(
        new_AGEMA_signal_2443), .CK(clk), .Q(new_AGEMA_signal_2444), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1257_s_current_state_reg ( .D(
        new_AGEMA_signal_2445), .CK(clk), .Q(new_AGEMA_signal_2446), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1259_s_current_state_reg ( .D(
        new_AGEMA_signal_2447), .CK(clk), .Q(new_AGEMA_signal_2448), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1261_s_current_state_reg ( .D(
        new_AGEMA_signal_2449), .CK(clk), .Q(new_AGEMA_signal_2450), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1263_s_current_state_reg ( .D(
        new_AGEMA_signal_2451), .CK(clk), .Q(new_AGEMA_signal_2452), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1265_s_current_state_reg ( .D(
        new_AGEMA_signal_2453), .CK(clk), .Q(new_AGEMA_signal_2454), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1267_s_current_state_reg ( .D(
        new_AGEMA_signal_2455), .CK(clk), .Q(new_AGEMA_signal_2456), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1269_s_current_state_reg ( .D(
        new_AGEMA_signal_2457), .CK(clk), .Q(new_AGEMA_signal_2458), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1271_s_current_state_reg ( .D(
        new_AGEMA_signal_2459), .CK(clk), .Q(new_AGEMA_signal_2460), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1273_s_current_state_reg ( .D(
        new_AGEMA_signal_2461), .CK(clk), .Q(new_AGEMA_signal_2462), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1275_s_current_state_reg ( .D(
        new_AGEMA_signal_2463), .CK(clk), .Q(new_AGEMA_signal_2464), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1277_s_current_state_reg ( .D(
        new_AGEMA_signal_2465), .CK(clk), .Q(new_AGEMA_signal_2466), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1279_s_current_state_reg ( .D(
        new_AGEMA_signal_2467), .CK(clk), .Q(new_AGEMA_signal_2468), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1281_s_current_state_reg ( .D(
        new_AGEMA_signal_2469), .CK(clk), .Q(new_AGEMA_signal_2470), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1283_s_current_state_reg ( .D(
        new_AGEMA_signal_2471), .CK(clk), .Q(new_AGEMA_signal_2472), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1285_s_current_state_reg ( .D(
        new_AGEMA_signal_2473), .CK(clk), .Q(new_AGEMA_signal_2474), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1287_s_current_state_reg ( .D(
        new_AGEMA_signal_2475), .CK(clk), .Q(new_AGEMA_signal_2476), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1289_s_current_state_reg ( .D(
        new_AGEMA_signal_2477), .CK(clk), .Q(new_AGEMA_signal_2478), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1291_s_current_state_reg ( .D(
        new_AGEMA_signal_2479), .CK(clk), .Q(new_AGEMA_signal_2480), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1293_s_current_state_reg ( .D(
        new_AGEMA_signal_2481), .CK(clk), .Q(new_AGEMA_signal_2482), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1295_s_current_state_reg ( .D(
        new_AGEMA_signal_2483), .CK(clk), .Q(new_AGEMA_signal_2484), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1297_s_current_state_reg ( .D(
        new_AGEMA_signal_2485), .CK(clk), .Q(new_AGEMA_signal_2486), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1299_s_current_state_reg ( .D(
        new_AGEMA_signal_2487), .CK(clk), .Q(new_AGEMA_signal_2488), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1301_s_current_state_reg ( .D(
        new_AGEMA_signal_2489), .CK(clk), .Q(new_AGEMA_signal_2490), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1303_s_current_state_reg ( .D(
        new_AGEMA_signal_2491), .CK(clk), .Q(new_AGEMA_signal_2492), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1305_s_current_state_reg ( .D(
        new_AGEMA_signal_2493), .CK(clk), .Q(new_AGEMA_signal_2494), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1307_s_current_state_reg ( .D(
        new_AGEMA_signal_2495), .CK(clk), .Q(new_AGEMA_signal_2496), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1309_s_current_state_reg ( .D(
        new_AGEMA_signal_2497), .CK(clk), .Q(new_AGEMA_signal_2498), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1311_s_current_state_reg ( .D(
        new_AGEMA_signal_2499), .CK(clk), .Q(new_AGEMA_signal_2500), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1313_s_current_state_reg ( .D(
        new_AGEMA_signal_2501), .CK(clk), .Q(new_AGEMA_signal_2502), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1315_s_current_state_reg ( .D(
        new_AGEMA_signal_2503), .CK(clk), .Q(new_AGEMA_signal_2504), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1317_s_current_state_reg ( .D(
        new_AGEMA_signal_2505), .CK(clk), .Q(new_AGEMA_signal_2506), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1319_s_current_state_reg ( .D(
        new_AGEMA_signal_2507), .CK(clk), .Q(new_AGEMA_signal_2508), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1321_s_current_state_reg ( .D(
        new_AGEMA_signal_2509), .CK(clk), .Q(new_AGEMA_signal_2510), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1323_s_current_state_reg ( .D(
        new_AGEMA_signal_2511), .CK(clk), .Q(new_AGEMA_signal_2512), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1325_s_current_state_reg ( .D(
        new_AGEMA_signal_2513), .CK(clk), .Q(new_AGEMA_signal_2514), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1327_s_current_state_reg ( .D(
        new_AGEMA_signal_2515), .CK(clk), .Q(new_AGEMA_signal_2516), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1329_s_current_state_reg ( .D(
        new_AGEMA_signal_2517), .CK(clk), .Q(new_AGEMA_signal_2518), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1331_s_current_state_reg ( .D(
        new_AGEMA_signal_2519), .CK(clk), .Q(new_AGEMA_signal_2520), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1333_s_current_state_reg ( .D(
        new_AGEMA_signal_2521), .CK(clk), .Q(new_AGEMA_signal_2522), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1335_s_current_state_reg ( .D(
        new_AGEMA_signal_2523), .CK(clk), .Q(new_AGEMA_signal_2524), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1337_s_current_state_reg ( .D(
        new_AGEMA_signal_2525), .CK(clk), .Q(new_AGEMA_signal_2526), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1339_s_current_state_reg ( .D(
        new_AGEMA_signal_2527), .CK(clk), .Q(new_AGEMA_signal_2528), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1341_s_current_state_reg ( .D(
        new_AGEMA_signal_2529), .CK(clk), .Q(new_AGEMA_signal_2530), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1343_s_current_state_reg ( .D(
        new_AGEMA_signal_2531), .CK(clk), .Q(new_AGEMA_signal_2532), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1345_s_current_state_reg ( .D(
        new_AGEMA_signal_2533), .CK(clk), .Q(new_AGEMA_signal_2534), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1347_s_current_state_reg ( .D(
        new_AGEMA_signal_2535), .CK(clk), .Q(new_AGEMA_signal_2536), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1349_s_current_state_reg ( .D(
        new_AGEMA_signal_2537), .CK(clk), .Q(new_AGEMA_signal_2538), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1351_s_current_state_reg ( .D(
        new_AGEMA_signal_2539), .CK(clk), .Q(new_AGEMA_signal_2540), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1353_s_current_state_reg ( .D(
        new_AGEMA_signal_2541), .CK(clk), .Q(new_AGEMA_signal_2542), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1355_s_current_state_reg ( .D(
        new_AGEMA_signal_2543), .CK(clk), .Q(new_AGEMA_signal_2544), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1357_s_current_state_reg ( .D(
        new_AGEMA_signal_2545), .CK(clk), .Q(new_AGEMA_signal_2546), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1359_s_current_state_reg ( .D(
        new_AGEMA_signal_2547), .CK(clk), .Q(new_AGEMA_signal_2548), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1361_s_current_state_reg ( .D(
        new_AGEMA_signal_2549), .CK(clk), .Q(new_AGEMA_signal_2550), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1363_s_current_state_reg ( .D(
        new_AGEMA_signal_2551), .CK(clk), .Q(new_AGEMA_signal_2552), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1365_s_current_state_reg ( .D(
        new_AGEMA_signal_2553), .CK(clk), .Q(new_AGEMA_signal_2554), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1367_s_current_state_reg ( .D(
        new_AGEMA_signal_2555), .CK(clk), .Q(new_AGEMA_signal_2556), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1369_s_current_state_reg ( .D(
        new_AGEMA_signal_2557), .CK(clk), .Q(new_AGEMA_signal_2558), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1371_s_current_state_reg ( .D(
        new_AGEMA_signal_2559), .CK(clk), .Q(new_AGEMA_signal_2560), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1373_s_current_state_reg ( .D(
        new_AGEMA_signal_2561), .CK(clk), .Q(new_AGEMA_signal_2562), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1375_s_current_state_reg ( .D(
        new_AGEMA_signal_2563), .CK(clk), .Q(new_AGEMA_signal_2564), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1377_s_current_state_reg ( .D(
        new_AGEMA_signal_2565), .CK(clk), .Q(new_AGEMA_signal_2566), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1379_s_current_state_reg ( .D(
        new_AGEMA_signal_2567), .CK(clk), .Q(new_AGEMA_signal_2568), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1381_s_current_state_reg ( .D(
        new_AGEMA_signal_2569), .CK(clk), .Q(new_AGEMA_signal_2570), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1383_s_current_state_reg ( .D(
        new_AGEMA_signal_2571), .CK(clk), .Q(new_AGEMA_signal_2572), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1385_s_current_state_reg ( .D(
        new_AGEMA_signal_2573), .CK(clk), .Q(new_AGEMA_signal_2574), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1387_s_current_state_reg ( .D(
        new_AGEMA_signal_2575), .CK(clk), .Q(new_AGEMA_signal_2576), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1389_s_current_state_reg ( .D(
        new_AGEMA_signal_2577), .CK(clk), .Q(new_AGEMA_signal_2578), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1391_s_current_state_reg ( .D(
        new_AGEMA_signal_2579), .CK(clk), .Q(new_AGEMA_signal_2580), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1393_s_current_state_reg ( .D(
        new_AGEMA_signal_2581), .CK(clk), .Q(new_AGEMA_signal_2582), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1395_s_current_state_reg ( .D(
        new_AGEMA_signal_2583), .CK(clk), .Q(new_AGEMA_signal_2584), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1397_s_current_state_reg ( .D(
        new_AGEMA_signal_2585), .CK(clk), .Q(new_AGEMA_signal_2586), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1399_s_current_state_reg ( .D(
        new_AGEMA_signal_2587), .CK(clk), .Q(new_AGEMA_signal_2588), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1401_s_current_state_reg ( .D(
        new_AGEMA_signal_2589), .CK(clk), .Q(new_AGEMA_signal_2590), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1403_s_current_state_reg ( .D(
        new_AGEMA_signal_2591), .CK(clk), .Q(new_AGEMA_signal_2592), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1405_s_current_state_reg ( .D(
        new_AGEMA_signal_2593), .CK(clk), .Q(new_AGEMA_signal_2594), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1407_s_current_state_reg ( .D(
        new_AGEMA_signal_2595), .CK(clk), .Q(new_AGEMA_signal_2596), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1409_s_current_state_reg ( .D(
        new_AGEMA_signal_2597), .CK(clk), .Q(new_AGEMA_signal_2598), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1411_s_current_state_reg ( .D(
        new_AGEMA_signal_2599), .CK(clk), .Q(new_AGEMA_signal_2600), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1413_s_current_state_reg ( .D(
        new_AGEMA_signal_2601), .CK(clk), .Q(new_AGEMA_signal_2602), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1415_s_current_state_reg ( .D(
        new_AGEMA_signal_2603), .CK(clk), .Q(new_AGEMA_signal_2604), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1417_s_current_state_reg ( .D(
        new_AGEMA_signal_2605), .CK(clk), .Q(new_AGEMA_signal_2606), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1419_s_current_state_reg ( .D(
        new_AGEMA_signal_2607), .CK(clk), .Q(new_AGEMA_signal_2608), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1421_s_current_state_reg ( .D(
        new_AGEMA_signal_2609), .CK(clk), .Q(new_AGEMA_signal_2610), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1423_s_current_state_reg ( .D(
        new_AGEMA_signal_2611), .CK(clk), .Q(new_AGEMA_signal_2612), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1425_s_current_state_reg ( .D(
        new_AGEMA_signal_2613), .CK(clk), .Q(new_AGEMA_signal_2614), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1427_s_current_state_reg ( .D(
        new_AGEMA_signal_2615), .CK(clk), .Q(new_AGEMA_signal_2616), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1429_s_current_state_reg ( .D(
        new_AGEMA_signal_2617), .CK(clk), .Q(new_AGEMA_signal_2618), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1431_s_current_state_reg ( .D(
        new_AGEMA_signal_2619), .CK(clk), .Q(new_AGEMA_signal_2620), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1433_s_current_state_reg ( .D(
        new_AGEMA_signal_2621), .CK(clk), .Q(new_AGEMA_signal_2622), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1435_s_current_state_reg ( .D(
        new_AGEMA_signal_2623), .CK(clk), .Q(new_AGEMA_signal_2624), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1437_s_current_state_reg ( .D(
        new_AGEMA_signal_2625), .CK(clk), .Q(new_AGEMA_signal_2626), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1439_s_current_state_reg ( .D(
        new_AGEMA_signal_2627), .CK(clk), .Q(new_AGEMA_signal_2628), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1441_s_current_state_reg ( .D(
        new_AGEMA_signal_2629), .CK(clk), .Q(new_AGEMA_signal_2630), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1443_s_current_state_reg ( .D(
        new_AGEMA_signal_2631), .CK(clk), .Q(new_AGEMA_signal_2632), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1445_s_current_state_reg ( .D(
        new_AGEMA_signal_2633), .CK(clk), .Q(new_AGEMA_signal_2634), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1447_s_current_state_reg ( .D(
        new_AGEMA_signal_2635), .CK(clk), .Q(new_AGEMA_signal_2636), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1449_s_current_state_reg ( .D(
        new_AGEMA_signal_2637), .CK(clk), .Q(new_AGEMA_signal_2638), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1451_s_current_state_reg ( .D(
        new_AGEMA_signal_2639), .CK(clk), .Q(new_AGEMA_signal_2640), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1453_s_current_state_reg ( .D(
        new_AGEMA_signal_2641), .CK(clk), .Q(new_AGEMA_signal_2642), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1457_s_current_state_reg ( .D(
        new_AGEMA_signal_2645), .CK(clk), .Q(new_AGEMA_signal_2646), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1461_s_current_state_reg ( .D(
        new_AGEMA_signal_2649), .CK(clk), .Q(new_AGEMA_signal_2650), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1465_s_current_state_reg ( .D(
        new_AGEMA_signal_2653), .CK(clk), .Q(new_AGEMA_signal_2654), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1469_s_current_state_reg ( .D(
        new_AGEMA_signal_2657), .CK(clk), .Q(new_AGEMA_signal_2658), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1473_s_current_state_reg ( .D(
        new_AGEMA_signal_2661), .CK(clk), .Q(new_AGEMA_signal_2662), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1477_s_current_state_reg ( .D(
        new_AGEMA_signal_2665), .CK(clk), .Q(new_AGEMA_signal_2666), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1481_s_current_state_reg ( .D(
        new_AGEMA_signal_2669), .CK(clk), .Q(new_AGEMA_signal_2670), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1485_s_current_state_reg ( .D(
        new_AGEMA_signal_2673), .CK(clk), .Q(new_AGEMA_signal_2674), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1489_s_current_state_reg ( .D(
        new_AGEMA_signal_2677), .CK(clk), .Q(new_AGEMA_signal_2678), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1493_s_current_state_reg ( .D(
        new_AGEMA_signal_2681), .CK(clk), .Q(new_AGEMA_signal_2682), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1497_s_current_state_reg ( .D(
        new_AGEMA_signal_2685), .CK(clk), .Q(new_AGEMA_signal_2686), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1501_s_current_state_reg ( .D(
        new_AGEMA_signal_2689), .CK(clk), .Q(new_AGEMA_signal_2690), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1505_s_current_state_reg ( .D(
        new_AGEMA_signal_2693), .CK(clk), .Q(new_AGEMA_signal_2694), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1509_s_current_state_reg ( .D(
        new_AGEMA_signal_2697), .CK(clk), .Q(new_AGEMA_signal_2698), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1513_s_current_state_reg ( .D(
        new_AGEMA_signal_2701), .CK(clk), .Q(new_AGEMA_signal_2702), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1517_s_current_state_reg ( .D(
        new_AGEMA_signal_2705), .CK(clk), .Q(new_AGEMA_signal_2706), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1521_s_current_state_reg ( .D(
        new_AGEMA_signal_2709), .CK(clk), .Q(new_AGEMA_signal_2710), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1525_s_current_state_reg ( .D(
        new_AGEMA_signal_2713), .CK(clk), .Q(new_AGEMA_signal_2714), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1529_s_current_state_reg ( .D(
        new_AGEMA_signal_2717), .CK(clk), .Q(new_AGEMA_signal_2718), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1533_s_current_state_reg ( .D(
        new_AGEMA_signal_2721), .CK(clk), .Q(new_AGEMA_signal_2722), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1537_s_current_state_reg ( .D(
        new_AGEMA_signal_2725), .CK(clk), .Q(new_AGEMA_signal_2726), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1541_s_current_state_reg ( .D(
        new_AGEMA_signal_2729), .CK(clk), .Q(new_AGEMA_signal_2730), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1545_s_current_state_reg ( .D(
        new_AGEMA_signal_2733), .CK(clk), .Q(new_AGEMA_signal_2734), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1549_s_current_state_reg ( .D(
        new_AGEMA_signal_2737), .CK(clk), .Q(new_AGEMA_signal_2738), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1553_s_current_state_reg ( .D(
        new_AGEMA_signal_2741), .CK(clk), .Q(new_AGEMA_signal_2742), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1557_s_current_state_reg ( .D(
        new_AGEMA_signal_2745), .CK(clk), .Q(new_AGEMA_signal_2746), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1561_s_current_state_reg ( .D(
        new_AGEMA_signal_2749), .CK(clk), .Q(new_AGEMA_signal_2750), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1565_s_current_state_reg ( .D(
        new_AGEMA_signal_2753), .CK(clk), .Q(new_AGEMA_signal_2754), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1569_s_current_state_reg ( .D(
        new_AGEMA_signal_2757), .CK(clk), .Q(new_AGEMA_signal_2758), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1573_s_current_state_reg ( .D(
        new_AGEMA_signal_2761), .CK(clk), .Q(new_AGEMA_signal_2762), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1577_s_current_state_reg ( .D(
        new_AGEMA_signal_2765), .CK(clk), .Q(new_AGEMA_signal_2766), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1581_s_current_state_reg ( .D(
        new_AGEMA_signal_2769), .CK(clk), .Q(new_AGEMA_signal_2770), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1585_s_current_state_reg ( .D(
        new_AGEMA_signal_2773), .CK(clk), .Q(new_AGEMA_signal_2774), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1589_s_current_state_reg ( .D(
        new_AGEMA_signal_2777), .CK(clk), .Q(new_AGEMA_signal_2778), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1593_s_current_state_reg ( .D(
        new_AGEMA_signal_2781), .CK(clk), .Q(new_AGEMA_signal_2782), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1597_s_current_state_reg ( .D(
        new_AGEMA_signal_2785), .CK(clk), .Q(new_AGEMA_signal_2786), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1601_s_current_state_reg ( .D(
        new_AGEMA_signal_2789), .CK(clk), .Q(new_AGEMA_signal_2790), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1605_s_current_state_reg ( .D(
        new_AGEMA_signal_2793), .CK(clk), .Q(new_AGEMA_signal_2794), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1609_s_current_state_reg ( .D(
        new_AGEMA_signal_2797), .CK(clk), .Q(new_AGEMA_signal_2798), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1613_s_current_state_reg ( .D(
        new_AGEMA_signal_2801), .CK(clk), .Q(new_AGEMA_signal_2802), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1617_s_current_state_reg ( .D(
        new_AGEMA_signal_2805), .CK(clk), .Q(new_AGEMA_signal_2806), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1621_s_current_state_reg ( .D(
        new_AGEMA_signal_2809), .CK(clk), .Q(new_AGEMA_signal_2810), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1625_s_current_state_reg ( .D(
        new_AGEMA_signal_2813), .CK(clk), .Q(new_AGEMA_signal_2814), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1629_s_current_state_reg ( .D(
        new_AGEMA_signal_2817), .CK(clk), .Q(new_AGEMA_signal_2818), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1633_s_current_state_reg ( .D(
        new_AGEMA_signal_2821), .CK(clk), .Q(new_AGEMA_signal_2822), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1637_s_current_state_reg ( .D(
        new_AGEMA_signal_2825), .CK(clk), .Q(new_AGEMA_signal_2826), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1641_s_current_state_reg ( .D(
        new_AGEMA_signal_2829), .CK(clk), .Q(new_AGEMA_signal_2830), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1645_s_current_state_reg ( .D(
        new_AGEMA_signal_2833), .CK(clk), .Q(new_AGEMA_signal_2834), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1649_s_current_state_reg ( .D(
        new_AGEMA_signal_2837), .CK(clk), .Q(new_AGEMA_signal_2838), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1653_s_current_state_reg ( .D(
        new_AGEMA_signal_2841), .CK(clk), .Q(new_AGEMA_signal_2842), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1657_s_current_state_reg ( .D(
        new_AGEMA_signal_2845), .CK(clk), .Q(new_AGEMA_signal_2846), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1661_s_current_state_reg ( .D(
        new_AGEMA_signal_2849), .CK(clk), .Q(new_AGEMA_signal_2850), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1665_s_current_state_reg ( .D(
        new_AGEMA_signal_2853), .CK(clk), .Q(new_AGEMA_signal_2854), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1669_s_current_state_reg ( .D(
        new_AGEMA_signal_2857), .CK(clk), .Q(new_AGEMA_signal_2858), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1673_s_current_state_reg ( .D(
        new_AGEMA_signal_2861), .CK(clk), .Q(new_AGEMA_signal_2862), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1677_s_current_state_reg ( .D(
        new_AGEMA_signal_2865), .CK(clk), .Q(new_AGEMA_signal_2866), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1681_s_current_state_reg ( .D(
        new_AGEMA_signal_2869), .CK(clk), .Q(new_AGEMA_signal_2870), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1685_s_current_state_reg ( .D(
        new_AGEMA_signal_2873), .CK(clk), .Q(new_AGEMA_signal_2874), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1689_s_current_state_reg ( .D(
        new_AGEMA_signal_2877), .CK(clk), .Q(new_AGEMA_signal_2878), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1693_s_current_state_reg ( .D(
        new_AGEMA_signal_2881), .CK(clk), .Q(new_AGEMA_signal_2882), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1697_s_current_state_reg ( .D(
        new_AGEMA_signal_2885), .CK(clk), .Q(new_AGEMA_signal_2886), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1701_s_current_state_reg ( .D(
        new_AGEMA_signal_2889), .CK(clk), .Q(new_AGEMA_signal_2890), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1705_s_current_state_reg ( .D(
        new_AGEMA_signal_2893), .CK(clk), .Q(new_AGEMA_signal_2894), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1709_s_current_state_reg ( .D(
        new_AGEMA_signal_2897), .CK(clk), .Q(new_AGEMA_signal_2898), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1713_s_current_state_reg ( .D(
        new_AGEMA_signal_2901), .CK(clk), .Q(new_AGEMA_signal_2902), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1715_s_current_state_reg ( .D(
        new_AGEMA_signal_2903), .CK(clk), .Q(new_AGEMA_signal_2904), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1721_s_current_state_reg ( .D(
        new_AGEMA_signal_2909), .CK(clk), .Q(new_AGEMA_signal_2910), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1723_s_current_state_reg ( .D(
        new_AGEMA_signal_2911), .CK(clk), .Q(new_AGEMA_signal_2912), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1725_s_current_state_reg ( .D(
        new_AGEMA_signal_2913), .CK(clk), .Q(new_AGEMA_signal_2914), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1729_s_current_state_reg ( .D(
        new_AGEMA_signal_2917), .CK(clk), .Q(new_AGEMA_signal_2918), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1737_s_current_state_reg ( .D(
        new_AGEMA_signal_2925), .CK(clk), .Q(new_AGEMA_signal_2926), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1739_s_current_state_reg ( .D(
        new_AGEMA_signal_2927), .CK(clk), .Q(new_AGEMA_signal_2928), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1745_s_current_state_reg ( .D(
        new_AGEMA_signal_2933), .CK(clk), .Q(new_AGEMA_signal_2934), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1747_s_current_state_reg ( .D(
        new_AGEMA_signal_2935), .CK(clk), .Q(new_AGEMA_signal_2936), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1749_s_current_state_reg ( .D(
        new_AGEMA_signal_2937), .CK(clk), .Q(new_AGEMA_signal_2938), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1753_s_current_state_reg ( .D(
        new_AGEMA_signal_2941), .CK(clk), .Q(new_AGEMA_signal_2942), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1761_s_current_state_reg ( .D(
        new_AGEMA_signal_2949), .CK(clk), .Q(new_AGEMA_signal_2950), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1763_s_current_state_reg ( .D(
        new_AGEMA_signal_2951), .CK(clk), .Q(new_AGEMA_signal_2952), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1769_s_current_state_reg ( .D(
        new_AGEMA_signal_2957), .CK(clk), .Q(new_AGEMA_signal_2958), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1771_s_current_state_reg ( .D(
        new_AGEMA_signal_2959), .CK(clk), .Q(new_AGEMA_signal_2960), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1773_s_current_state_reg ( .D(
        new_AGEMA_signal_2961), .CK(clk), .Q(new_AGEMA_signal_2962), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1777_s_current_state_reg ( .D(
        new_AGEMA_signal_2965), .CK(clk), .Q(new_AGEMA_signal_2966), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1785_s_current_state_reg ( .D(
        new_AGEMA_signal_2973), .CK(clk), .Q(new_AGEMA_signal_2974), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1787_s_current_state_reg ( .D(
        new_AGEMA_signal_2975), .CK(clk), .Q(new_AGEMA_signal_2976), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1793_s_current_state_reg ( .D(
        new_AGEMA_signal_2981), .CK(clk), .Q(new_AGEMA_signal_2982), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1795_s_current_state_reg ( .D(
        new_AGEMA_signal_2983), .CK(clk), .Q(new_AGEMA_signal_2984), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1797_s_current_state_reg ( .D(
        new_AGEMA_signal_2985), .CK(clk), .Q(new_AGEMA_signal_2986), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1801_s_current_state_reg ( .D(
        new_AGEMA_signal_2989), .CK(clk), .Q(new_AGEMA_signal_2990), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1809_s_current_state_reg ( .D(
        new_AGEMA_signal_2997), .CK(clk), .Q(new_AGEMA_signal_2998), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1811_s_current_state_reg ( .D(
        new_AGEMA_signal_2999), .CK(clk), .Q(new_AGEMA_signal_3000), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1817_s_current_state_reg ( .D(
        new_AGEMA_signal_3005), .CK(clk), .Q(new_AGEMA_signal_3006), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1819_s_current_state_reg ( .D(
        new_AGEMA_signal_3007), .CK(clk), .Q(new_AGEMA_signal_3008), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1821_s_current_state_reg ( .D(
        new_AGEMA_signal_3009), .CK(clk), .Q(new_AGEMA_signal_3010), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1825_s_current_state_reg ( .D(
        new_AGEMA_signal_3013), .CK(clk), .Q(new_AGEMA_signal_3014), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1833_s_current_state_reg ( .D(
        new_AGEMA_signal_3021), .CK(clk), .Q(new_AGEMA_signal_3022), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1835_s_current_state_reg ( .D(
        new_AGEMA_signal_3023), .CK(clk), .Q(new_AGEMA_signal_3024), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1841_s_current_state_reg ( .D(
        new_AGEMA_signal_3029), .CK(clk), .Q(new_AGEMA_signal_3030), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1843_s_current_state_reg ( .D(
        new_AGEMA_signal_3031), .CK(clk), .Q(new_AGEMA_signal_3032), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1845_s_current_state_reg ( .D(
        new_AGEMA_signal_3033), .CK(clk), .Q(new_AGEMA_signal_3034), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1849_s_current_state_reg ( .D(
        new_AGEMA_signal_3037), .CK(clk), .Q(new_AGEMA_signal_3038), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1857_s_current_state_reg ( .D(
        new_AGEMA_signal_3045), .CK(clk), .Q(new_AGEMA_signal_3046), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1859_s_current_state_reg ( .D(
        new_AGEMA_signal_3047), .CK(clk), .Q(new_AGEMA_signal_3048), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1865_s_current_state_reg ( .D(
        new_AGEMA_signal_3053), .CK(clk), .Q(new_AGEMA_signal_3054), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1867_s_current_state_reg ( .D(
        new_AGEMA_signal_3055), .CK(clk), .Q(new_AGEMA_signal_3056), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1869_s_current_state_reg ( .D(
        new_AGEMA_signal_3057), .CK(clk), .Q(new_AGEMA_signal_3058), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1873_s_current_state_reg ( .D(
        new_AGEMA_signal_3061), .CK(clk), .Q(new_AGEMA_signal_3062), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1881_s_current_state_reg ( .D(
        new_AGEMA_signal_3069), .CK(clk), .Q(new_AGEMA_signal_3070), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1883_s_current_state_reg ( .D(
        new_AGEMA_signal_3071), .CK(clk), .Q(new_AGEMA_signal_3072), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1889_s_current_state_reg ( .D(
        new_AGEMA_signal_3077), .CK(clk), .Q(new_AGEMA_signal_3078), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1891_s_current_state_reg ( .D(
        new_AGEMA_signal_3079), .CK(clk), .Q(new_AGEMA_signal_3080), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1893_s_current_state_reg ( .D(
        new_AGEMA_signal_3081), .CK(clk), .Q(new_AGEMA_signal_3082), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1897_s_current_state_reg ( .D(
        new_AGEMA_signal_3085), .CK(clk), .Q(new_AGEMA_signal_3086), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1905_s_current_state_reg ( .D(
        new_AGEMA_signal_3093), .CK(clk), .Q(new_AGEMA_signal_3094), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1907_s_current_state_reg ( .D(
        new_AGEMA_signal_3095), .CK(clk), .Q(new_AGEMA_signal_3096), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1913_s_current_state_reg ( .D(
        new_AGEMA_signal_3101), .CK(clk), .Q(new_AGEMA_signal_3102), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1915_s_current_state_reg ( .D(
        new_AGEMA_signal_3103), .CK(clk), .Q(new_AGEMA_signal_3104), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1917_s_current_state_reg ( .D(
        new_AGEMA_signal_3105), .CK(clk), .Q(new_AGEMA_signal_3106), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1921_s_current_state_reg ( .D(
        new_AGEMA_signal_3109), .CK(clk), .Q(new_AGEMA_signal_3110), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1929_s_current_state_reg ( .D(
        new_AGEMA_signal_3117), .CK(clk), .Q(new_AGEMA_signal_3118), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1931_s_current_state_reg ( .D(
        new_AGEMA_signal_3119), .CK(clk), .Q(new_AGEMA_signal_3120), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1937_s_current_state_reg ( .D(
        new_AGEMA_signal_3125), .CK(clk), .Q(new_AGEMA_signal_3126), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1939_s_current_state_reg ( .D(
        new_AGEMA_signal_3127), .CK(clk), .Q(new_AGEMA_signal_3128), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1941_s_current_state_reg ( .D(
        new_AGEMA_signal_3129), .CK(clk), .Q(new_AGEMA_signal_3130), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1945_s_current_state_reg ( .D(
        new_AGEMA_signal_3133), .CK(clk), .Q(new_AGEMA_signal_3134), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1953_s_current_state_reg ( .D(
        new_AGEMA_signal_3141), .CK(clk), .Q(new_AGEMA_signal_3142), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1955_s_current_state_reg ( .D(
        new_AGEMA_signal_3143), .CK(clk), .Q(new_AGEMA_signal_3144), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1961_s_current_state_reg ( .D(
        new_AGEMA_signal_3149), .CK(clk), .Q(new_AGEMA_signal_3150), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1963_s_current_state_reg ( .D(
        new_AGEMA_signal_3151), .CK(clk), .Q(new_AGEMA_signal_3152), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1965_s_current_state_reg ( .D(
        new_AGEMA_signal_3153), .CK(clk), .Q(new_AGEMA_signal_3154), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1969_s_current_state_reg ( .D(
        new_AGEMA_signal_3157), .CK(clk), .Q(new_AGEMA_signal_3158), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1977_s_current_state_reg ( .D(
        new_AGEMA_signal_3165), .CK(clk), .Q(new_AGEMA_signal_3166), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1979_s_current_state_reg ( .D(
        new_AGEMA_signal_3167), .CK(clk), .Q(new_AGEMA_signal_3168), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1985_s_current_state_reg ( .D(
        new_AGEMA_signal_3173), .CK(clk), .Q(new_AGEMA_signal_3174), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1987_s_current_state_reg ( .D(
        new_AGEMA_signal_3175), .CK(clk), .Q(new_AGEMA_signal_3176), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1989_s_current_state_reg ( .D(
        new_AGEMA_signal_3177), .CK(clk), .Q(new_AGEMA_signal_3178), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1993_s_current_state_reg ( .D(
        new_AGEMA_signal_3181), .CK(clk), .Q(new_AGEMA_signal_3182), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2001_s_current_state_reg ( .D(
        new_AGEMA_signal_3189), .CK(clk), .Q(new_AGEMA_signal_3190), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2003_s_current_state_reg ( .D(
        new_AGEMA_signal_3191), .CK(clk), .Q(new_AGEMA_signal_3192), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2009_s_current_state_reg ( .D(
        new_AGEMA_signal_3197), .CK(clk), .Q(new_AGEMA_signal_3198), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2011_s_current_state_reg ( .D(
        new_AGEMA_signal_3199), .CK(clk), .Q(new_AGEMA_signal_3200), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2013_s_current_state_reg ( .D(
        new_AGEMA_signal_3201), .CK(clk), .Q(new_AGEMA_signal_3202), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2017_s_current_state_reg ( .D(
        new_AGEMA_signal_3205), .CK(clk), .Q(new_AGEMA_signal_3206), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2025_s_current_state_reg ( .D(
        new_AGEMA_signal_3213), .CK(clk), .Q(new_AGEMA_signal_3214), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2027_s_current_state_reg ( .D(
        new_AGEMA_signal_3215), .CK(clk), .Q(new_AGEMA_signal_3216), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2033_s_current_state_reg ( .D(
        new_AGEMA_signal_3221), .CK(clk), .Q(new_AGEMA_signal_3222), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2035_s_current_state_reg ( .D(
        new_AGEMA_signal_3223), .CK(clk), .Q(new_AGEMA_signal_3224), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2037_s_current_state_reg ( .D(
        new_AGEMA_signal_3225), .CK(clk), .Q(new_AGEMA_signal_3226), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2041_s_current_state_reg ( .D(
        new_AGEMA_signal_3229), .CK(clk), .Q(new_AGEMA_signal_3230), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2049_s_current_state_reg ( .D(
        new_AGEMA_signal_3237), .CK(clk), .Q(new_AGEMA_signal_3238), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2051_s_current_state_reg ( .D(
        new_AGEMA_signal_3239), .CK(clk), .Q(new_AGEMA_signal_3240), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2057_s_current_state_reg ( .D(
        new_AGEMA_signal_3245), .CK(clk), .Q(new_AGEMA_signal_3246), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2059_s_current_state_reg ( .D(
        new_AGEMA_signal_3247), .CK(clk), .Q(new_AGEMA_signal_3248), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2061_s_current_state_reg ( .D(
        new_AGEMA_signal_3249), .CK(clk), .Q(new_AGEMA_signal_3250), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2065_s_current_state_reg ( .D(
        new_AGEMA_signal_3253), .CK(clk), .Q(new_AGEMA_signal_3254), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2073_s_current_state_reg ( .D(
        new_AGEMA_signal_3261), .CK(clk), .Q(new_AGEMA_signal_3262), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2075_s_current_state_reg ( .D(
        new_AGEMA_signal_3263), .CK(clk), .Q(new_AGEMA_signal_3264), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2081_s_current_state_reg ( .D(
        new_AGEMA_signal_3269), .CK(clk), .Q(new_AGEMA_signal_3270), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2083_s_current_state_reg ( .D(
        new_AGEMA_signal_3271), .CK(clk), .Q(new_AGEMA_signal_3272), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2085_s_current_state_reg ( .D(
        new_AGEMA_signal_3273), .CK(clk), .Q(new_AGEMA_signal_3274), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2089_s_current_state_reg ( .D(
        new_AGEMA_signal_3277), .CK(clk), .Q(new_AGEMA_signal_3278), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2097_s_current_state_reg ( .D(
        new_AGEMA_signal_3285), .CK(clk), .Q(new_AGEMA_signal_3286), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2101_s_current_state_reg ( .D(
        new_AGEMA_signal_3289), .CK(clk), .Q(new_AGEMA_signal_3290), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2105_s_current_state_reg ( .D(
        new_AGEMA_signal_3293), .CK(clk), .Q(new_AGEMA_signal_3294), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2109_s_current_state_reg ( .D(
        new_AGEMA_signal_3297), .CK(clk), .Q(new_AGEMA_signal_3298), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2113_s_current_state_reg ( .D(
        new_AGEMA_signal_3301), .CK(clk), .Q(new_AGEMA_signal_3302), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2117_s_current_state_reg ( .D(
        new_AGEMA_signal_3305), .CK(clk), .Q(new_AGEMA_signal_3306), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2121_s_current_state_reg ( .D(
        new_AGEMA_signal_3309), .CK(clk), .Q(new_AGEMA_signal_3310), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2125_s_current_state_reg ( .D(
        new_AGEMA_signal_3313), .CK(clk), .Q(new_AGEMA_signal_3314), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2129_s_current_state_reg ( .D(
        new_AGEMA_signal_3317), .CK(clk), .Q(new_AGEMA_signal_3318), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2133_s_current_state_reg ( .D(
        new_AGEMA_signal_3321), .CK(clk), .Q(new_AGEMA_signal_3322), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2137_s_current_state_reg ( .D(
        new_AGEMA_signal_3325), .CK(clk), .Q(new_AGEMA_signal_3326), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2141_s_current_state_reg ( .D(
        new_AGEMA_signal_3329), .CK(clk), .Q(new_AGEMA_signal_3330), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2145_s_current_state_reg ( .D(
        new_AGEMA_signal_3333), .CK(clk), .Q(new_AGEMA_signal_3334), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2149_s_current_state_reg ( .D(
        new_AGEMA_signal_3337), .CK(clk), .Q(new_AGEMA_signal_3338), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2153_s_current_state_reg ( .D(
        new_AGEMA_signal_3341), .CK(clk), .Q(new_AGEMA_signal_3342), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2157_s_current_state_reg ( .D(
        new_AGEMA_signal_3345), .CK(clk), .Q(new_AGEMA_signal_3346), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2161_s_current_state_reg ( .D(
        new_AGEMA_signal_3349), .CK(clk), .Q(new_AGEMA_signal_3350), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2165_s_current_state_reg ( .D(
        new_AGEMA_signal_3353), .CK(clk), .Q(new_AGEMA_signal_3354), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2169_s_current_state_reg ( .D(
        new_AGEMA_signal_3357), .CK(clk), .Q(new_AGEMA_signal_3358), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2173_s_current_state_reg ( .D(
        new_AGEMA_signal_3361), .CK(clk), .Q(new_AGEMA_signal_3362), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2177_s_current_state_reg ( .D(
        new_AGEMA_signal_3365), .CK(clk), .Q(new_AGEMA_signal_3366), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2181_s_current_state_reg ( .D(
        new_AGEMA_signal_3369), .CK(clk), .Q(new_AGEMA_signal_3370), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2185_s_current_state_reg ( .D(
        new_AGEMA_signal_3373), .CK(clk), .Q(new_AGEMA_signal_3374), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2189_s_current_state_reg ( .D(
        new_AGEMA_signal_3377), .CK(clk), .Q(new_AGEMA_signal_3378), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2193_s_current_state_reg ( .D(
        new_AGEMA_signal_3381), .CK(clk), .Q(new_AGEMA_signal_3382), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2197_s_current_state_reg ( .D(
        new_AGEMA_signal_3385), .CK(clk), .Q(new_AGEMA_signal_3386), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2201_s_current_state_reg ( .D(
        new_AGEMA_signal_3389), .CK(clk), .Q(new_AGEMA_signal_3390), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2205_s_current_state_reg ( .D(
        new_AGEMA_signal_3393), .CK(clk), .Q(new_AGEMA_signal_3394), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2209_s_current_state_reg ( .D(
        new_AGEMA_signal_3397), .CK(clk), .Q(new_AGEMA_signal_3398), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2213_s_current_state_reg ( .D(
        new_AGEMA_signal_3401), .CK(clk), .Q(new_AGEMA_signal_3402), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2217_s_current_state_reg ( .D(
        new_AGEMA_signal_3405), .CK(clk), .Q(new_AGEMA_signal_3406), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2221_s_current_state_reg ( .D(
        new_AGEMA_signal_3409), .CK(clk), .Q(new_AGEMA_signal_3410), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2225_s_current_state_reg ( .D(
        new_AGEMA_signal_3413), .CK(clk), .Q(new_AGEMA_signal_3414), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2229_s_current_state_reg ( .D(
        new_AGEMA_signal_3417), .CK(clk), .Q(new_AGEMA_signal_3418), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2233_s_current_state_reg ( .D(
        new_AGEMA_signal_3421), .CK(clk), .Q(new_AGEMA_signal_3422), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2237_s_current_state_reg ( .D(
        new_AGEMA_signal_3425), .CK(clk), .Q(new_AGEMA_signal_3426), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2369_s_current_state_reg ( .D(
        new_AGEMA_signal_3557), .CK(clk), .Q(new_AGEMA_signal_3558), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2373_s_current_state_reg ( .D(
        new_AGEMA_signal_3561), .CK(clk), .Q(new_AGEMA_signal_3562), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2377_s_current_state_reg ( .D(
        new_AGEMA_signal_3565), .CK(clk), .Q(new_AGEMA_signal_3566), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2381_s_current_state_reg ( .D(
        new_AGEMA_signal_3569), .CK(clk), .Q(new_AGEMA_signal_3570), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2385_s_current_state_reg ( .D(
        new_AGEMA_signal_3573), .CK(clk), .Q(new_AGEMA_signal_3574), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2389_s_current_state_reg ( .D(
        new_AGEMA_signal_3577), .CK(clk), .Q(new_AGEMA_signal_3578), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2393_s_current_state_reg ( .D(
        new_AGEMA_signal_3581), .CK(clk), .Q(new_AGEMA_signal_3582), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2397_s_current_state_reg ( .D(
        new_AGEMA_signal_3585), .CK(clk), .Q(new_AGEMA_signal_3586), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2401_s_current_state_reg ( .D(
        new_AGEMA_signal_3589), .CK(clk), .Q(new_AGEMA_signal_3590), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2405_s_current_state_reg ( .D(
        new_AGEMA_signal_3593), .CK(clk), .Q(new_AGEMA_signal_3594), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2409_s_current_state_reg ( .D(
        new_AGEMA_signal_3597), .CK(clk), .Q(new_AGEMA_signal_3598), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2413_s_current_state_reg ( .D(
        new_AGEMA_signal_3601), .CK(clk), .Q(new_AGEMA_signal_3602), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2417_s_current_state_reg ( .D(
        new_AGEMA_signal_3605), .CK(clk), .Q(new_AGEMA_signal_3606), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2421_s_current_state_reg ( .D(
        new_AGEMA_signal_3609), .CK(clk), .Q(new_AGEMA_signal_3610), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2425_s_current_state_reg ( .D(
        new_AGEMA_signal_3613), .CK(clk), .Q(new_AGEMA_signal_3614), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2429_s_current_state_reg ( .D(
        new_AGEMA_signal_3617), .CK(clk), .Q(new_AGEMA_signal_3618), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2433_s_current_state_reg ( .D(
        new_AGEMA_signal_3621), .CK(clk), .Q(new_AGEMA_signal_3622), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2437_s_current_state_reg ( .D(
        new_AGEMA_signal_3625), .CK(clk), .Q(new_AGEMA_signal_3626), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2441_s_current_state_reg ( .D(
        new_AGEMA_signal_3629), .CK(clk), .Q(new_AGEMA_signal_3630), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2445_s_current_state_reg ( .D(
        new_AGEMA_signal_3633), .CK(clk), .Q(new_AGEMA_signal_3634), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2449_s_current_state_reg ( .D(
        new_AGEMA_signal_3637), .CK(clk), .Q(new_AGEMA_signal_3638), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2453_s_current_state_reg ( .D(
        new_AGEMA_signal_3641), .CK(clk), .Q(new_AGEMA_signal_3642), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2457_s_current_state_reg ( .D(
        new_AGEMA_signal_3645), .CK(clk), .Q(new_AGEMA_signal_3646), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2461_s_current_state_reg ( .D(
        new_AGEMA_signal_3649), .CK(clk), .Q(new_AGEMA_signal_3650), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2465_s_current_state_reg ( .D(
        new_AGEMA_signal_3653), .CK(clk), .Q(new_AGEMA_signal_3654), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2469_s_current_state_reg ( .D(
        new_AGEMA_signal_3657), .CK(clk), .Q(new_AGEMA_signal_3658), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2473_s_current_state_reg ( .D(
        new_AGEMA_signal_3661), .CK(clk), .Q(new_AGEMA_signal_3662), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2477_s_current_state_reg ( .D(
        new_AGEMA_signal_3665), .CK(clk), .Q(new_AGEMA_signal_3666), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2481_s_current_state_reg ( .D(
        new_AGEMA_signal_3669), .CK(clk), .Q(new_AGEMA_signal_3670), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2485_s_current_state_reg ( .D(
        new_AGEMA_signal_3673), .CK(clk), .Q(new_AGEMA_signal_3674), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2489_s_current_state_reg ( .D(
        new_AGEMA_signal_3677), .CK(clk), .Q(new_AGEMA_signal_3678), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2493_s_current_state_reg ( .D(
        new_AGEMA_signal_3681), .CK(clk), .Q(new_AGEMA_signal_3682), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2497_s_current_state_reg ( .D(
        new_AGEMA_signal_3685), .CK(clk), .Q(new_AGEMA_signal_3686), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2501_s_current_state_reg ( .D(
        new_AGEMA_signal_3689), .CK(clk), .Q(new_AGEMA_signal_3690), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2505_s_current_state_reg ( .D(
        new_AGEMA_signal_3693), .CK(clk), .Q(new_AGEMA_signal_3694), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2509_s_current_state_reg ( .D(
        new_AGEMA_signal_3697), .CK(clk), .Q(new_AGEMA_signal_3698), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2513_s_current_state_reg ( .D(
        new_AGEMA_signal_3701), .CK(clk), .Q(new_AGEMA_signal_3702), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2517_s_current_state_reg ( .D(
        new_AGEMA_signal_3705), .CK(clk), .Q(new_AGEMA_signal_3706), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2521_s_current_state_reg ( .D(
        new_AGEMA_signal_3709), .CK(clk), .Q(new_AGEMA_signal_3710), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2525_s_current_state_reg ( .D(
        new_AGEMA_signal_3713), .CK(clk), .Q(new_AGEMA_signal_3714), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2529_s_current_state_reg ( .D(
        new_AGEMA_signal_3717), .CK(clk), .Q(new_AGEMA_signal_3718), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2533_s_current_state_reg ( .D(
        new_AGEMA_signal_3721), .CK(clk), .Q(new_AGEMA_signal_3722), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2537_s_current_state_reg ( .D(
        new_AGEMA_signal_3725), .CK(clk), .Q(new_AGEMA_signal_3726), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2541_s_current_state_reg ( .D(
        new_AGEMA_signal_3729), .CK(clk), .Q(new_AGEMA_signal_3730), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2545_s_current_state_reg ( .D(
        new_AGEMA_signal_3733), .CK(clk), .Q(new_AGEMA_signal_3734), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2549_s_current_state_reg ( .D(
        new_AGEMA_signal_3737), .CK(clk), .Q(new_AGEMA_signal_3738), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2553_s_current_state_reg ( .D(
        new_AGEMA_signal_3741), .CK(clk), .Q(new_AGEMA_signal_3742), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2557_s_current_state_reg ( .D(
        new_AGEMA_signal_3745), .CK(clk), .Q(new_AGEMA_signal_3746), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2561_s_current_state_reg ( .D(
        new_AGEMA_signal_3749), .CK(clk), .Q(new_AGEMA_signal_3750), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2565_s_current_state_reg ( .D(
        new_AGEMA_signal_3753), .CK(clk), .Q(new_AGEMA_signal_3754), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2569_s_current_state_reg ( .D(
        new_AGEMA_signal_3757), .CK(clk), .Q(new_AGEMA_signal_3758), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2573_s_current_state_reg ( .D(
        new_AGEMA_signal_3761), .CK(clk), .Q(new_AGEMA_signal_3762), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2577_s_current_state_reg ( .D(
        new_AGEMA_signal_3765), .CK(clk), .Q(new_AGEMA_signal_3766), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2581_s_current_state_reg ( .D(
        new_AGEMA_signal_3769), .CK(clk), .Q(new_AGEMA_signal_3770), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2585_s_current_state_reg ( .D(
        new_AGEMA_signal_3773), .CK(clk), .Q(new_AGEMA_signal_3774), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2589_s_current_state_reg ( .D(
        new_AGEMA_signal_3777), .CK(clk), .Q(new_AGEMA_signal_3778), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2593_s_current_state_reg ( .D(
        new_AGEMA_signal_3781), .CK(clk), .Q(new_AGEMA_signal_3782), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2597_s_current_state_reg ( .D(
        new_AGEMA_signal_3785), .CK(clk), .Q(new_AGEMA_signal_3786), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2601_s_current_state_reg ( .D(
        new_AGEMA_signal_3789), .CK(clk), .Q(new_AGEMA_signal_3790), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2605_s_current_state_reg ( .D(
        new_AGEMA_signal_3793), .CK(clk), .Q(new_AGEMA_signal_3794), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2609_s_current_state_reg ( .D(
        new_AGEMA_signal_3797), .CK(clk), .Q(new_AGEMA_signal_3798), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2613_s_current_state_reg ( .D(
        new_AGEMA_signal_3801), .CK(clk), .Q(new_AGEMA_signal_3802), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2617_s_current_state_reg ( .D(
        new_AGEMA_signal_3805), .CK(clk), .Q(new_AGEMA_signal_3806), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2621_s_current_state_reg ( .D(
        new_AGEMA_signal_3809), .CK(clk), .Q(new_AGEMA_signal_3810), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2625_s_current_state_reg ( .D(
        new_AGEMA_signal_3813), .CK(clk), .Q(new_AGEMA_signal_3814), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2629_s_current_state_reg ( .D(
        new_AGEMA_signal_3817), .CK(clk), .Q(new_AGEMA_signal_3818), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2633_s_current_state_reg ( .D(
        new_AGEMA_signal_3821), .CK(clk), .Q(new_AGEMA_signal_3822), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2637_s_current_state_reg ( .D(
        new_AGEMA_signal_3825), .CK(clk), .Q(new_AGEMA_signal_3826), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2641_s_current_state_reg ( .D(
        new_AGEMA_signal_3829), .CK(clk), .Q(new_AGEMA_signal_3830), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2645_s_current_state_reg ( .D(
        new_AGEMA_signal_3833), .CK(clk), .Q(new_AGEMA_signal_3834), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2649_s_current_state_reg ( .D(
        new_AGEMA_signal_3837), .CK(clk), .Q(new_AGEMA_signal_3838), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2653_s_current_state_reg ( .D(
        new_AGEMA_signal_3841), .CK(clk), .Q(new_AGEMA_signal_3842), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2657_s_current_state_reg ( .D(
        new_AGEMA_signal_3845), .CK(clk), .Q(new_AGEMA_signal_3846), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2661_s_current_state_reg ( .D(
        new_AGEMA_signal_3849), .CK(clk), .Q(new_AGEMA_signal_3850), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2665_s_current_state_reg ( .D(
        new_AGEMA_signal_3853), .CK(clk), .Q(new_AGEMA_signal_3854), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2669_s_current_state_reg ( .D(
        new_AGEMA_signal_3857), .CK(clk), .Q(new_AGEMA_signal_3858), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2673_s_current_state_reg ( .D(
        new_AGEMA_signal_3861), .CK(clk), .Q(new_AGEMA_signal_3862), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2677_s_current_state_reg ( .D(
        new_AGEMA_signal_3865), .CK(clk), .Q(new_AGEMA_signal_3866), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2681_s_current_state_reg ( .D(
        new_AGEMA_signal_3869), .CK(clk), .Q(new_AGEMA_signal_3870), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2685_s_current_state_reg ( .D(
        new_AGEMA_signal_3873), .CK(clk), .Q(new_AGEMA_signal_3874), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2689_s_current_state_reg ( .D(
        new_AGEMA_signal_3877), .CK(clk), .Q(new_AGEMA_signal_3878), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2693_s_current_state_reg ( .D(
        new_AGEMA_signal_3881), .CK(clk), .Q(new_AGEMA_signal_3882), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2697_s_current_state_reg ( .D(
        new_AGEMA_signal_3885), .CK(clk), .Q(new_AGEMA_signal_3886), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2701_s_current_state_reg ( .D(
        new_AGEMA_signal_3889), .CK(clk), .Q(new_AGEMA_signal_3890), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2705_s_current_state_reg ( .D(
        new_AGEMA_signal_3893), .CK(clk), .Q(new_AGEMA_signal_3894), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2709_s_current_state_reg ( .D(
        new_AGEMA_signal_3897), .CK(clk), .Q(new_AGEMA_signal_3898), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2713_s_current_state_reg ( .D(
        new_AGEMA_signal_3901), .CK(clk), .Q(new_AGEMA_signal_3902), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2717_s_current_state_reg ( .D(
        new_AGEMA_signal_3905), .CK(clk), .Q(new_AGEMA_signal_3906), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2721_s_current_state_reg ( .D(
        new_AGEMA_signal_3909), .CK(clk), .Q(new_AGEMA_signal_3910), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2725_s_current_state_reg ( .D(
        new_AGEMA_signal_3913), .CK(clk), .Q(new_AGEMA_signal_3914), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2729_s_current_state_reg ( .D(
        new_AGEMA_signal_3917), .CK(clk), .Q(new_AGEMA_signal_3918), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2733_s_current_state_reg ( .D(
        new_AGEMA_signal_3921), .CK(clk), .Q(new_AGEMA_signal_3922), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2737_s_current_state_reg ( .D(
        new_AGEMA_signal_3925), .CK(clk), .Q(new_AGEMA_signal_3926), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2741_s_current_state_reg ( .D(
        new_AGEMA_signal_3929), .CK(clk), .Q(new_AGEMA_signal_3930), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2745_s_current_state_reg ( .D(
        new_AGEMA_signal_3933), .CK(clk), .Q(new_AGEMA_signal_3934), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2749_s_current_state_reg ( .D(
        new_AGEMA_signal_3937), .CK(clk), .Q(new_AGEMA_signal_3938), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2753_s_current_state_reg ( .D(
        new_AGEMA_signal_3941), .CK(clk), .Q(new_AGEMA_signal_3942), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2757_s_current_state_reg ( .D(
        new_AGEMA_signal_3945), .CK(clk), .Q(new_AGEMA_signal_3946), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2761_s_current_state_reg ( .D(
        new_AGEMA_signal_3949), .CK(clk), .Q(new_AGEMA_signal_3950), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2765_s_current_state_reg ( .D(
        new_AGEMA_signal_3953), .CK(clk), .Q(new_AGEMA_signal_3954), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2769_s_current_state_reg ( .D(
        new_AGEMA_signal_3957), .CK(clk), .Q(new_AGEMA_signal_3958), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2773_s_current_state_reg ( .D(
        new_AGEMA_signal_3961), .CK(clk), .Q(new_AGEMA_signal_3962), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2777_s_current_state_reg ( .D(
        new_AGEMA_signal_3965), .CK(clk), .Q(new_AGEMA_signal_3966), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2781_s_current_state_reg ( .D(
        new_AGEMA_signal_3969), .CK(clk), .Q(new_AGEMA_signal_3970), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2785_s_current_state_reg ( .D(
        new_AGEMA_signal_3973), .CK(clk), .Q(new_AGEMA_signal_3974), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2789_s_current_state_reg ( .D(
        new_AGEMA_signal_3977), .CK(clk), .Q(new_AGEMA_signal_3978), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2793_s_current_state_reg ( .D(
        new_AGEMA_signal_3981), .CK(clk), .Q(new_AGEMA_signal_3982), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2797_s_current_state_reg ( .D(
        new_AGEMA_signal_3985), .CK(clk), .Q(new_AGEMA_signal_3986), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2801_s_current_state_reg ( .D(
        new_AGEMA_signal_3989), .CK(clk), .Q(new_AGEMA_signal_3990), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2805_s_current_state_reg ( .D(
        new_AGEMA_signal_3993), .CK(clk), .Q(new_AGEMA_signal_3994), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2809_s_current_state_reg ( .D(
        new_AGEMA_signal_3997), .CK(clk), .Q(new_AGEMA_signal_3998), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2813_s_current_state_reg ( .D(
        new_AGEMA_signal_4001), .CK(clk), .Q(new_AGEMA_signal_4002), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2817_s_current_state_reg ( .D(
        new_AGEMA_signal_4005), .CK(clk), .Q(new_AGEMA_signal_4006), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2821_s_current_state_reg ( .D(
        new_AGEMA_signal_4009), .CK(clk), .Q(new_AGEMA_signal_4010), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2825_s_current_state_reg ( .D(
        new_AGEMA_signal_4013), .CK(clk), .Q(new_AGEMA_signal_4014), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2829_s_current_state_reg ( .D(
        new_AGEMA_signal_4017), .CK(clk), .Q(new_AGEMA_signal_4018), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2833_s_current_state_reg ( .D(
        new_AGEMA_signal_4021), .CK(clk), .Q(new_AGEMA_signal_4022), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2837_s_current_state_reg ( .D(
        new_AGEMA_signal_4025), .CK(clk), .Q(new_AGEMA_signal_4026), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2841_s_current_state_reg ( .D(
        new_AGEMA_signal_4029), .CK(clk), .Q(new_AGEMA_signal_4030), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2845_s_current_state_reg ( .D(
        new_AGEMA_signal_4033), .CK(clk), .Q(new_AGEMA_signal_4034), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2849_s_current_state_reg ( .D(
        new_AGEMA_signal_4037), .CK(clk), .Q(new_AGEMA_signal_4038), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2853_s_current_state_reg ( .D(
        new_AGEMA_signal_4041), .CK(clk), .Q(new_AGEMA_signal_4042), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2857_s_current_state_reg ( .D(
        new_AGEMA_signal_4045), .CK(clk), .Q(new_AGEMA_signal_4046), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2861_s_current_state_reg ( .D(
        new_AGEMA_signal_4049), .CK(clk), .Q(new_AGEMA_signal_4050), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2865_s_current_state_reg ( .D(
        new_AGEMA_signal_4053), .CK(clk), .Q(new_AGEMA_signal_4054), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2869_s_current_state_reg ( .D(
        new_AGEMA_signal_4057), .CK(clk), .Q(new_AGEMA_signal_4058), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2873_s_current_state_reg ( .D(
        new_AGEMA_signal_4061), .CK(clk), .Q(new_AGEMA_signal_4062), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2877_s_current_state_reg ( .D(
        new_AGEMA_signal_4065), .CK(clk), .Q(new_AGEMA_signal_4066), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2881_s_current_state_reg ( .D(
        new_AGEMA_signal_4069), .CK(clk), .Q(new_AGEMA_signal_4070), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2885_s_current_state_reg ( .D(
        new_AGEMA_signal_4073), .CK(clk), .Q(new_AGEMA_signal_4074), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2889_s_current_state_reg ( .D(
        new_AGEMA_signal_4077), .CK(clk), .Q(new_AGEMA_signal_4078), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2893_s_current_state_reg ( .D(
        new_AGEMA_signal_4081), .CK(clk), .Q(new_AGEMA_signal_4082), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2897_s_current_state_reg ( .D(
        new_AGEMA_signal_4085), .CK(clk), .Q(new_AGEMA_signal_4086), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2901_s_current_state_reg ( .D(
        new_AGEMA_signal_4089), .CK(clk), .Q(new_AGEMA_signal_4090), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1454_s_current_state_reg ( .D(
        new_AGEMA_signal_2190), .CK(clk), .Q(new_AGEMA_signal_2643), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1458_s_current_state_reg ( .D(
        new_AGEMA_signal_2646), .CK(clk), .Q(new_AGEMA_signal_2647), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1462_s_current_state_reg ( .D(
        new_AGEMA_signal_2650), .CK(clk), .Q(new_AGEMA_signal_2651), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1466_s_current_state_reg ( .D(
        new_AGEMA_signal_2654), .CK(clk), .Q(new_AGEMA_signal_2655), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1470_s_current_state_reg ( .D(
        new_AGEMA_signal_2658), .CK(clk), .Q(new_AGEMA_signal_2659), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1474_s_current_state_reg ( .D(
        new_AGEMA_signal_2662), .CK(clk), .Q(new_AGEMA_signal_2663), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1478_s_current_state_reg ( .D(
        new_AGEMA_signal_2666), .CK(clk), .Q(new_AGEMA_signal_2667), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1482_s_current_state_reg ( .D(
        new_AGEMA_signal_2670), .CK(clk), .Q(new_AGEMA_signal_2671), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1486_s_current_state_reg ( .D(
        new_AGEMA_signal_2674), .CK(clk), .Q(new_AGEMA_signal_2675), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1490_s_current_state_reg ( .D(
        new_AGEMA_signal_2678), .CK(clk), .Q(new_AGEMA_signal_2679), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1494_s_current_state_reg ( .D(
        new_AGEMA_signal_2682), .CK(clk), .Q(new_AGEMA_signal_2683), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1498_s_current_state_reg ( .D(
        new_AGEMA_signal_2686), .CK(clk), .Q(new_AGEMA_signal_2687), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1502_s_current_state_reg ( .D(
        new_AGEMA_signal_2690), .CK(clk), .Q(new_AGEMA_signal_2691), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1506_s_current_state_reg ( .D(
        new_AGEMA_signal_2694), .CK(clk), .Q(new_AGEMA_signal_2695), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1510_s_current_state_reg ( .D(
        new_AGEMA_signal_2698), .CK(clk), .Q(new_AGEMA_signal_2699), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1514_s_current_state_reg ( .D(
        new_AGEMA_signal_2702), .CK(clk), .Q(new_AGEMA_signal_2703), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1518_s_current_state_reg ( .D(
        new_AGEMA_signal_2706), .CK(clk), .Q(new_AGEMA_signal_2707), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1522_s_current_state_reg ( .D(
        new_AGEMA_signal_2710), .CK(clk), .Q(new_AGEMA_signal_2711), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1526_s_current_state_reg ( .D(
        new_AGEMA_signal_2714), .CK(clk), .Q(new_AGEMA_signal_2715), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1530_s_current_state_reg ( .D(
        new_AGEMA_signal_2718), .CK(clk), .Q(new_AGEMA_signal_2719), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1534_s_current_state_reg ( .D(
        new_AGEMA_signal_2722), .CK(clk), .Q(new_AGEMA_signal_2723), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1538_s_current_state_reg ( .D(
        new_AGEMA_signal_2726), .CK(clk), .Q(new_AGEMA_signal_2727), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1542_s_current_state_reg ( .D(
        new_AGEMA_signal_2730), .CK(clk), .Q(new_AGEMA_signal_2731), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1546_s_current_state_reg ( .D(
        new_AGEMA_signal_2734), .CK(clk), .Q(new_AGEMA_signal_2735), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1550_s_current_state_reg ( .D(
        new_AGEMA_signal_2738), .CK(clk), .Q(new_AGEMA_signal_2739), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1554_s_current_state_reg ( .D(
        new_AGEMA_signal_2742), .CK(clk), .Q(new_AGEMA_signal_2743), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1558_s_current_state_reg ( .D(
        new_AGEMA_signal_2746), .CK(clk), .Q(new_AGEMA_signal_2747), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1562_s_current_state_reg ( .D(
        new_AGEMA_signal_2750), .CK(clk), .Q(new_AGEMA_signal_2751), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1566_s_current_state_reg ( .D(
        new_AGEMA_signal_2754), .CK(clk), .Q(new_AGEMA_signal_2755), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1570_s_current_state_reg ( .D(
        new_AGEMA_signal_2758), .CK(clk), .Q(new_AGEMA_signal_2759), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1574_s_current_state_reg ( .D(
        new_AGEMA_signal_2762), .CK(clk), .Q(new_AGEMA_signal_2763), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1578_s_current_state_reg ( .D(
        new_AGEMA_signal_2766), .CK(clk), .Q(new_AGEMA_signal_2767), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1582_s_current_state_reg ( .D(
        new_AGEMA_signal_2770), .CK(clk), .Q(new_AGEMA_signal_2771), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1586_s_current_state_reg ( .D(
        new_AGEMA_signal_2774), .CK(clk), .Q(new_AGEMA_signal_2775), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1590_s_current_state_reg ( .D(
        new_AGEMA_signal_2778), .CK(clk), .Q(new_AGEMA_signal_2779), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1594_s_current_state_reg ( .D(
        new_AGEMA_signal_2782), .CK(clk), .Q(new_AGEMA_signal_2783), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1598_s_current_state_reg ( .D(
        new_AGEMA_signal_2786), .CK(clk), .Q(new_AGEMA_signal_2787), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1602_s_current_state_reg ( .D(
        new_AGEMA_signal_2790), .CK(clk), .Q(new_AGEMA_signal_2791), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1606_s_current_state_reg ( .D(
        new_AGEMA_signal_2794), .CK(clk), .Q(new_AGEMA_signal_2795), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1610_s_current_state_reg ( .D(
        new_AGEMA_signal_2798), .CK(clk), .Q(new_AGEMA_signal_2799), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1614_s_current_state_reg ( .D(
        new_AGEMA_signal_2802), .CK(clk), .Q(new_AGEMA_signal_2803), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1618_s_current_state_reg ( .D(
        new_AGEMA_signal_2806), .CK(clk), .Q(new_AGEMA_signal_2807), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1622_s_current_state_reg ( .D(
        new_AGEMA_signal_2810), .CK(clk), .Q(new_AGEMA_signal_2811), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1626_s_current_state_reg ( .D(
        new_AGEMA_signal_2814), .CK(clk), .Q(new_AGEMA_signal_2815), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1630_s_current_state_reg ( .D(
        new_AGEMA_signal_2818), .CK(clk), .Q(new_AGEMA_signal_2819), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1634_s_current_state_reg ( .D(
        new_AGEMA_signal_2822), .CK(clk), .Q(new_AGEMA_signal_2823), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1638_s_current_state_reg ( .D(
        new_AGEMA_signal_2826), .CK(clk), .Q(new_AGEMA_signal_2827), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1642_s_current_state_reg ( .D(
        new_AGEMA_signal_2830), .CK(clk), .Q(new_AGEMA_signal_2831), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1646_s_current_state_reg ( .D(
        new_AGEMA_signal_2834), .CK(clk), .Q(new_AGEMA_signal_2835), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1650_s_current_state_reg ( .D(
        new_AGEMA_signal_2838), .CK(clk), .Q(new_AGEMA_signal_2839), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1654_s_current_state_reg ( .D(
        new_AGEMA_signal_2842), .CK(clk), .Q(new_AGEMA_signal_2843), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1658_s_current_state_reg ( .D(
        new_AGEMA_signal_2846), .CK(clk), .Q(new_AGEMA_signal_2847), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1662_s_current_state_reg ( .D(
        new_AGEMA_signal_2850), .CK(clk), .Q(new_AGEMA_signal_2851), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1666_s_current_state_reg ( .D(
        new_AGEMA_signal_2854), .CK(clk), .Q(new_AGEMA_signal_2855), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1670_s_current_state_reg ( .D(
        new_AGEMA_signal_2858), .CK(clk), .Q(new_AGEMA_signal_2859), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1674_s_current_state_reg ( .D(
        new_AGEMA_signal_2862), .CK(clk), .Q(new_AGEMA_signal_2863), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1678_s_current_state_reg ( .D(
        new_AGEMA_signal_2866), .CK(clk), .Q(new_AGEMA_signal_2867), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1682_s_current_state_reg ( .D(
        new_AGEMA_signal_2870), .CK(clk), .Q(new_AGEMA_signal_2871), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1686_s_current_state_reg ( .D(
        new_AGEMA_signal_2874), .CK(clk), .Q(new_AGEMA_signal_2875), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1690_s_current_state_reg ( .D(
        new_AGEMA_signal_2878), .CK(clk), .Q(new_AGEMA_signal_2879), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1694_s_current_state_reg ( .D(
        new_AGEMA_signal_2882), .CK(clk), .Q(new_AGEMA_signal_2883), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1698_s_current_state_reg ( .D(
        new_AGEMA_signal_2886), .CK(clk), .Q(new_AGEMA_signal_2887), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1702_s_current_state_reg ( .D(
        new_AGEMA_signal_2890), .CK(clk), .Q(new_AGEMA_signal_2891), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1706_s_current_state_reg ( .D(
        new_AGEMA_signal_2894), .CK(clk), .Q(new_AGEMA_signal_2895), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1710_s_current_state_reg ( .D(
        new_AGEMA_signal_2898), .CK(clk), .Q(new_AGEMA_signal_2899), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1716_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_T2), .CK(clk), .Q(new_AGEMA_signal_2905), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1718_s_current_state_reg ( .D(
        new_AGEMA_signal_1549), .CK(clk), .Q(new_AGEMA_signal_2907), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1726_s_current_state_reg ( .D(
        new_AGEMA_signal_2914), .CK(clk), .Q(new_AGEMA_signal_2915), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1730_s_current_state_reg ( .D(
        new_AGEMA_signal_2918), .CK(clk), .Q(new_AGEMA_signal_2919), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1732_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_YY_1_), .CK(clk), .Q(new_AGEMA_signal_2921), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1734_s_current_state_reg ( .D(
        new_AGEMA_signal_1724), .CK(clk), .Q(new_AGEMA_signal_2923), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1740_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_T2), .CK(clk), .Q(new_AGEMA_signal_2929), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1742_s_current_state_reg ( .D(
        new_AGEMA_signal_1552), .CK(clk), .Q(new_AGEMA_signal_2931), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1750_s_current_state_reg ( .D(
        new_AGEMA_signal_2938), .CK(clk), .Q(new_AGEMA_signal_2939), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1754_s_current_state_reg ( .D(
        new_AGEMA_signal_2942), .CK(clk), .Q(new_AGEMA_signal_2943), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1756_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_YY_1_), .CK(clk), .Q(new_AGEMA_signal_2945), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1758_s_current_state_reg ( .D(
        new_AGEMA_signal_1726), .CK(clk), .Q(new_AGEMA_signal_2947), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1764_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_T2), .CK(clk), .Q(new_AGEMA_signal_2953), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1766_s_current_state_reg ( .D(
        new_AGEMA_signal_1555), .CK(clk), .Q(new_AGEMA_signal_2955), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1774_s_current_state_reg ( .D(
        new_AGEMA_signal_2962), .CK(clk), .Q(new_AGEMA_signal_2963), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1778_s_current_state_reg ( .D(
        new_AGEMA_signal_2966), .CK(clk), .Q(new_AGEMA_signal_2967), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1780_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_YY_1_), .CK(clk), .Q(new_AGEMA_signal_2969), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1782_s_current_state_reg ( .D(
        new_AGEMA_signal_1728), .CK(clk), .Q(new_AGEMA_signal_2971), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1788_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_T2), .CK(clk), .Q(new_AGEMA_signal_2977), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1790_s_current_state_reg ( .D(
        new_AGEMA_signal_1558), .CK(clk), .Q(new_AGEMA_signal_2979), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1798_s_current_state_reg ( .D(
        new_AGEMA_signal_2986), .CK(clk), .Q(new_AGEMA_signal_2987), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1802_s_current_state_reg ( .D(
        new_AGEMA_signal_2990), .CK(clk), .Q(new_AGEMA_signal_2991), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1804_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_YY_1_), .CK(clk), .Q(new_AGEMA_signal_2993), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1806_s_current_state_reg ( .D(
        new_AGEMA_signal_1730), .CK(clk), .Q(new_AGEMA_signal_2995), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1812_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_T2), .CK(clk), .Q(new_AGEMA_signal_3001), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1814_s_current_state_reg ( .D(
        new_AGEMA_signal_1561), .CK(clk), .Q(new_AGEMA_signal_3003), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1822_s_current_state_reg ( .D(
        new_AGEMA_signal_3010), .CK(clk), .Q(new_AGEMA_signal_3011), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1826_s_current_state_reg ( .D(
        new_AGEMA_signal_3014), .CK(clk), .Q(new_AGEMA_signal_3015), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1828_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3017), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1830_s_current_state_reg ( .D(
        new_AGEMA_signal_1732), .CK(clk), .Q(new_AGEMA_signal_3019), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1836_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_T2), .CK(clk), .Q(new_AGEMA_signal_3025), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1838_s_current_state_reg ( .D(
        new_AGEMA_signal_1564), .CK(clk), .Q(new_AGEMA_signal_3027), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1846_s_current_state_reg ( .D(
        new_AGEMA_signal_3034), .CK(clk), .Q(new_AGEMA_signal_3035), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1850_s_current_state_reg ( .D(
        new_AGEMA_signal_3038), .CK(clk), .Q(new_AGEMA_signal_3039), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1852_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3041), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1854_s_current_state_reg ( .D(
        new_AGEMA_signal_1734), .CK(clk), .Q(new_AGEMA_signal_3043), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1860_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_T2), .CK(clk), .Q(new_AGEMA_signal_3049), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1862_s_current_state_reg ( .D(
        new_AGEMA_signal_1567), .CK(clk), .Q(new_AGEMA_signal_3051), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1870_s_current_state_reg ( .D(
        new_AGEMA_signal_3058), .CK(clk), .Q(new_AGEMA_signal_3059), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1874_s_current_state_reg ( .D(
        new_AGEMA_signal_3062), .CK(clk), .Q(new_AGEMA_signal_3063), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1876_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3065), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1878_s_current_state_reg ( .D(
        new_AGEMA_signal_1736), .CK(clk), .Q(new_AGEMA_signal_3067), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1884_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_T2), .CK(clk), .Q(new_AGEMA_signal_3073), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1886_s_current_state_reg ( .D(
        new_AGEMA_signal_1570), .CK(clk), .Q(new_AGEMA_signal_3075), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1894_s_current_state_reg ( .D(
        new_AGEMA_signal_3082), .CK(clk), .Q(new_AGEMA_signal_3083), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1898_s_current_state_reg ( .D(
        new_AGEMA_signal_3086), .CK(clk), .Q(new_AGEMA_signal_3087), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1900_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3089), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1902_s_current_state_reg ( .D(
        new_AGEMA_signal_1738), .CK(clk), .Q(new_AGEMA_signal_3091), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1908_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_T2), .CK(clk), .Q(new_AGEMA_signal_3097), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1910_s_current_state_reg ( .D(
        new_AGEMA_signal_1573), .CK(clk), .Q(new_AGEMA_signal_3099), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1918_s_current_state_reg ( .D(
        new_AGEMA_signal_3106), .CK(clk), .Q(new_AGEMA_signal_3107), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1922_s_current_state_reg ( .D(
        new_AGEMA_signal_3110), .CK(clk), .Q(new_AGEMA_signal_3111), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1924_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3113), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1926_s_current_state_reg ( .D(
        new_AGEMA_signal_1740), .CK(clk), .Q(new_AGEMA_signal_3115), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1932_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_T2), .CK(clk), .Q(new_AGEMA_signal_3121), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1934_s_current_state_reg ( .D(
        new_AGEMA_signal_1576), .CK(clk), .Q(new_AGEMA_signal_3123), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1942_s_current_state_reg ( .D(
        new_AGEMA_signal_3130), .CK(clk), .Q(new_AGEMA_signal_3131), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1946_s_current_state_reg ( .D(
        new_AGEMA_signal_3134), .CK(clk), .Q(new_AGEMA_signal_3135), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1948_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3137), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1950_s_current_state_reg ( .D(
        new_AGEMA_signal_1742), .CK(clk), .Q(new_AGEMA_signal_3139), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1956_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_T2), .CK(clk), .Q(new_AGEMA_signal_3145), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1958_s_current_state_reg ( .D(
        new_AGEMA_signal_1579), .CK(clk), .Q(new_AGEMA_signal_3147), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1966_s_current_state_reg ( .D(
        new_AGEMA_signal_3154), .CK(clk), .Q(new_AGEMA_signal_3155), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1970_s_current_state_reg ( .D(
        new_AGEMA_signal_3158), .CK(clk), .Q(new_AGEMA_signal_3159), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1972_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3161), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1974_s_current_state_reg ( .D(
        new_AGEMA_signal_1744), .CK(clk), .Q(new_AGEMA_signal_3163), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1980_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_T2), .CK(clk), .Q(new_AGEMA_signal_3169), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1982_s_current_state_reg ( .D(
        new_AGEMA_signal_1582), .CK(clk), .Q(new_AGEMA_signal_3171), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1990_s_current_state_reg ( .D(
        new_AGEMA_signal_3178), .CK(clk), .Q(new_AGEMA_signal_3179), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1994_s_current_state_reg ( .D(
        new_AGEMA_signal_3182), .CK(clk), .Q(new_AGEMA_signal_3183), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1996_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3185), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1998_s_current_state_reg ( .D(
        new_AGEMA_signal_1746), .CK(clk), .Q(new_AGEMA_signal_3187), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2004_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_T2), .CK(clk), .Q(new_AGEMA_signal_3193), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2006_s_current_state_reg ( .D(
        new_AGEMA_signal_1585), .CK(clk), .Q(new_AGEMA_signal_3195), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2014_s_current_state_reg ( .D(
        new_AGEMA_signal_3202), .CK(clk), .Q(new_AGEMA_signal_3203), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2018_s_current_state_reg ( .D(
        new_AGEMA_signal_3206), .CK(clk), .Q(new_AGEMA_signal_3207), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2020_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3209), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2022_s_current_state_reg ( .D(
        new_AGEMA_signal_1748), .CK(clk), .Q(new_AGEMA_signal_3211), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2028_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_T2), .CK(clk), .Q(new_AGEMA_signal_3217), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2030_s_current_state_reg ( .D(
        new_AGEMA_signal_1588), .CK(clk), .Q(new_AGEMA_signal_3219), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2038_s_current_state_reg ( .D(
        new_AGEMA_signal_3226), .CK(clk), .Q(new_AGEMA_signal_3227), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2042_s_current_state_reg ( .D(
        new_AGEMA_signal_3230), .CK(clk), .Q(new_AGEMA_signal_3231), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2044_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3233), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2046_s_current_state_reg ( .D(
        new_AGEMA_signal_1750), .CK(clk), .Q(new_AGEMA_signal_3235), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2052_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_T2), .CK(clk), .Q(new_AGEMA_signal_3241), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2054_s_current_state_reg ( .D(
        new_AGEMA_signal_1591), .CK(clk), .Q(new_AGEMA_signal_3243), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2062_s_current_state_reg ( .D(
        new_AGEMA_signal_3250), .CK(clk), .Q(new_AGEMA_signal_3251), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2066_s_current_state_reg ( .D(
        new_AGEMA_signal_3254), .CK(clk), .Q(new_AGEMA_signal_3255), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2068_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3257), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2070_s_current_state_reg ( .D(
        new_AGEMA_signal_1752), .CK(clk), .Q(new_AGEMA_signal_3259), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2076_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_T2), .CK(clk), .Q(new_AGEMA_signal_3265), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2078_s_current_state_reg ( .D(
        new_AGEMA_signal_1594), .CK(clk), .Q(new_AGEMA_signal_3267), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2086_s_current_state_reg ( .D(
        new_AGEMA_signal_3274), .CK(clk), .Q(new_AGEMA_signal_3275), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2090_s_current_state_reg ( .D(
        new_AGEMA_signal_3278), .CK(clk), .Q(new_AGEMA_signal_3279), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2092_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_YY_1_), .CK(clk), .Q(new_AGEMA_signal_3281), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2094_s_current_state_reg ( .D(
        new_AGEMA_signal_1754), .CK(clk), .Q(new_AGEMA_signal_3283), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2098_s_current_state_reg ( .D(
        new_AGEMA_signal_3286), .CK(clk), .Q(new_AGEMA_signal_3287), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2102_s_current_state_reg ( .D(
        new_AGEMA_signal_3290), .CK(clk), .Q(new_AGEMA_signal_3291), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2106_s_current_state_reg ( .D(
        new_AGEMA_signal_3294), .CK(clk), .Q(new_AGEMA_signal_3295), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2110_s_current_state_reg ( .D(
        new_AGEMA_signal_3298), .CK(clk), .Q(new_AGEMA_signal_3299), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2114_s_current_state_reg ( .D(
        new_AGEMA_signal_3302), .CK(clk), .Q(new_AGEMA_signal_3303), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2118_s_current_state_reg ( .D(
        new_AGEMA_signal_3306), .CK(clk), .Q(new_AGEMA_signal_3307), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2122_s_current_state_reg ( .D(
        new_AGEMA_signal_3310), .CK(clk), .Q(new_AGEMA_signal_3311), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2126_s_current_state_reg ( .D(
        new_AGEMA_signal_3314), .CK(clk), .Q(new_AGEMA_signal_3315), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2130_s_current_state_reg ( .D(
        new_AGEMA_signal_3318), .CK(clk), .Q(new_AGEMA_signal_3319), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2134_s_current_state_reg ( .D(
        new_AGEMA_signal_3322), .CK(clk), .Q(new_AGEMA_signal_3323), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2138_s_current_state_reg ( .D(
        new_AGEMA_signal_3326), .CK(clk), .Q(new_AGEMA_signal_3327), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2142_s_current_state_reg ( .D(
        new_AGEMA_signal_3330), .CK(clk), .Q(new_AGEMA_signal_3331), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2146_s_current_state_reg ( .D(
        new_AGEMA_signal_3334), .CK(clk), .Q(new_AGEMA_signal_3335), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2150_s_current_state_reg ( .D(
        new_AGEMA_signal_3338), .CK(clk), .Q(new_AGEMA_signal_3339), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2154_s_current_state_reg ( .D(
        new_AGEMA_signal_3342), .CK(clk), .Q(new_AGEMA_signal_3343), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2158_s_current_state_reg ( .D(
        new_AGEMA_signal_3346), .CK(clk), .Q(new_AGEMA_signal_3347), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2162_s_current_state_reg ( .D(
        new_AGEMA_signal_3350), .CK(clk), .Q(new_AGEMA_signal_3351), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2166_s_current_state_reg ( .D(
        new_AGEMA_signal_3354), .CK(clk), .Q(new_AGEMA_signal_3355), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2170_s_current_state_reg ( .D(
        new_AGEMA_signal_3358), .CK(clk), .Q(new_AGEMA_signal_3359), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2174_s_current_state_reg ( .D(
        new_AGEMA_signal_3362), .CK(clk), .Q(new_AGEMA_signal_3363), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2178_s_current_state_reg ( .D(
        new_AGEMA_signal_3366), .CK(clk), .Q(new_AGEMA_signal_3367), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2182_s_current_state_reg ( .D(
        new_AGEMA_signal_3370), .CK(clk), .Q(new_AGEMA_signal_3371), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2186_s_current_state_reg ( .D(
        new_AGEMA_signal_3374), .CK(clk), .Q(new_AGEMA_signal_3375), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2190_s_current_state_reg ( .D(
        new_AGEMA_signal_3378), .CK(clk), .Q(new_AGEMA_signal_3379), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2194_s_current_state_reg ( .D(
        new_AGEMA_signal_3382), .CK(clk), .Q(new_AGEMA_signal_3383), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2198_s_current_state_reg ( .D(
        new_AGEMA_signal_3386), .CK(clk), .Q(new_AGEMA_signal_3387), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2202_s_current_state_reg ( .D(
        new_AGEMA_signal_3390), .CK(clk), .Q(new_AGEMA_signal_3391), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2206_s_current_state_reg ( .D(
        new_AGEMA_signal_3394), .CK(clk), .Q(new_AGEMA_signal_3395), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2210_s_current_state_reg ( .D(
        new_AGEMA_signal_3398), .CK(clk), .Q(new_AGEMA_signal_3399), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2214_s_current_state_reg ( .D(
        new_AGEMA_signal_3402), .CK(clk), .Q(new_AGEMA_signal_3403), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2218_s_current_state_reg ( .D(
        new_AGEMA_signal_3406), .CK(clk), .Q(new_AGEMA_signal_3407), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2222_s_current_state_reg ( .D(
        new_AGEMA_signal_3410), .CK(clk), .Q(new_AGEMA_signal_3411), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2226_s_current_state_reg ( .D(
        new_AGEMA_signal_3414), .CK(clk), .Q(new_AGEMA_signal_3415), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2230_s_current_state_reg ( .D(
        new_AGEMA_signal_3418), .CK(clk), .Q(new_AGEMA_signal_3419), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2234_s_current_state_reg ( .D(
        new_AGEMA_signal_3422), .CK(clk), .Q(new_AGEMA_signal_3423), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2238_s_current_state_reg ( .D(
        new_AGEMA_signal_3426), .CK(clk), .Q(new_AGEMA_signal_3427), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2240_s_current_state_reg ( .D(StateRegInput[63]), 
        .CK(clk), .Q(new_AGEMA_signal_3429), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2242_s_current_state_reg ( .D(
        new_AGEMA_signal_2103), .CK(clk), .Q(new_AGEMA_signal_3431), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2244_s_current_state_reg ( .D(StateRegInput[62]), 
        .CK(clk), .Q(new_AGEMA_signal_3433), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2246_s_current_state_reg ( .D(
        new_AGEMA_signal_2060), .CK(clk), .Q(new_AGEMA_signal_3435), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2248_s_current_state_reg ( .D(StateRegInput[59]), 
        .CK(clk), .Q(new_AGEMA_signal_3437), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2250_s_current_state_reg ( .D(
        new_AGEMA_signal_2006), .CK(clk), .Q(new_AGEMA_signal_3439), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2252_s_current_state_reg ( .D(StateRegInput[58]), 
        .CK(clk), .Q(new_AGEMA_signal_3441), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2254_s_current_state_reg ( .D(
        new_AGEMA_signal_1946), .CK(clk), .Q(new_AGEMA_signal_3443), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2256_s_current_state_reg ( .D(StateRegInput[55]), 
        .CK(clk), .Q(new_AGEMA_signal_3445), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2258_s_current_state_reg ( .D(
        new_AGEMA_signal_2004), .CK(clk), .Q(new_AGEMA_signal_3447), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2260_s_current_state_reg ( .D(StateRegInput[54]), 
        .CK(clk), .Q(new_AGEMA_signal_3449), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2262_s_current_state_reg ( .D(
        new_AGEMA_signal_1944), .CK(clk), .Q(new_AGEMA_signal_3451), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2264_s_current_state_reg ( .D(StateRegInput[51]), 
        .CK(clk), .Q(new_AGEMA_signal_3453), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2266_s_current_state_reg ( .D(
        new_AGEMA_signal_2002), .CK(clk), .Q(new_AGEMA_signal_3455), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2268_s_current_state_reg ( .D(StateRegInput[50]), 
        .CK(clk), .Q(new_AGEMA_signal_3457), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2270_s_current_state_reg ( .D(
        new_AGEMA_signal_1942), .CK(clk), .Q(new_AGEMA_signal_3459), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2272_s_current_state_reg ( .D(StateRegInput[47]), 
        .CK(clk), .Q(new_AGEMA_signal_3461), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2274_s_current_state_reg ( .D(
        new_AGEMA_signal_2000), .CK(clk), .Q(new_AGEMA_signal_3463), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2276_s_current_state_reg ( .D(StateRegInput[46]), 
        .CK(clk), .Q(new_AGEMA_signal_3465), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2278_s_current_state_reg ( .D(
        new_AGEMA_signal_1940), .CK(clk), .Q(new_AGEMA_signal_3467), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2280_s_current_state_reg ( .D(StateRegInput[43]), 
        .CK(clk), .Q(new_AGEMA_signal_3469), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2282_s_current_state_reg ( .D(
        new_AGEMA_signal_1878), .CK(clk), .Q(new_AGEMA_signal_3471), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2284_s_current_state_reg ( .D(StateRegInput[42]), 
        .CK(clk), .Q(new_AGEMA_signal_3473), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2286_s_current_state_reg ( .D(
        new_AGEMA_signal_1825), .CK(clk), .Q(new_AGEMA_signal_3475), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2288_s_current_state_reg ( .D(StateRegInput[39]), 
        .CK(clk), .Q(new_AGEMA_signal_3477), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2290_s_current_state_reg ( .D(
        new_AGEMA_signal_1876), .CK(clk), .Q(new_AGEMA_signal_3479), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2292_s_current_state_reg ( .D(StateRegInput[38]), 
        .CK(clk), .Q(new_AGEMA_signal_3481), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2294_s_current_state_reg ( .D(
        new_AGEMA_signal_1823), .CK(clk), .Q(new_AGEMA_signal_3483), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2296_s_current_state_reg ( .D(StateRegInput[35]), 
        .CK(clk), .Q(new_AGEMA_signal_3485), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2298_s_current_state_reg ( .D(
        new_AGEMA_signal_1874), .CK(clk), .Q(new_AGEMA_signal_3487), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2300_s_current_state_reg ( .D(StateRegInput[34]), 
        .CK(clk), .Q(new_AGEMA_signal_3489), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2302_s_current_state_reg ( .D(
        new_AGEMA_signal_1821), .CK(clk), .Q(new_AGEMA_signal_3491), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2304_s_current_state_reg ( .D(StateRegInput[31]), 
        .CK(clk), .Q(new_AGEMA_signal_3493), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2306_s_current_state_reg ( .D(
        new_AGEMA_signal_1992), .CK(clk), .Q(new_AGEMA_signal_3495), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2308_s_current_state_reg ( .D(StateRegInput[30]), 
        .CK(clk), .Q(new_AGEMA_signal_3497), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2310_s_current_state_reg ( .D(
        new_AGEMA_signal_1932), .CK(clk), .Q(new_AGEMA_signal_3499), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2312_s_current_state_reg ( .D(StateRegInput[27]), 
        .CK(clk), .Q(new_AGEMA_signal_3501), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2314_s_current_state_reg ( .D(
        new_AGEMA_signal_2091), .CK(clk), .Q(new_AGEMA_signal_3503), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2316_s_current_state_reg ( .D(StateRegInput[26]), 
        .CK(clk), .Q(new_AGEMA_signal_3505), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2318_s_current_state_reg ( .D(
        new_AGEMA_signal_2048), .CK(clk), .Q(new_AGEMA_signal_3507), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2320_s_current_state_reg ( .D(StateRegInput[23]), 
        .CK(clk), .Q(new_AGEMA_signal_3509), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2322_s_current_state_reg ( .D(
        new_AGEMA_signal_1990), .CK(clk), .Q(new_AGEMA_signal_3511), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2324_s_current_state_reg ( .D(StateRegInput[22]), 
        .CK(clk), .Q(new_AGEMA_signal_3513), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2326_s_current_state_reg ( .D(
        new_AGEMA_signal_1930), .CK(clk), .Q(new_AGEMA_signal_3515), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2328_s_current_state_reg ( .D(StateRegInput[19]), 
        .CK(clk), .Q(new_AGEMA_signal_3517), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2330_s_current_state_reg ( .D(
        new_AGEMA_signal_1988), .CK(clk), .Q(new_AGEMA_signal_3519), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2332_s_current_state_reg ( .D(StateRegInput[18]), 
        .CK(clk), .Q(new_AGEMA_signal_3521), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2334_s_current_state_reg ( .D(
        new_AGEMA_signal_1928), .CK(clk), .Q(new_AGEMA_signal_3523), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2336_s_current_state_reg ( .D(StateRegInput[15]), 
        .CK(clk), .Q(new_AGEMA_signal_3525), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2338_s_current_state_reg ( .D(
        new_AGEMA_signal_2085), .CK(clk), .Q(new_AGEMA_signal_3527), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2340_s_current_state_reg ( .D(StateRegInput[14]), 
        .CK(clk), .Q(new_AGEMA_signal_3529), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2342_s_current_state_reg ( .D(
        new_AGEMA_signal_2042), .CK(clk), .Q(new_AGEMA_signal_3531), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2344_s_current_state_reg ( .D(StateRegInput[11]), 
        .CK(clk), .Q(new_AGEMA_signal_3533), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2346_s_current_state_reg ( .D(
        new_AGEMA_signal_1986), .CK(clk), .Q(new_AGEMA_signal_3535), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2348_s_current_state_reg ( .D(StateRegInput[10]), 
        .CK(clk), .Q(new_AGEMA_signal_3537), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2350_s_current_state_reg ( .D(
        new_AGEMA_signal_1926), .CK(clk), .Q(new_AGEMA_signal_3539), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2352_s_current_state_reg ( .D(StateRegInput[7]), 
        .CK(clk), .Q(new_AGEMA_signal_3541), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2354_s_current_state_reg ( .D(
        new_AGEMA_signal_1984), .CK(clk), .Q(new_AGEMA_signal_3543), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2356_s_current_state_reg ( .D(StateRegInput[6]), 
        .CK(clk), .Q(new_AGEMA_signal_3545), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2358_s_current_state_reg ( .D(
        new_AGEMA_signal_1924), .CK(clk), .Q(new_AGEMA_signal_3547), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2360_s_current_state_reg ( .D(StateRegInput[3]), 
        .CK(clk), .Q(new_AGEMA_signal_3549), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2362_s_current_state_reg ( .D(
        new_AGEMA_signal_1982), .CK(clk), .Q(new_AGEMA_signal_3551), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2364_s_current_state_reg ( .D(StateRegInput[2]), 
        .CK(clk), .Q(new_AGEMA_signal_3553), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2366_s_current_state_reg ( .D(
        new_AGEMA_signal_1922), .CK(clk), .Q(new_AGEMA_signal_3555), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2370_s_current_state_reg ( .D(
        new_AGEMA_signal_3558), .CK(clk), .Q(new_AGEMA_signal_3559), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2374_s_current_state_reg ( .D(
        new_AGEMA_signal_3562), .CK(clk), .Q(new_AGEMA_signal_3563), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2378_s_current_state_reg ( .D(
        new_AGEMA_signal_3566), .CK(clk), .Q(new_AGEMA_signal_3567), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2382_s_current_state_reg ( .D(
        new_AGEMA_signal_3570), .CK(clk), .Q(new_AGEMA_signal_3571), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2386_s_current_state_reg ( .D(
        new_AGEMA_signal_3574), .CK(clk), .Q(new_AGEMA_signal_3575), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2390_s_current_state_reg ( .D(
        new_AGEMA_signal_3578), .CK(clk), .Q(new_AGEMA_signal_3579), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2394_s_current_state_reg ( .D(
        new_AGEMA_signal_3582), .CK(clk), .Q(new_AGEMA_signal_3583), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2398_s_current_state_reg ( .D(
        new_AGEMA_signal_3586), .CK(clk), .Q(new_AGEMA_signal_3587), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2402_s_current_state_reg ( .D(
        new_AGEMA_signal_3590), .CK(clk), .Q(new_AGEMA_signal_3591), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2406_s_current_state_reg ( .D(
        new_AGEMA_signal_3594), .CK(clk), .Q(new_AGEMA_signal_3595), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2410_s_current_state_reg ( .D(
        new_AGEMA_signal_3598), .CK(clk), .Q(new_AGEMA_signal_3599), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2414_s_current_state_reg ( .D(
        new_AGEMA_signal_3602), .CK(clk), .Q(new_AGEMA_signal_3603), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2418_s_current_state_reg ( .D(
        new_AGEMA_signal_3606), .CK(clk), .Q(new_AGEMA_signal_3607), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2422_s_current_state_reg ( .D(
        new_AGEMA_signal_3610), .CK(clk), .Q(new_AGEMA_signal_3611), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2426_s_current_state_reg ( .D(
        new_AGEMA_signal_3614), .CK(clk), .Q(new_AGEMA_signal_3615), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2430_s_current_state_reg ( .D(
        new_AGEMA_signal_3618), .CK(clk), .Q(new_AGEMA_signal_3619), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2434_s_current_state_reg ( .D(
        new_AGEMA_signal_3622), .CK(clk), .Q(new_AGEMA_signal_3623), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2438_s_current_state_reg ( .D(
        new_AGEMA_signal_3626), .CK(clk), .Q(new_AGEMA_signal_3627), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2442_s_current_state_reg ( .D(
        new_AGEMA_signal_3630), .CK(clk), .Q(new_AGEMA_signal_3631), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2446_s_current_state_reg ( .D(
        new_AGEMA_signal_3634), .CK(clk), .Q(new_AGEMA_signal_3635), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2450_s_current_state_reg ( .D(
        new_AGEMA_signal_3638), .CK(clk), .Q(new_AGEMA_signal_3639), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2454_s_current_state_reg ( .D(
        new_AGEMA_signal_3642), .CK(clk), .Q(new_AGEMA_signal_3643), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2458_s_current_state_reg ( .D(
        new_AGEMA_signal_3646), .CK(clk), .Q(new_AGEMA_signal_3647), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2462_s_current_state_reg ( .D(
        new_AGEMA_signal_3650), .CK(clk), .Q(new_AGEMA_signal_3651), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2466_s_current_state_reg ( .D(
        new_AGEMA_signal_3654), .CK(clk), .Q(new_AGEMA_signal_3655), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2470_s_current_state_reg ( .D(
        new_AGEMA_signal_3658), .CK(clk), .Q(new_AGEMA_signal_3659), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2474_s_current_state_reg ( .D(
        new_AGEMA_signal_3662), .CK(clk), .Q(new_AGEMA_signal_3663), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2478_s_current_state_reg ( .D(
        new_AGEMA_signal_3666), .CK(clk), .Q(new_AGEMA_signal_3667), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2482_s_current_state_reg ( .D(
        new_AGEMA_signal_3670), .CK(clk), .Q(new_AGEMA_signal_3671), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2486_s_current_state_reg ( .D(
        new_AGEMA_signal_3674), .CK(clk), .Q(new_AGEMA_signal_3675), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2490_s_current_state_reg ( .D(
        new_AGEMA_signal_3678), .CK(clk), .Q(new_AGEMA_signal_3679), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2494_s_current_state_reg ( .D(
        new_AGEMA_signal_3682), .CK(clk), .Q(new_AGEMA_signal_3683), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2498_s_current_state_reg ( .D(
        new_AGEMA_signal_3686), .CK(clk), .Q(new_AGEMA_signal_3687), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2502_s_current_state_reg ( .D(
        new_AGEMA_signal_3690), .CK(clk), .Q(new_AGEMA_signal_3691), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2506_s_current_state_reg ( .D(
        new_AGEMA_signal_3694), .CK(clk), .Q(new_AGEMA_signal_3695), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2510_s_current_state_reg ( .D(
        new_AGEMA_signal_3698), .CK(clk), .Q(new_AGEMA_signal_3699), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2514_s_current_state_reg ( .D(
        new_AGEMA_signal_3702), .CK(clk), .Q(new_AGEMA_signal_3703), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2518_s_current_state_reg ( .D(
        new_AGEMA_signal_3706), .CK(clk), .Q(new_AGEMA_signal_3707), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2522_s_current_state_reg ( .D(
        new_AGEMA_signal_3710), .CK(clk), .Q(new_AGEMA_signal_3711), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2526_s_current_state_reg ( .D(
        new_AGEMA_signal_3714), .CK(clk), .Q(new_AGEMA_signal_3715), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2530_s_current_state_reg ( .D(
        new_AGEMA_signal_3718), .CK(clk), .Q(new_AGEMA_signal_3719), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2534_s_current_state_reg ( .D(
        new_AGEMA_signal_3722), .CK(clk), .Q(new_AGEMA_signal_3723), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2538_s_current_state_reg ( .D(
        new_AGEMA_signal_3726), .CK(clk), .Q(new_AGEMA_signal_3727), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2542_s_current_state_reg ( .D(
        new_AGEMA_signal_3730), .CK(clk), .Q(new_AGEMA_signal_3731), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2546_s_current_state_reg ( .D(
        new_AGEMA_signal_3734), .CK(clk), .Q(new_AGEMA_signal_3735), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2550_s_current_state_reg ( .D(
        new_AGEMA_signal_3738), .CK(clk), .Q(new_AGEMA_signal_3739), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2554_s_current_state_reg ( .D(
        new_AGEMA_signal_3742), .CK(clk), .Q(new_AGEMA_signal_3743), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2558_s_current_state_reg ( .D(
        new_AGEMA_signal_3746), .CK(clk), .Q(new_AGEMA_signal_3747), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2562_s_current_state_reg ( .D(
        new_AGEMA_signal_3750), .CK(clk), .Q(new_AGEMA_signal_3751), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2566_s_current_state_reg ( .D(
        new_AGEMA_signal_3754), .CK(clk), .Q(new_AGEMA_signal_3755), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2570_s_current_state_reg ( .D(
        new_AGEMA_signal_3758), .CK(clk), .Q(new_AGEMA_signal_3759), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2574_s_current_state_reg ( .D(
        new_AGEMA_signal_3762), .CK(clk), .Q(new_AGEMA_signal_3763), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2578_s_current_state_reg ( .D(
        new_AGEMA_signal_3766), .CK(clk), .Q(new_AGEMA_signal_3767), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2582_s_current_state_reg ( .D(
        new_AGEMA_signal_3770), .CK(clk), .Q(new_AGEMA_signal_3771), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2586_s_current_state_reg ( .D(
        new_AGEMA_signal_3774), .CK(clk), .Q(new_AGEMA_signal_3775), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2590_s_current_state_reg ( .D(
        new_AGEMA_signal_3778), .CK(clk), .Q(new_AGEMA_signal_3779), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2594_s_current_state_reg ( .D(
        new_AGEMA_signal_3782), .CK(clk), .Q(new_AGEMA_signal_3783), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2598_s_current_state_reg ( .D(
        new_AGEMA_signal_3786), .CK(clk), .Q(new_AGEMA_signal_3787), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2602_s_current_state_reg ( .D(
        new_AGEMA_signal_3790), .CK(clk), .Q(new_AGEMA_signal_3791), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2606_s_current_state_reg ( .D(
        new_AGEMA_signal_3794), .CK(clk), .Q(new_AGEMA_signal_3795), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2610_s_current_state_reg ( .D(
        new_AGEMA_signal_3798), .CK(clk), .Q(new_AGEMA_signal_3799), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2614_s_current_state_reg ( .D(
        new_AGEMA_signal_3802), .CK(clk), .Q(new_AGEMA_signal_3803), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2618_s_current_state_reg ( .D(
        new_AGEMA_signal_3806), .CK(clk), .Q(new_AGEMA_signal_3807), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2622_s_current_state_reg ( .D(
        new_AGEMA_signal_3810), .CK(clk), .Q(new_AGEMA_signal_3811), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2626_s_current_state_reg ( .D(
        new_AGEMA_signal_3814), .CK(clk), .Q(new_AGEMA_signal_3815), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2630_s_current_state_reg ( .D(
        new_AGEMA_signal_3818), .CK(clk), .Q(new_AGEMA_signal_3819), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2634_s_current_state_reg ( .D(
        new_AGEMA_signal_3822), .CK(clk), .Q(new_AGEMA_signal_3823), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2638_s_current_state_reg ( .D(
        new_AGEMA_signal_3826), .CK(clk), .Q(new_AGEMA_signal_3827), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2642_s_current_state_reg ( .D(
        new_AGEMA_signal_3830), .CK(clk), .Q(new_AGEMA_signal_3831), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2646_s_current_state_reg ( .D(
        new_AGEMA_signal_3834), .CK(clk), .Q(new_AGEMA_signal_3835), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2650_s_current_state_reg ( .D(
        new_AGEMA_signal_3838), .CK(clk), .Q(new_AGEMA_signal_3839), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2654_s_current_state_reg ( .D(
        new_AGEMA_signal_3842), .CK(clk), .Q(new_AGEMA_signal_3843), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2658_s_current_state_reg ( .D(
        new_AGEMA_signal_3846), .CK(clk), .Q(new_AGEMA_signal_3847), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2662_s_current_state_reg ( .D(
        new_AGEMA_signal_3850), .CK(clk), .Q(new_AGEMA_signal_3851), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2666_s_current_state_reg ( .D(
        new_AGEMA_signal_3854), .CK(clk), .Q(new_AGEMA_signal_3855), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2670_s_current_state_reg ( .D(
        new_AGEMA_signal_3858), .CK(clk), .Q(new_AGEMA_signal_3859), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2674_s_current_state_reg ( .D(
        new_AGEMA_signal_3862), .CK(clk), .Q(new_AGEMA_signal_3863), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2678_s_current_state_reg ( .D(
        new_AGEMA_signal_3866), .CK(clk), .Q(new_AGEMA_signal_3867), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2682_s_current_state_reg ( .D(
        new_AGEMA_signal_3870), .CK(clk), .Q(new_AGEMA_signal_3871), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2686_s_current_state_reg ( .D(
        new_AGEMA_signal_3874), .CK(clk), .Q(new_AGEMA_signal_3875), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2690_s_current_state_reg ( .D(
        new_AGEMA_signal_3878), .CK(clk), .Q(new_AGEMA_signal_3879), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2694_s_current_state_reg ( .D(
        new_AGEMA_signal_3882), .CK(clk), .Q(new_AGEMA_signal_3883), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2698_s_current_state_reg ( .D(
        new_AGEMA_signal_3886), .CK(clk), .Q(new_AGEMA_signal_3887), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2702_s_current_state_reg ( .D(
        new_AGEMA_signal_3890), .CK(clk), .Q(new_AGEMA_signal_3891), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2706_s_current_state_reg ( .D(
        new_AGEMA_signal_3894), .CK(clk), .Q(new_AGEMA_signal_3895), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2710_s_current_state_reg ( .D(
        new_AGEMA_signal_3898), .CK(clk), .Q(new_AGEMA_signal_3899), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2714_s_current_state_reg ( .D(
        new_AGEMA_signal_3902), .CK(clk), .Q(new_AGEMA_signal_3903), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2718_s_current_state_reg ( .D(
        new_AGEMA_signal_3906), .CK(clk), .Q(new_AGEMA_signal_3907), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2722_s_current_state_reg ( .D(
        new_AGEMA_signal_3910), .CK(clk), .Q(new_AGEMA_signal_3911), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2726_s_current_state_reg ( .D(
        new_AGEMA_signal_3914), .CK(clk), .Q(new_AGEMA_signal_3915), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2730_s_current_state_reg ( .D(
        new_AGEMA_signal_3918), .CK(clk), .Q(new_AGEMA_signal_3919), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2734_s_current_state_reg ( .D(
        new_AGEMA_signal_3922), .CK(clk), .Q(new_AGEMA_signal_3923), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2738_s_current_state_reg ( .D(
        new_AGEMA_signal_3926), .CK(clk), .Q(new_AGEMA_signal_3927), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2742_s_current_state_reg ( .D(
        new_AGEMA_signal_3930), .CK(clk), .Q(new_AGEMA_signal_3931), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2746_s_current_state_reg ( .D(
        new_AGEMA_signal_3934), .CK(clk), .Q(new_AGEMA_signal_3935), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2750_s_current_state_reg ( .D(
        new_AGEMA_signal_3938), .CK(clk), .Q(new_AGEMA_signal_3939), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2754_s_current_state_reg ( .D(
        new_AGEMA_signal_3942), .CK(clk), .Q(new_AGEMA_signal_3943), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2758_s_current_state_reg ( .D(
        new_AGEMA_signal_3946), .CK(clk), .Q(new_AGEMA_signal_3947), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2762_s_current_state_reg ( .D(
        new_AGEMA_signal_3950), .CK(clk), .Q(new_AGEMA_signal_3951), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2766_s_current_state_reg ( .D(
        new_AGEMA_signal_3954), .CK(clk), .Q(new_AGEMA_signal_3955), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2770_s_current_state_reg ( .D(
        new_AGEMA_signal_3958), .CK(clk), .Q(new_AGEMA_signal_3959), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2774_s_current_state_reg ( .D(
        new_AGEMA_signal_3962), .CK(clk), .Q(new_AGEMA_signal_3963), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2778_s_current_state_reg ( .D(
        new_AGEMA_signal_3966), .CK(clk), .Q(new_AGEMA_signal_3967), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2782_s_current_state_reg ( .D(
        new_AGEMA_signal_3970), .CK(clk), .Q(new_AGEMA_signal_3971), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2786_s_current_state_reg ( .D(
        new_AGEMA_signal_3974), .CK(clk), .Q(new_AGEMA_signal_3975), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2790_s_current_state_reg ( .D(
        new_AGEMA_signal_3978), .CK(clk), .Q(new_AGEMA_signal_3979), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2794_s_current_state_reg ( .D(
        new_AGEMA_signal_3982), .CK(clk), .Q(new_AGEMA_signal_3983), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2798_s_current_state_reg ( .D(
        new_AGEMA_signal_3986), .CK(clk), .Q(new_AGEMA_signal_3987), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2802_s_current_state_reg ( .D(
        new_AGEMA_signal_3990), .CK(clk), .Q(new_AGEMA_signal_3991), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2806_s_current_state_reg ( .D(
        new_AGEMA_signal_3994), .CK(clk), .Q(new_AGEMA_signal_3995), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2810_s_current_state_reg ( .D(
        new_AGEMA_signal_3998), .CK(clk), .Q(new_AGEMA_signal_3999), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2814_s_current_state_reg ( .D(
        new_AGEMA_signal_4002), .CK(clk), .Q(new_AGEMA_signal_4003), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2818_s_current_state_reg ( .D(
        new_AGEMA_signal_4006), .CK(clk), .Q(new_AGEMA_signal_4007), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2822_s_current_state_reg ( .D(
        new_AGEMA_signal_4010), .CK(clk), .Q(new_AGEMA_signal_4011), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2826_s_current_state_reg ( .D(
        new_AGEMA_signal_4014), .CK(clk), .Q(new_AGEMA_signal_4015), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2830_s_current_state_reg ( .D(
        new_AGEMA_signal_4018), .CK(clk), .Q(new_AGEMA_signal_4019), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2834_s_current_state_reg ( .D(
        new_AGEMA_signal_4022), .CK(clk), .Q(new_AGEMA_signal_4023), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2838_s_current_state_reg ( .D(
        new_AGEMA_signal_4026), .CK(clk), .Q(new_AGEMA_signal_4027), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2842_s_current_state_reg ( .D(
        new_AGEMA_signal_4030), .CK(clk), .Q(new_AGEMA_signal_4031), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2846_s_current_state_reg ( .D(
        new_AGEMA_signal_4034), .CK(clk), .Q(new_AGEMA_signal_4035), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2850_s_current_state_reg ( .D(
        new_AGEMA_signal_4038), .CK(clk), .Q(new_AGEMA_signal_4039), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2854_s_current_state_reg ( .D(
        new_AGEMA_signal_4042), .CK(clk), .Q(new_AGEMA_signal_4043), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2858_s_current_state_reg ( .D(
        new_AGEMA_signal_4046), .CK(clk), .Q(new_AGEMA_signal_4047), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2862_s_current_state_reg ( .D(
        new_AGEMA_signal_4050), .CK(clk), .Q(new_AGEMA_signal_4051), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2866_s_current_state_reg ( .D(
        new_AGEMA_signal_4054), .CK(clk), .Q(new_AGEMA_signal_4055), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2870_s_current_state_reg ( .D(
        new_AGEMA_signal_4058), .CK(clk), .Q(new_AGEMA_signal_4059), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2874_s_current_state_reg ( .D(
        new_AGEMA_signal_4062), .CK(clk), .Q(new_AGEMA_signal_4063), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2878_s_current_state_reg ( .D(
        new_AGEMA_signal_4066), .CK(clk), .Q(new_AGEMA_signal_4067), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2882_s_current_state_reg ( .D(
        new_AGEMA_signal_4070), .CK(clk), .Q(new_AGEMA_signal_4071), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2886_s_current_state_reg ( .D(
        new_AGEMA_signal_4074), .CK(clk), .Q(new_AGEMA_signal_4075), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2890_s_current_state_reg ( .D(
        new_AGEMA_signal_4078), .CK(clk), .Q(new_AGEMA_signal_4079), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2894_s_current_state_reg ( .D(
        new_AGEMA_signal_4082), .CK(clk), .Q(new_AGEMA_signal_4083), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2898_s_current_state_reg ( .D(
        new_AGEMA_signal_4086), .CK(clk), .Q(new_AGEMA_signal_4087), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2902_s_current_state_reg ( .D(
        new_AGEMA_signal_4090), .CK(clk), .Q(new_AGEMA_signal_4091), .QN() );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_0_U1 ( .A(MCOutput[0]), .B(
        new_AGEMA_signal_2648), .S(n35), .Z(StateRegInput[0]) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2027), .B(
        new_AGEMA_signal_2652), .S(n35), .Z(new_AGEMA_signal_2036) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_0_U1 ( .A(MCOutput[1]), .B(
        new_AGEMA_signal_2656), .S(n36), .Z(StateRegInput[1]) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2073), .B(
        new_AGEMA_signal_2660), .S(n36), .Z(new_AGEMA_signal_2079) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_0_U1 ( .A(MCOutput[4]), .B(
        new_AGEMA_signal_2664), .S(new_AGEMA_signal_2644), .Z(StateRegInput[4]) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2029), .B(
        new_AGEMA_signal_2668), .S(new_AGEMA_signal_2644), .Z(
        new_AGEMA_signal_2038) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_0_U1 ( .A(MCOutput[5]), .B(
        new_AGEMA_signal_2672), .S(new_AGEMA_signal_2644), .Z(StateRegInput[5]) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2074), .B(
        new_AGEMA_signal_2676), .S(new_AGEMA_signal_2644), .Z(
        new_AGEMA_signal_2081) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_0_U1 ( .A(MCOutput[8]), .B(
        new_AGEMA_signal_2680), .S(new_AGEMA_signal_2644), .Z(StateRegInput[8]) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2031), .B(
        new_AGEMA_signal_2684), .S(new_AGEMA_signal_2644), .Z(
        new_AGEMA_signal_2040) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_0_U1 ( .A(MCOutput[9]), .B(
        new_AGEMA_signal_2688), .S(new_AGEMA_signal_2644), .Z(StateRegInput[9]) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2075), .B(
        new_AGEMA_signal_2692), .S(new_AGEMA_signal_2644), .Z(
        new_AGEMA_signal_2083) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_0_U1 ( .A(MCOutput[12]), .B(
        new_AGEMA_signal_2696), .S(new_AGEMA_signal_2644), .Z(
        StateRegInput[12]) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2108), .B(
        new_AGEMA_signal_2700), .S(new_AGEMA_signal_2644), .Z(
        new_AGEMA_signal_2111) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_0_U1 ( .A(MCOutput[13]), .B(
        new_AGEMA_signal_2704), .S(n34), .Z(StateRegInput[13]) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2118), .B(
        new_AGEMA_signal_2708), .S(n34), .Z(new_AGEMA_signal_2120) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_0_U1 ( .A(MCOutput[16]), .B(
        new_AGEMA_signal_2712), .S(n34), .Z(StateRegInput[16]) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2019), .B(
        new_AGEMA_signal_2716), .S(n34), .Z(new_AGEMA_signal_2044) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_0_U1 ( .A(MCOutput[17]), .B(
        new_AGEMA_signal_2720), .S(n34), .Z(StateRegInput[17]) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2068), .B(
        new_AGEMA_signal_2724), .S(n34), .Z(new_AGEMA_signal_2087) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_0_U1 ( .A(MCOutput[20]), .B(
        new_AGEMA_signal_2728), .S(n34), .Z(StateRegInput[20]) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2021), .B(
        new_AGEMA_signal_2732), .S(n34), .Z(new_AGEMA_signal_2046) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_0_U1 ( .A(MCOutput[21]), .B(
        new_AGEMA_signal_2736), .S(n34), .Z(StateRegInput[21]) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2069), .B(
        new_AGEMA_signal_2740), .S(n34), .Z(new_AGEMA_signal_2089) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_0_U1 ( .A(MCOutput[24]), .B(
        new_AGEMA_signal_2744), .S(n34), .Z(StateRegInput[24]) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2106), .B(
        new_AGEMA_signal_2748), .S(n34), .Z(new_AGEMA_signal_2113) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_0_U1 ( .A(MCOutput[25]), .B(
        new_AGEMA_signal_2752), .S(n34), .Z(StateRegInput[25]) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2117), .B(
        new_AGEMA_signal_2756), .S(n34), .Z(new_AGEMA_signal_2122) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_0_U1 ( .A(MCOutput[28]), .B(
        new_AGEMA_signal_2760), .S(n35), .Z(StateRegInput[28]) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2025), .B(
        new_AGEMA_signal_2764), .S(n35), .Z(new_AGEMA_signal_2050) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_0_U1 ( .A(MCOutput[29]), .B(
        new_AGEMA_signal_2768), .S(n35), .Z(StateRegInput[29]) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2072), .B(
        new_AGEMA_signal_2772), .S(n35), .Z(new_AGEMA_signal_2093) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_0_U1 ( .A(MCOutput[32]), .B(
        new_AGEMA_signal_2776), .S(n35), .Z(StateRegInput[32]) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1892), .B(
        new_AGEMA_signal_2780), .S(n35), .Z(new_AGEMA_signal_1934) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_0_U1 ( .A(MCOutput[33]), .B(
        new_AGEMA_signal_2784), .S(n35), .Z(StateRegInput[33]) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1954), .B(
        new_AGEMA_signal_2788), .S(n35), .Z(new_AGEMA_signal_1994) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_0_U1 ( .A(MCOutput[36]), .B(
        new_AGEMA_signal_2792), .S(n35), .Z(StateRegInput[36]) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1894), .B(
        new_AGEMA_signal_2796), .S(n35), .Z(new_AGEMA_signal_1936) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_0_U1 ( .A(MCOutput[37]), .B(
        new_AGEMA_signal_2800), .S(n35), .Z(StateRegInput[37]) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1955), .B(
        new_AGEMA_signal_2804), .S(n35), .Z(new_AGEMA_signal_1996) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_0_U1 ( .A(MCOutput[40]), .B(
        new_AGEMA_signal_2808), .S(n35), .Z(StateRegInput[40]) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1896), .B(
        new_AGEMA_signal_2812), .S(n35), .Z(new_AGEMA_signal_1938) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_0_U1 ( .A(MCOutput[41]), .B(
        new_AGEMA_signal_2816), .S(n36), .Z(StateRegInput[41]) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1956), .B(
        new_AGEMA_signal_2820), .S(n36), .Z(new_AGEMA_signal_1998) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_0_U1 ( .A(MCOutput[44]), .B(
        new_AGEMA_signal_2824), .S(n36), .Z(StateRegInput[44]) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2009), .B(
        new_AGEMA_signal_2828), .S(n36), .Z(new_AGEMA_signal_2052) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_0_U1 ( .A(MCOutput[45]), .B(
        new_AGEMA_signal_2832), .S(n36), .Z(StateRegInput[45]) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2062), .B(
        new_AGEMA_signal_2836), .S(n36), .Z(new_AGEMA_signal_2095) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_0_U1 ( .A(MCOutput[48]), .B(
        new_AGEMA_signal_2840), .S(n36), .Z(StateRegInput[48]) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2011), .B(
        new_AGEMA_signal_2844), .S(n36), .Z(new_AGEMA_signal_2054) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_0_U1 ( .A(MCOutput[49]), .B(
        new_AGEMA_signal_2848), .S(n36), .Z(StateRegInput[49]) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2063), .B(
        new_AGEMA_signal_2852), .S(n36), .Z(new_AGEMA_signal_2097) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_0_U1 ( .A(MCOutput[52]), .B(
        new_AGEMA_signal_2856), .S(n36), .Z(StateRegInput[52]) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2013), .B(
        new_AGEMA_signal_2860), .S(n36), .Z(new_AGEMA_signal_2056) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_0_U1 ( .A(MCOutput[53]), .B(
        new_AGEMA_signal_2864), .S(n36), .Z(StateRegInput[53]) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2064), .B(
        new_AGEMA_signal_2868), .S(n36), .Z(new_AGEMA_signal_2099) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_0_U1 ( .A(MCOutput[56]), .B(
        new_AGEMA_signal_2872), .S(new_AGEMA_signal_2644), .Z(
        StateRegInput[56]) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2015), .B(
        new_AGEMA_signal_2876), .S(new_AGEMA_signal_2644), .Z(
        new_AGEMA_signal_2058) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_0_U1 ( .A(MCOutput[57]), .B(
        new_AGEMA_signal_2880), .S(new_AGEMA_signal_2644), .Z(
        StateRegInput[57]) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2065), .B(
        new_AGEMA_signal_2884), .S(new_AGEMA_signal_2644), .Z(
        new_AGEMA_signal_2101) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_0_U1 ( .A(MCOutput[60]), .B(
        new_AGEMA_signal_2888), .S(new_AGEMA_signal_2644), .Z(
        StateRegInput[60]) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2104), .B(
        new_AGEMA_signal_2892), .S(new_AGEMA_signal_2644), .Z(
        new_AGEMA_signal_2115) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_0_U1 ( .A(MCOutput[61]), .B(
        new_AGEMA_signal_2896), .S(new_AGEMA_signal_2644), .Z(
        StateRegInput[61]) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2116), .B(
        new_AGEMA_signal_2900), .S(new_AGEMA_signal_2644), .Z(
        new_AGEMA_signal_2124) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U14 ( .A(Fresh[32]), .B(
        SubCellInst_SboxInst_0_Q2), .Z(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U13 ( .A(Fresh[32]), .B(
        new_AGEMA_signal_1596), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U10 ( .A1(new_AGEMA_signal_2904), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U9 ( .A1(new_AGEMA_signal_2902), .A2(
        SubCellInst_SboxInst_0_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U8 ( .A(Fresh[32]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U7 ( .A1(new_AGEMA_signal_1596), .A2(
        new_AGEMA_signal_2904), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_0_Q2), 
        .A2(new_AGEMA_signal_2902), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n8), .B(
        SubCellInst_SboxInst_0_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1661) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n7), .B(
        SubCellInst_SboxInst_0_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_0_T1) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2902), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2904), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_T1), .B(new_AGEMA_signal_2906), .Z(
        SubCellInst_SboxInst_0_L0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1661), 
        .B(new_AGEMA_signal_2908), .Z(new_AGEMA_signal_1725) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U14 ( .A(Fresh[33]), .B(
        SubCellInst_SboxInst_0_Q7), .Z(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U13 ( .A(Fresh[33]), .B(
        new_AGEMA_signal_1597), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U10 ( .A1(new_AGEMA_signal_2912), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U9 ( .A1(new_AGEMA_signal_2910), .A2(
        SubCellInst_SboxInst_0_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U8 ( .A(Fresh[33]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U7 ( .A1(new_AGEMA_signal_1597), .A2(
        new_AGEMA_signal_2912), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_0_Q7), 
        .A2(new_AGEMA_signal_2910), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n8), .B(
        SubCellInst_SboxInst_0_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1662) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n7), .B(
        SubCellInst_SboxInst_0_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_0_T3) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2910), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2912), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L0), .B(new_AGEMA_signal_2916), .Z(
        SubCellInst_SboxInst_0_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1725), 
        .B(new_AGEMA_signal_2920), .Z(new_AGEMA_signal_1768) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L0), .B(SubCellInst_SboxInst_0_T3), .Z(
        ShiftRowsOutput[4]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1725), 
        .B(new_AGEMA_signal_1662), .Z(new_AGEMA_signal_1769) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_2922), .B(SubCellInst_SboxInst_0_YY_3), .ZN(ShiftRowsOutput[5]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2924), .B(new_AGEMA_signal_1768), .Z(new_AGEMA_signal_1826) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U14 ( .A(Fresh[34]), .B(
        SubCellInst_SboxInst_1_Q2), .Z(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U13 ( .A(Fresh[34]), .B(
        new_AGEMA_signal_1600), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U10 ( .A1(new_AGEMA_signal_2928), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U9 ( .A1(new_AGEMA_signal_2926), .A2(
        SubCellInst_SboxInst_1_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U8 ( .A(Fresh[34]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U7 ( .A1(new_AGEMA_signal_1600), .A2(
        new_AGEMA_signal_2928), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_1_Q2), 
        .A2(new_AGEMA_signal_2926), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n8), .B(
        SubCellInst_SboxInst_1_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1665) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n7), .B(
        SubCellInst_SboxInst_1_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_1_T1) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2926), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2928), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_T1), .B(new_AGEMA_signal_2930), .Z(
        SubCellInst_SboxInst_1_L0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1665), 
        .B(new_AGEMA_signal_2932), .Z(new_AGEMA_signal_1727) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U14 ( .A(Fresh[35]), .B(
        SubCellInst_SboxInst_1_Q7), .Z(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U13 ( .A(Fresh[35]), .B(
        new_AGEMA_signal_1601), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U10 ( .A1(new_AGEMA_signal_2936), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U9 ( .A1(new_AGEMA_signal_2934), .A2(
        SubCellInst_SboxInst_1_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U8 ( .A(Fresh[35]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U7 ( .A1(new_AGEMA_signal_1601), .A2(
        new_AGEMA_signal_2936), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_1_Q7), 
        .A2(new_AGEMA_signal_2934), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n8), .B(
        SubCellInst_SboxInst_1_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1666) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n7), .B(
        SubCellInst_SboxInst_1_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_1_T3) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2934), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2936), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L0), .B(new_AGEMA_signal_2940), .Z(
        SubCellInst_SboxInst_1_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1727), 
        .B(new_AGEMA_signal_2944), .Z(new_AGEMA_signal_1770) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L0), .B(SubCellInst_SboxInst_1_T3), .Z(
        ShiftRowsOutput[8]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1727), 
        .B(new_AGEMA_signal_1666), .Z(new_AGEMA_signal_1771) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_2946), .B(SubCellInst_SboxInst_1_YY_3), .ZN(ShiftRowsOutput[9]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2948), .B(new_AGEMA_signal_1770), .Z(new_AGEMA_signal_1827) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U14 ( .A(Fresh[36]), .B(
        SubCellInst_SboxInst_2_Q2), .Z(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U13 ( .A(Fresh[36]), .B(
        new_AGEMA_signal_1604), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U10 ( .A1(new_AGEMA_signal_2952), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U9 ( .A1(new_AGEMA_signal_2950), .A2(
        SubCellInst_SboxInst_2_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U8 ( .A(Fresh[36]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U7 ( .A1(new_AGEMA_signal_1604), .A2(
        new_AGEMA_signal_2952), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_2_Q2), 
        .A2(new_AGEMA_signal_2950), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n8), .B(
        SubCellInst_SboxInst_2_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1669) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n7), .B(
        SubCellInst_SboxInst_2_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_2_T1) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2950), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2952), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_T1), .B(new_AGEMA_signal_2954), .Z(
        SubCellInst_SboxInst_2_L0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1669), 
        .B(new_AGEMA_signal_2956), .Z(new_AGEMA_signal_1729) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U14 ( .A(Fresh[37]), .B(
        SubCellInst_SboxInst_2_Q7), .Z(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U13 ( .A(Fresh[37]), .B(
        new_AGEMA_signal_1605), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U10 ( .A1(new_AGEMA_signal_2960), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U9 ( .A1(new_AGEMA_signal_2958), .A2(
        SubCellInst_SboxInst_2_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U8 ( .A(Fresh[37]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U7 ( .A1(new_AGEMA_signal_1605), .A2(
        new_AGEMA_signal_2960), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_2_Q7), 
        .A2(new_AGEMA_signal_2958), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n8), .B(
        SubCellInst_SboxInst_2_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1670) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n7), .B(
        SubCellInst_SboxInst_2_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_2_T3) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2958), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2960), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L0), .B(new_AGEMA_signal_2964), .Z(
        SubCellInst_SboxInst_2_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1729), 
        .B(new_AGEMA_signal_2968), .Z(new_AGEMA_signal_1772) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L0), .B(SubCellInst_SboxInst_2_T3), .Z(
        ShiftRowsOutput[12]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1729), 
        .B(new_AGEMA_signal_1670), .Z(new_AGEMA_signal_1773) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_2970), .B(SubCellInst_SboxInst_2_YY_3), .ZN(ShiftRowsOutput[13]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2972), .B(new_AGEMA_signal_1772), .Z(new_AGEMA_signal_1828) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U14 ( .A(Fresh[38]), .B(
        SubCellInst_SboxInst_3_Q2), .Z(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U13 ( .A(Fresh[38]), .B(
        new_AGEMA_signal_1608), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U10 ( .A1(new_AGEMA_signal_2976), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U9 ( .A1(new_AGEMA_signal_2974), .A2(
        SubCellInst_SboxInst_3_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U8 ( .A(Fresh[38]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U7 ( .A1(new_AGEMA_signal_1608), .A2(
        new_AGEMA_signal_2976), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_3_Q2), 
        .A2(new_AGEMA_signal_2974), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n8), .B(
        SubCellInst_SboxInst_3_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1673) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n7), .B(
        SubCellInst_SboxInst_3_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_3_T1) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2974), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2976), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_T1), .B(new_AGEMA_signal_2978), .Z(
        SubCellInst_SboxInst_3_L0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1673), 
        .B(new_AGEMA_signal_2980), .Z(new_AGEMA_signal_1731) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U14 ( .A(Fresh[39]), .B(
        SubCellInst_SboxInst_3_Q7), .Z(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U13 ( .A(Fresh[39]), .B(
        new_AGEMA_signal_1609), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U10 ( .A1(new_AGEMA_signal_2984), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U9 ( .A1(new_AGEMA_signal_2982), .A2(
        SubCellInst_SboxInst_3_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U8 ( .A(Fresh[39]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U7 ( .A1(new_AGEMA_signal_1609), .A2(
        new_AGEMA_signal_2984), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_3_Q7), 
        .A2(new_AGEMA_signal_2982), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n8), .B(
        SubCellInst_SboxInst_3_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1674) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n7), .B(
        SubCellInst_SboxInst_3_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_3_T3) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2982), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2984), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L0), .B(new_AGEMA_signal_2988), .Z(
        SubCellInst_SboxInst_3_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1731), 
        .B(new_AGEMA_signal_2992), .Z(new_AGEMA_signal_1774) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L0), .B(SubCellInst_SboxInst_3_T3), .Z(
        ShiftRowsOutput[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1731), 
        .B(new_AGEMA_signal_1674), .Z(new_AGEMA_signal_1775) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_2994), .B(SubCellInst_SboxInst_3_YY_3), .ZN(ShiftRowsOutput[1]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2996), .B(new_AGEMA_signal_1774), .Z(new_AGEMA_signal_1829) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U14 ( .A(Fresh[40]), .B(
        SubCellInst_SboxInst_4_Q2), .Z(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U13 ( .A(Fresh[40]), .B(
        new_AGEMA_signal_1612), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U10 ( .A1(new_AGEMA_signal_3000), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U9 ( .A1(new_AGEMA_signal_2998), .A2(
        SubCellInst_SboxInst_4_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U8 ( .A(Fresh[40]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U7 ( .A1(new_AGEMA_signal_1612), .A2(
        new_AGEMA_signal_3000), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_4_Q2), 
        .A2(new_AGEMA_signal_2998), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n8), .B(
        SubCellInst_SboxInst_4_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1677) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n7), .B(
        SubCellInst_SboxInst_4_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_4_T1) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2998), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3000), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_T1), .B(new_AGEMA_signal_3002), .Z(
        SubCellInst_SboxInst_4_L0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1677), 
        .B(new_AGEMA_signal_3004), .Z(new_AGEMA_signal_1733) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U14 ( .A(Fresh[41]), .B(
        SubCellInst_SboxInst_4_Q7), .Z(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U13 ( .A(Fresh[41]), .B(
        new_AGEMA_signal_1613), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U10 ( .A1(new_AGEMA_signal_3008), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U9 ( .A1(new_AGEMA_signal_3006), .A2(
        SubCellInst_SboxInst_4_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U8 ( .A(Fresh[41]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U7 ( .A1(new_AGEMA_signal_1613), .A2(
        new_AGEMA_signal_3008), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_4_Q7), 
        .A2(new_AGEMA_signal_3006), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n8), .B(
        SubCellInst_SboxInst_4_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1678) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n7), .B(
        SubCellInst_SboxInst_4_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_4_T3) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3006), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3008), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L0), .B(new_AGEMA_signal_3012), .Z(
        SubCellInst_SboxInst_4_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1733), 
        .B(new_AGEMA_signal_3016), .Z(new_AGEMA_signal_1776) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L0), .B(SubCellInst_SboxInst_4_T3), .Z(
        ShiftRowsOutput[24]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1733), 
        .B(new_AGEMA_signal_1678), .Z(new_AGEMA_signal_1777) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_3018), .B(SubCellInst_SboxInst_4_YY_3), .ZN(ShiftRowsOutput[25]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3020), .B(new_AGEMA_signal_1776), .Z(new_AGEMA_signal_1830) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U14 ( .A(Fresh[42]), .B(
        SubCellInst_SboxInst_5_Q2), .Z(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U13 ( .A(Fresh[42]), .B(
        new_AGEMA_signal_1616), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U10 ( .A1(new_AGEMA_signal_3024), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U9 ( .A1(new_AGEMA_signal_3022), .A2(
        SubCellInst_SboxInst_5_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U8 ( .A(Fresh[42]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U7 ( .A1(new_AGEMA_signal_1616), .A2(
        new_AGEMA_signal_3024), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_5_Q2), 
        .A2(new_AGEMA_signal_3022), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n8), .B(
        SubCellInst_SboxInst_5_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1681) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n7), .B(
        SubCellInst_SboxInst_5_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_5_T1) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3022), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3024), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_T1), .B(new_AGEMA_signal_3026), .Z(
        SubCellInst_SboxInst_5_L0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1681), 
        .B(new_AGEMA_signal_3028), .Z(new_AGEMA_signal_1735) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U14 ( .A(Fresh[43]), .B(
        SubCellInst_SboxInst_5_Q7), .Z(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U13 ( .A(Fresh[43]), .B(
        new_AGEMA_signal_1617), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U10 ( .A1(new_AGEMA_signal_3032), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U9 ( .A1(new_AGEMA_signal_3030), .A2(
        SubCellInst_SboxInst_5_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U8 ( .A(Fresh[43]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U7 ( .A1(new_AGEMA_signal_1617), .A2(
        new_AGEMA_signal_3032), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_5_Q7), 
        .A2(new_AGEMA_signal_3030), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n8), .B(
        SubCellInst_SboxInst_5_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1682) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n7), .B(
        SubCellInst_SboxInst_5_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_5_T3) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3030), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3032), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L0), .B(new_AGEMA_signal_3036), .Z(
        SubCellInst_SboxInst_5_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1735), 
        .B(new_AGEMA_signal_3040), .Z(new_AGEMA_signal_1778) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L0), .B(SubCellInst_SboxInst_5_T3), .Z(
        ShiftRowsOutput[28]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1735), 
        .B(new_AGEMA_signal_1682), .Z(new_AGEMA_signal_1779) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_3042), .B(SubCellInst_SboxInst_5_YY_3), .ZN(ShiftRowsOutput[29]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3044), .B(new_AGEMA_signal_1778), .Z(new_AGEMA_signal_1831) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U14 ( .A(Fresh[44]), .B(
        SubCellInst_SboxInst_6_Q2), .Z(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U13 ( .A(Fresh[44]), .B(
        new_AGEMA_signal_1620), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U10 ( .A1(new_AGEMA_signal_3048), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U9 ( .A1(new_AGEMA_signal_3046), .A2(
        SubCellInst_SboxInst_6_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U8 ( .A(Fresh[44]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U7 ( .A1(new_AGEMA_signal_1620), .A2(
        new_AGEMA_signal_3048), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_6_Q2), 
        .A2(new_AGEMA_signal_3046), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n8), .B(
        SubCellInst_SboxInst_6_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1685) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n7), .B(
        SubCellInst_SboxInst_6_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_6_T1) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3046), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3048), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_T1), .B(new_AGEMA_signal_3050), .Z(
        SubCellInst_SboxInst_6_L0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1685), 
        .B(new_AGEMA_signal_3052), .Z(new_AGEMA_signal_1737) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U14 ( .A(Fresh[45]), .B(
        SubCellInst_SboxInst_6_Q7), .Z(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U13 ( .A(Fresh[45]), .B(
        new_AGEMA_signal_1621), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U10 ( .A1(new_AGEMA_signal_3056), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U9 ( .A1(new_AGEMA_signal_3054), .A2(
        SubCellInst_SboxInst_6_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U8 ( .A(Fresh[45]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U7 ( .A1(new_AGEMA_signal_1621), .A2(
        new_AGEMA_signal_3056), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_6_Q7), 
        .A2(new_AGEMA_signal_3054), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n8), .B(
        SubCellInst_SboxInst_6_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1686) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n7), .B(
        SubCellInst_SboxInst_6_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_6_T3) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3054), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3056), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L0), .B(new_AGEMA_signal_3060), .Z(
        SubCellInst_SboxInst_6_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1737), 
        .B(new_AGEMA_signal_3064), .Z(new_AGEMA_signal_1780) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L0), .B(SubCellInst_SboxInst_6_T3), .Z(
        ShiftRowsOutput[16]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1737), 
        .B(new_AGEMA_signal_1686), .Z(new_AGEMA_signal_1781) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_3066), .B(SubCellInst_SboxInst_6_YY_3), .ZN(ShiftRowsOutput[17]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3068), .B(new_AGEMA_signal_1780), .Z(new_AGEMA_signal_1832) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U14 ( .A(Fresh[46]), .B(
        SubCellInst_SboxInst_7_Q2), .Z(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U13 ( .A(Fresh[46]), .B(
        new_AGEMA_signal_1624), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U10 ( .A1(new_AGEMA_signal_3072), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U9 ( .A1(new_AGEMA_signal_3070), .A2(
        SubCellInst_SboxInst_7_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U8 ( .A(Fresh[46]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U7 ( .A1(new_AGEMA_signal_1624), .A2(
        new_AGEMA_signal_3072), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_7_Q2), 
        .A2(new_AGEMA_signal_3070), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n8), .B(
        SubCellInst_SboxInst_7_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1689) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n7), .B(
        SubCellInst_SboxInst_7_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_7_T1) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3070), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3072), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_T1), .B(new_AGEMA_signal_3074), .Z(
        SubCellInst_SboxInst_7_L0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1689), 
        .B(new_AGEMA_signal_3076), .Z(new_AGEMA_signal_1739) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U14 ( .A(Fresh[47]), .B(
        SubCellInst_SboxInst_7_Q7), .Z(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U13 ( .A(Fresh[47]), .B(
        new_AGEMA_signal_1625), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U10 ( .A1(new_AGEMA_signal_3080), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U9 ( .A1(new_AGEMA_signal_3078), .A2(
        SubCellInst_SboxInst_7_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U8 ( .A(Fresh[47]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U7 ( .A1(new_AGEMA_signal_1625), .A2(
        new_AGEMA_signal_3080), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_7_Q7), 
        .A2(new_AGEMA_signal_3078), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n8), .B(
        SubCellInst_SboxInst_7_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1690) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n7), .B(
        SubCellInst_SboxInst_7_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_7_T3) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3078), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3080), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L0), .B(new_AGEMA_signal_3084), .Z(
        SubCellInst_SboxInst_7_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1739), 
        .B(new_AGEMA_signal_3088), .Z(new_AGEMA_signal_1782) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L0), .B(SubCellInst_SboxInst_7_T3), .Z(
        ShiftRowsOutput[20]) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1739), 
        .B(new_AGEMA_signal_1690), .Z(new_AGEMA_signal_1783) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_3090), .B(SubCellInst_SboxInst_7_YY_3), .ZN(SubCellOutput_29) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3092), .B(new_AGEMA_signal_1782), .Z(new_AGEMA_signal_1879) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U14 ( .A(Fresh[48]), .B(
        SubCellInst_SboxInst_8_Q2), .Z(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U13 ( .A(Fresh[48]), .B(
        new_AGEMA_signal_1628), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U10 ( .A1(new_AGEMA_signal_3096), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U9 ( .A1(new_AGEMA_signal_3094), .A2(
        SubCellInst_SboxInst_8_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U8 ( .A(Fresh[48]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U7 ( .A1(new_AGEMA_signal_1628), .A2(
        new_AGEMA_signal_3096), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_8_Q2), 
        .A2(new_AGEMA_signal_3094), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n8), .B(
        SubCellInst_SboxInst_8_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1693) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n7), .B(
        SubCellInst_SboxInst_8_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_8_T1) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3094), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3096), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_T1), .B(new_AGEMA_signal_3098), .Z(
        SubCellInst_SboxInst_8_L0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1693), 
        .B(new_AGEMA_signal_3100), .Z(new_AGEMA_signal_1741) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U14 ( .A(Fresh[49]), .B(
        SubCellInst_SboxInst_8_Q7), .Z(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U13 ( .A(Fresh[49]), .B(
        new_AGEMA_signal_1629), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U10 ( .A1(new_AGEMA_signal_3104), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U9 ( .A1(new_AGEMA_signal_3102), .A2(
        SubCellInst_SboxInst_8_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U8 ( .A(Fresh[49]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U7 ( .A1(new_AGEMA_signal_1629), .A2(
        new_AGEMA_signal_3104), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_8_Q7), 
        .A2(new_AGEMA_signal_3102), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n8), .B(
        SubCellInst_SboxInst_8_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1694) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n7), .B(
        SubCellInst_SboxInst_8_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_8_T3) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3102), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3104), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L0), .B(new_AGEMA_signal_3108), .Z(
        SubCellInst_SboxInst_8_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1741), 
        .B(new_AGEMA_signal_3112), .Z(new_AGEMA_signal_1784) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L0), .B(SubCellInst_SboxInst_8_T3), .Z(
        AddRoundConstantOutput[32]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1741), 
        .B(new_AGEMA_signal_1694), .Z(new_AGEMA_signal_1785) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_3114), .B(SubCellInst_SboxInst_8_YY_3), .ZN(AddRoundConstantOutput[33]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3116), .B(new_AGEMA_signal_1784), .Z(new_AGEMA_signal_1834) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U14 ( .A(Fresh[50]), .B(
        SubCellInst_SboxInst_9_Q2), .Z(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U13 ( .A(Fresh[50]), .B(
        new_AGEMA_signal_1632), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U10 ( .A1(new_AGEMA_signal_3120), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U9 ( .A1(new_AGEMA_signal_3118), .A2(
        SubCellInst_SboxInst_9_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U8 ( .A(Fresh[50]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U7 ( .A1(new_AGEMA_signal_1632), .A2(
        new_AGEMA_signal_3120), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_9_Q2), 
        .A2(new_AGEMA_signal_3118), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n8), .B(
        SubCellInst_SboxInst_9_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1697) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n7), .B(
        SubCellInst_SboxInst_9_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_9_T1) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3118), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3120), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_T1), .B(new_AGEMA_signal_3122), .Z(
        SubCellInst_SboxInst_9_L0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1697), 
        .B(new_AGEMA_signal_3124), .Z(new_AGEMA_signal_1743) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U14 ( .A(Fresh[51]), .B(
        SubCellInst_SboxInst_9_Q7), .Z(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U13 ( .A(Fresh[51]), .B(
        new_AGEMA_signal_1633), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U10 ( .A1(new_AGEMA_signal_3128), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U9 ( .A1(new_AGEMA_signal_3126), .A2(
        SubCellInst_SboxInst_9_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U8 ( .A(Fresh[51]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U7 ( .A1(new_AGEMA_signal_1633), .A2(
        new_AGEMA_signal_3128), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_9_Q7), 
        .A2(new_AGEMA_signal_3126), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n8), .B(
        SubCellInst_SboxInst_9_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1698) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n7), .B(
        SubCellInst_SboxInst_9_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_9_T3) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3126), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3128), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L0), .B(new_AGEMA_signal_3132), .Z(
        SubCellInst_SboxInst_9_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1743), 
        .B(new_AGEMA_signal_3136), .Z(new_AGEMA_signal_1786) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L0), .B(SubCellInst_SboxInst_9_T3), .Z(
        AddRoundConstantOutput[36]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1743), 
        .B(new_AGEMA_signal_1698), .Z(new_AGEMA_signal_1787) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_3138), .B(SubCellInst_SboxInst_9_YY_3), .ZN(AddRoundConstantOutput[37]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3140), .B(new_AGEMA_signal_1786), .Z(new_AGEMA_signal_1835) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U14 ( .A(Fresh[52]), .B(
        SubCellInst_SboxInst_10_Q2), .Z(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U13 ( .A(Fresh[52]), .B(
        new_AGEMA_signal_1636), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U10 ( .A1(new_AGEMA_signal_3144), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U9 ( .A1(new_AGEMA_signal_3142), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U8 ( .A(Fresh[52]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U7 ( .A1(new_AGEMA_signal_1636), 
        .A2(new_AGEMA_signal_3144), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_10_Q2), 
        .A2(new_AGEMA_signal_3142), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n8), .B(
        SubCellInst_SboxInst_10_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1701)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n7), .B(
        SubCellInst_SboxInst_10_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_10_T1) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3142), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3144), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_T1), .B(new_AGEMA_signal_3146), .Z(
        SubCellInst_SboxInst_10_L0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1701), 
        .B(new_AGEMA_signal_3148), .Z(new_AGEMA_signal_1745) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U14 ( .A(Fresh[53]), .B(
        SubCellInst_SboxInst_10_Q7), .Z(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U13 ( .A(Fresh[53]), .B(
        new_AGEMA_signal_1637), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U10 ( .A1(new_AGEMA_signal_3152), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U9 ( .A1(new_AGEMA_signal_3150), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U8 ( .A(Fresh[53]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U7 ( .A1(new_AGEMA_signal_1637), 
        .A2(new_AGEMA_signal_3152), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_10_Q7), 
        .A2(new_AGEMA_signal_3150), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n8), .B(
        SubCellInst_SboxInst_10_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1702)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n7), .B(
        SubCellInst_SboxInst_10_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_10_T3) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3150), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3152), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L0), .B(new_AGEMA_signal_3156), .Z(
        SubCellInst_SboxInst_10_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1745), 
        .B(new_AGEMA_signal_3160), .Z(new_AGEMA_signal_1788) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L0), .B(SubCellInst_SboxInst_10_T3), .Z(
        AddRoundConstantOutput[40]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1745), .B(new_AGEMA_signal_1702), .Z(new_AGEMA_signal_1789) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_3162), .B(SubCellInst_SboxInst_10_YY_3), .ZN(
        AddRoundConstantOutput[41]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3164), .B(new_AGEMA_signal_1788), .Z(
        new_AGEMA_signal_1836) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U14 ( .A(Fresh[54]), .B(
        SubCellInst_SboxInst_11_Q2), .Z(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U13 ( .A(Fresh[54]), .B(
        new_AGEMA_signal_1640), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U10 ( .A1(new_AGEMA_signal_3168), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U9 ( .A1(new_AGEMA_signal_3166), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U8 ( .A(Fresh[54]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U7 ( .A1(new_AGEMA_signal_1640), 
        .A2(new_AGEMA_signal_3168), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_11_Q2), 
        .A2(new_AGEMA_signal_3166), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n8), .B(
        SubCellInst_SboxInst_11_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1705)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n7), .B(
        SubCellInst_SboxInst_11_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_11_T1) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3166), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3168), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_T1), .B(new_AGEMA_signal_3170), .Z(
        SubCellInst_SboxInst_11_L0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1705), 
        .B(new_AGEMA_signal_3172), .Z(new_AGEMA_signal_1747) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U14 ( .A(Fresh[55]), .B(
        SubCellInst_SboxInst_11_Q7), .Z(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U13 ( .A(Fresh[55]), .B(
        new_AGEMA_signal_1641), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U10 ( .A1(new_AGEMA_signal_3176), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U9 ( .A1(new_AGEMA_signal_3174), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U8 ( .A(Fresh[55]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U7 ( .A1(new_AGEMA_signal_1641), 
        .A2(new_AGEMA_signal_3176), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_11_Q7), 
        .A2(new_AGEMA_signal_3174), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n8), .B(
        SubCellInst_SboxInst_11_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1706)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n7), .B(
        SubCellInst_SboxInst_11_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_11_T3) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3174), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3176), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L0), .B(new_AGEMA_signal_3180), .Z(
        SubCellInst_SboxInst_11_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1747), 
        .B(new_AGEMA_signal_3184), .Z(new_AGEMA_signal_1790) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L0), .B(SubCellInst_SboxInst_11_T3), .Z(
        SubCellOutput_44) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1747), .B(new_AGEMA_signal_1706), .Z(new_AGEMA_signal_1791) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_3186), .B(SubCellInst_SboxInst_11_YY_3), .ZN(
        SubCellOutput_45) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3188), .B(new_AGEMA_signal_1790), .Z(
        new_AGEMA_signal_1837) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U14 ( .A(Fresh[56]), .B(
        SubCellInst_SboxInst_12_Q2), .Z(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U13 ( .A(Fresh[56]), .B(
        new_AGEMA_signal_1644), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U10 ( .A1(new_AGEMA_signal_3192), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U9 ( .A1(new_AGEMA_signal_3190), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U8 ( .A(Fresh[56]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U7 ( .A1(new_AGEMA_signal_1644), 
        .A2(new_AGEMA_signal_3192), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_12_Q2), 
        .A2(new_AGEMA_signal_3190), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n8), .B(
        SubCellInst_SboxInst_12_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1709)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n7), .B(
        SubCellInst_SboxInst_12_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_12_T1) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3190), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3192), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_T1), .B(new_AGEMA_signal_3194), .Z(
        SubCellInst_SboxInst_12_L0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1709), 
        .B(new_AGEMA_signal_3196), .Z(new_AGEMA_signal_1749) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U14 ( .A(Fresh[57]), .B(
        SubCellInst_SboxInst_12_Q7), .Z(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U13 ( .A(Fresh[57]), .B(
        new_AGEMA_signal_1645), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U10 ( .A1(new_AGEMA_signal_3200), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U9 ( .A1(new_AGEMA_signal_3198), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U8 ( .A(Fresh[57]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U7 ( .A1(new_AGEMA_signal_1645), 
        .A2(new_AGEMA_signal_3200), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_12_Q7), 
        .A2(new_AGEMA_signal_3198), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n8), .B(
        SubCellInst_SboxInst_12_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1710)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n7), .B(
        SubCellInst_SboxInst_12_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_12_T3) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3198), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3200), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L0), .B(new_AGEMA_signal_3204), .Z(
        SubCellInst_SboxInst_12_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1749), 
        .B(new_AGEMA_signal_3208), .Z(new_AGEMA_signal_1792) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L0), .B(SubCellInst_SboxInst_12_T3), .Z(
        AddRoundConstantOutput[48]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1749), .B(new_AGEMA_signal_1710), .Z(new_AGEMA_signal_1793) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_3210), .B(SubCellInst_SboxInst_12_YY_3), .ZN(
        AddRoundConstantOutput[49]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3212), .B(new_AGEMA_signal_1792), .Z(
        new_AGEMA_signal_1838) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U14 ( .A(Fresh[58]), .B(
        SubCellInst_SboxInst_13_Q2), .Z(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U13 ( .A(Fresh[58]), .B(
        new_AGEMA_signal_1648), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U10 ( .A1(new_AGEMA_signal_3216), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U9 ( .A1(new_AGEMA_signal_3214), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U8 ( .A(Fresh[58]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U7 ( .A1(new_AGEMA_signal_1648), 
        .A2(new_AGEMA_signal_3216), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_13_Q2), 
        .A2(new_AGEMA_signal_3214), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n8), .B(
        SubCellInst_SboxInst_13_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1713)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n7), .B(
        SubCellInst_SboxInst_13_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_13_T1) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3214), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3216), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_T1), .B(new_AGEMA_signal_3218), .Z(
        SubCellInst_SboxInst_13_L0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1713), 
        .B(new_AGEMA_signal_3220), .Z(new_AGEMA_signal_1751) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U14 ( .A(Fresh[59]), .B(
        SubCellInst_SboxInst_13_Q7), .Z(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U13 ( .A(Fresh[59]), .B(
        new_AGEMA_signal_1649), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U10 ( .A1(new_AGEMA_signal_3224), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U9 ( .A1(new_AGEMA_signal_3222), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U8 ( .A(Fresh[59]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U7 ( .A1(new_AGEMA_signal_1649), 
        .A2(new_AGEMA_signal_3224), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_13_Q7), 
        .A2(new_AGEMA_signal_3222), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n8), .B(
        SubCellInst_SboxInst_13_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1714)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n7), .B(
        SubCellInst_SboxInst_13_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_13_T3) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3222), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3224), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L0), .B(new_AGEMA_signal_3228), .Z(
        SubCellInst_SboxInst_13_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1751), 
        .B(new_AGEMA_signal_3232), .Z(new_AGEMA_signal_1794) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L0), .B(SubCellInst_SboxInst_13_T3), .Z(
        AddRoundConstantOutput[52]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1751), .B(new_AGEMA_signal_1714), .Z(new_AGEMA_signal_1795) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_3234), .B(SubCellInst_SboxInst_13_YY_3), .ZN(
        AddRoundConstantOutput[53]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3236), .B(new_AGEMA_signal_1794), .Z(
        new_AGEMA_signal_1839) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U14 ( .A(Fresh[60]), .B(
        SubCellInst_SboxInst_14_Q2), .Z(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U13 ( .A(Fresh[60]), .B(
        new_AGEMA_signal_1652), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U10 ( .A1(new_AGEMA_signal_3240), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U9 ( .A1(new_AGEMA_signal_3238), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U8 ( .A(Fresh[60]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U7 ( .A1(new_AGEMA_signal_1652), 
        .A2(new_AGEMA_signal_3240), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_14_Q2), 
        .A2(new_AGEMA_signal_3238), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n8), .B(
        SubCellInst_SboxInst_14_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1717)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n7), .B(
        SubCellInst_SboxInst_14_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_14_T1) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3238), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3240), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_T1), .B(new_AGEMA_signal_3242), .Z(
        SubCellInst_SboxInst_14_L0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1717), 
        .B(new_AGEMA_signal_3244), .Z(new_AGEMA_signal_1753) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U14 ( .A(Fresh[61]), .B(
        SubCellInst_SboxInst_14_Q7), .Z(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U13 ( .A(Fresh[61]), .B(
        new_AGEMA_signal_1653), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U10 ( .A1(new_AGEMA_signal_3248), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U9 ( .A1(new_AGEMA_signal_3246), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U8 ( .A(Fresh[61]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U7 ( .A1(new_AGEMA_signal_1653), 
        .A2(new_AGEMA_signal_3248), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_14_Q7), 
        .A2(new_AGEMA_signal_3246), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n8), .B(
        SubCellInst_SboxInst_14_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1718)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n7), .B(
        SubCellInst_SboxInst_14_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_14_T3) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3246), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3248), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L0), .B(new_AGEMA_signal_3252), .Z(
        SubCellInst_SboxInst_14_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1753), 
        .B(new_AGEMA_signal_3256), .Z(new_AGEMA_signal_1796) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L0), .B(SubCellInst_SboxInst_14_T3), .Z(
        AddRoundConstantOutput[56]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1753), .B(new_AGEMA_signal_1718), .Z(new_AGEMA_signal_1797) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_3258), .B(SubCellInst_SboxInst_14_YY_3), .ZN(
        AddRoundConstantOutput[57]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3260), .B(new_AGEMA_signal_1796), .Z(
        new_AGEMA_signal_1840) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U14 ( .A(Fresh[62]), .B(
        SubCellInst_SboxInst_15_Q2), .Z(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U13 ( .A(Fresh[62]), .B(
        new_AGEMA_signal_1656), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U10 ( .A1(new_AGEMA_signal_3264), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U9 ( .A1(new_AGEMA_signal_3262), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U8 ( .A(Fresh[62]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U7 ( .A1(new_AGEMA_signal_1656), 
        .A2(new_AGEMA_signal_3264), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_15_Q2), 
        .A2(new_AGEMA_signal_3262), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n8), .B(
        SubCellInst_SboxInst_15_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1721)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n7), .B(
        SubCellInst_SboxInst_15_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_15_T1) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3262), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3264), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_T1), .B(new_AGEMA_signal_3266), .Z(
        SubCellInst_SboxInst_15_L0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1721), 
        .B(new_AGEMA_signal_3268), .Z(new_AGEMA_signal_1755) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U14 ( .A(Fresh[63]), .B(
        SubCellInst_SboxInst_15_Q7), .Z(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U13 ( .A(Fresh[63]), .B(
        new_AGEMA_signal_1657), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U10 ( .A1(new_AGEMA_signal_3272), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U9 ( .A1(new_AGEMA_signal_3270), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U8 ( .A(Fresh[63]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U7 ( .A1(new_AGEMA_signal_1657), 
        .A2(new_AGEMA_signal_3272), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_15_Q7), 
        .A2(new_AGEMA_signal_3270), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n8), .B(
        SubCellInst_SboxInst_15_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1722)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n7), .B(
        SubCellInst_SboxInst_15_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_15_T3) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3270), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3272), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L0), .B(new_AGEMA_signal_3276), .Z(
        SubCellInst_SboxInst_15_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1755), 
        .B(new_AGEMA_signal_3280), .Z(new_AGEMA_signal_1798) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L0), .B(SubCellInst_SboxInst_15_T3), .Z(
        SubCellOutput[60]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1755), .B(new_AGEMA_signal_1722), .Z(new_AGEMA_signal_1799) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_3282), .B(SubCellInst_SboxInst_15_YY_3), .ZN(
        SubCellOutput[61]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3284), .B(new_AGEMA_signal_1798), .Z(
        new_AGEMA_signal_1841) );
  INV_X1 AddConstXOR_U2_U1 ( .A(SubCellOutput_29), .ZN(ShiftRowsOutput[21]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_0_n1), .B(new_AGEMA_signal_3288), 
        .ZN(AddRoundConstantOutput[60]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1842), .B(1'b0), .Z(new_AGEMA_signal_1880) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[60]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_0_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1799), .Z(new_AGEMA_signal_1842) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_1_n1), .B(new_AGEMA_signal_3292), 
        .ZN(AddRoundConstantOutput[61]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1881), .B(1'b0), .Z(new_AGEMA_signal_1947) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[61]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_1_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1841), .Z(new_AGEMA_signal_1881) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_0_n1), .B(new_AGEMA_signal_3296), 
        .ZN(AddRoundConstantOutput[44]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1844), .B(1'b0), .Z(new_AGEMA_signal_1882) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_44), .ZN(AddConstXOR_AddConstXOR_XORInst_1_0_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1791), .Z(new_AGEMA_signal_1844) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_1_n1), .B(new_AGEMA_signal_3300), 
        .ZN(AddRoundConstantOutput[45]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1883), .B(1'b0), .Z(new_AGEMA_signal_1948) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_45), .ZN(AddConstXOR_AddConstXOR_XORInst_1_1_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1837), .Z(new_AGEMA_signal_1883) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_0_n1), .B(new_AGEMA_signal_3304), .ZN(
        ShiftRowsOutput[44]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1846), .B(new_AGEMA_signal_3308), .Z(
        new_AGEMA_signal_1884) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[32]), .ZN(AddRoundTweakeyXOR_XORInst_0_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1785), .Z(new_AGEMA_signal_1846) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_1_n1), .B(new_AGEMA_signal_3312), .ZN(
        ShiftRowsOutput[45]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1885), .B(new_AGEMA_signal_3316), .Z(
        new_AGEMA_signal_1949) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[33]), .ZN(AddRoundTweakeyXOR_XORInst_0_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1834), .Z(new_AGEMA_signal_1885) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_0_n1), .B(new_AGEMA_signal_3320), .ZN(
        ShiftRowsOutput[32]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1848), .B(new_AGEMA_signal_3324), .Z(
        new_AGEMA_signal_1886) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[36]), .ZN(AddRoundTweakeyXOR_XORInst_1_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1787), .Z(new_AGEMA_signal_1848) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_1_n1), .B(new_AGEMA_signal_3328), .ZN(
        ShiftRowsOutput[33]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1887), .B(new_AGEMA_signal_3332), .Z(
        new_AGEMA_signal_1950) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[37]), .ZN(AddRoundTweakeyXOR_XORInst_1_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1835), .Z(new_AGEMA_signal_1887) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_0_n1), .B(new_AGEMA_signal_3336), .ZN(
        ShiftRowsOutput[36]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1850), .B(new_AGEMA_signal_3340), .Z(
        new_AGEMA_signal_1888) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[40]), .ZN(AddRoundTweakeyXOR_XORInst_2_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1789), .Z(new_AGEMA_signal_1850) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_1_n1), .B(new_AGEMA_signal_3344), .ZN(
        ShiftRowsOutput[37]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1889), .B(new_AGEMA_signal_3348), .Z(
        new_AGEMA_signal_1951) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[41]), .ZN(AddRoundTweakeyXOR_XORInst_2_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1836), .Z(new_AGEMA_signal_1889) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_0_n1), .B(new_AGEMA_signal_3352), .ZN(
        ShiftRowsOutput[40]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1952), .B(new_AGEMA_signal_3356), .Z(
        new_AGEMA_signal_2007) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[44]), .ZN(AddRoundTweakeyXOR_XORInst_3_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1882), .Z(new_AGEMA_signal_1952) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_1_n1), .B(new_AGEMA_signal_3360), .ZN(
        ShiftRowsOutput[41]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2008), .B(new_AGEMA_signal_3364), .Z(
        new_AGEMA_signal_2061) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[45]), .ZN(AddRoundTweakeyXOR_XORInst_3_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1948), .Z(new_AGEMA_signal_2008) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_0_n1), .B(new_AGEMA_signal_3368), .ZN(
        MCOutput[32]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1853), .B(new_AGEMA_signal_3372), .Z(
        new_AGEMA_signal_1892) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[48]), .ZN(AddRoundTweakeyXOR_XORInst_4_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1793), .Z(new_AGEMA_signal_1853) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_1_n1), .B(new_AGEMA_signal_3376), .ZN(
        MCOutput[33]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1893), .B(new_AGEMA_signal_3380), .Z(
        new_AGEMA_signal_1954) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[49]), .ZN(AddRoundTweakeyXOR_XORInst_4_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1838), .Z(new_AGEMA_signal_1893) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_0_n1), .B(new_AGEMA_signal_3384), .ZN(
        MCOutput[36]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1855), .B(new_AGEMA_signal_3388), .Z(
        new_AGEMA_signal_1894) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[52]), .ZN(AddRoundTweakeyXOR_XORInst_5_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1795), .Z(new_AGEMA_signal_1855) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_1_n1), .B(new_AGEMA_signal_3392), .ZN(
        MCOutput[37]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1895), .B(new_AGEMA_signal_3396), .Z(
        new_AGEMA_signal_1955) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[53]), .ZN(AddRoundTweakeyXOR_XORInst_5_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1839), .Z(new_AGEMA_signal_1895) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_0_n1), .B(new_AGEMA_signal_3400), .ZN(
        MCOutput[40]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1857), .B(new_AGEMA_signal_3404), .Z(
        new_AGEMA_signal_1896) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[56]), .ZN(AddRoundTweakeyXOR_XORInst_6_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1797), .Z(new_AGEMA_signal_1857) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_1_n1), .B(new_AGEMA_signal_3408), .ZN(
        MCOutput[41]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1897), .B(new_AGEMA_signal_3412), .Z(
        new_AGEMA_signal_1956) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[57]), .ZN(AddRoundTweakeyXOR_XORInst_6_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1840), .Z(new_AGEMA_signal_1897) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_0_n1), .B(new_AGEMA_signal_3416), .ZN(
        MCOutput[44]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1957), .B(new_AGEMA_signal_3420), .Z(
        new_AGEMA_signal_2009) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[60]), .ZN(AddRoundTweakeyXOR_XORInst_7_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1880), .Z(new_AGEMA_signal_1957) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_1_n1), .B(new_AGEMA_signal_3424), .ZN(
        MCOutput[45]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2010), .B(new_AGEMA_signal_3428), .Z(
        new_AGEMA_signal_2062) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[61]), .ZN(AddRoundTweakeyXOR_XORInst_7_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1947), .Z(new_AGEMA_signal_2010) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_0_n2), 
        .B(MCInst_MCR0_XORInst_0_0_n1), .ZN(MCOutput[48]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1959), .B(
        new_AGEMA_signal_1860), .Z(new_AGEMA_signal_2011) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[16]), .B(
        ShiftRowsOutput[0]), .ZN(MCInst_MCR0_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1781), .B(
        new_AGEMA_signal_1775), .Z(new_AGEMA_signal_1860) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[32]), 
        .Z(MCInst_MCR0_XORInst_0_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1892), .Z(new_AGEMA_signal_1959) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_1_n2), 
        .B(MCInst_MCR0_XORInst_0_1_n1), .ZN(MCOutput[49]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2012), .B(
        new_AGEMA_signal_1900), .Z(new_AGEMA_signal_2063) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[17]), .B(
        ShiftRowsOutput[1]), .ZN(MCInst_MCR0_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1832), .B(
        new_AGEMA_signal_1829), .Z(new_AGEMA_signal_1900) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[33]), 
        .Z(MCInst_MCR0_XORInst_0_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1954), .Z(new_AGEMA_signal_2012) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_0_n2), 
        .B(MCInst_MCR0_XORInst_1_0_n1), .ZN(MCOutput[52]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1961), .B(
        new_AGEMA_signal_1862), .Z(new_AGEMA_signal_2013) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[20]), .B(
        ShiftRowsOutput[4]), .ZN(MCInst_MCR0_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1783), .B(
        new_AGEMA_signal_1769), .Z(new_AGEMA_signal_1862) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[36]), 
        .Z(MCInst_MCR0_XORInst_1_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1894), .Z(new_AGEMA_signal_1961) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_1_n2), 
        .B(MCInst_MCR0_XORInst_1_1_n1), .ZN(MCOutput[53]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2014), .B(
        new_AGEMA_signal_1962), .Z(new_AGEMA_signal_2064) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[21]), .B(
        ShiftRowsOutput[5]), .ZN(MCInst_MCR0_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1879), .B(
        new_AGEMA_signal_1826), .Z(new_AGEMA_signal_1962) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[37]), 
        .Z(MCInst_MCR0_XORInst_1_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1955), .Z(new_AGEMA_signal_2014) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_0_n2), 
        .B(MCInst_MCR0_XORInst_2_0_n1), .ZN(MCOutput[56]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1964), .B(
        new_AGEMA_signal_1864), .Z(new_AGEMA_signal_2015) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[24]), .B(
        ShiftRowsOutput[8]), .ZN(MCInst_MCR0_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1777), .B(
        new_AGEMA_signal_1771), .Z(new_AGEMA_signal_1864) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[40]), 
        .Z(MCInst_MCR0_XORInst_2_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1896), .Z(new_AGEMA_signal_1964) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_1_n2), 
        .B(MCInst_MCR0_XORInst_2_1_n1), .ZN(MCOutput[57]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2016), .B(
        new_AGEMA_signal_1905), .Z(new_AGEMA_signal_2065) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[25]), .B(
        ShiftRowsOutput[9]), .ZN(MCInst_MCR0_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1830), .B(
        new_AGEMA_signal_1827), .Z(new_AGEMA_signal_1905) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[41]), 
        .Z(MCInst_MCR0_XORInst_2_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1956), .Z(new_AGEMA_signal_2016) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_0_n2), 
        .B(MCInst_MCR0_XORInst_3_0_n1), .ZN(MCOutput[60]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2066), .B(
        new_AGEMA_signal_1866), .Z(new_AGEMA_signal_2104) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[28]), .B(
        ShiftRowsOutput[12]), .ZN(MCInst_MCR0_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1779), .B(
        new_AGEMA_signal_1773), .Z(new_AGEMA_signal_1866) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[44]), 
        .Z(MCInst_MCR0_XORInst_3_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2009), .Z(new_AGEMA_signal_2066) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_1_n2), 
        .B(MCInst_MCR0_XORInst_3_1_n1), .ZN(MCOutput[61]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2105), .B(
        new_AGEMA_signal_1908), .Z(new_AGEMA_signal_2116) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[29]), .B(
        ShiftRowsOutput[13]), .ZN(MCInst_MCR0_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1831), .B(
        new_AGEMA_signal_1828), .Z(new_AGEMA_signal_1908) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[45]), 
        .Z(MCInst_MCR0_XORInst_3_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2062), .Z(new_AGEMA_signal_2105) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_0_n1), 
        .B(ShiftRowsOutput[16]), .ZN(MCOutput[16]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1967), .B(
        new_AGEMA_signal_1781), .Z(new_AGEMA_signal_2019) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[32]), .ZN(MCInst_MCR2_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1886), .Z(new_AGEMA_signal_1967) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_1_n1), 
        .B(ShiftRowsOutput[17]), .ZN(MCOutput[17]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2020), .B(
        new_AGEMA_signal_1832), .Z(new_AGEMA_signal_2068) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[33]), .ZN(MCInst_MCR2_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1950), .Z(new_AGEMA_signal_2020) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_0_n1), 
        .B(ShiftRowsOutput[20]), .ZN(MCOutput[20]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1969), .B(
        new_AGEMA_signal_1783), .Z(new_AGEMA_signal_2021) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[36]), .ZN(MCInst_MCR2_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1888), .Z(new_AGEMA_signal_1969) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_1_n1), 
        .B(ShiftRowsOutput[21]), .ZN(MCOutput[21]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2022), .B(
        new_AGEMA_signal_1879), .Z(new_AGEMA_signal_2069) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[37]), .ZN(MCInst_MCR2_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1951), .Z(new_AGEMA_signal_2022) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_0_n1), 
        .B(ShiftRowsOutput[24]), .ZN(MCOutput[24]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2070), .B(
        new_AGEMA_signal_1777), .Z(new_AGEMA_signal_2106) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[40]), .ZN(MCInst_MCR2_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2007), .Z(new_AGEMA_signal_2070) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_1_n1), 
        .B(ShiftRowsOutput[25]), .ZN(MCOutput[25]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2107), .B(
        new_AGEMA_signal_1830), .Z(new_AGEMA_signal_2117) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[41]), .ZN(MCInst_MCR2_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2061), .Z(new_AGEMA_signal_2107) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_0_n1), 
        .B(ShiftRowsOutput[28]), .ZN(MCOutput[28]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1972), .B(
        new_AGEMA_signal_1779), .Z(new_AGEMA_signal_2025) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[44]), .ZN(MCInst_MCR2_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1884), .Z(new_AGEMA_signal_1972) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_1_n1), 
        .B(ShiftRowsOutput[29]), .ZN(MCOutput[29]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2026), .B(
        new_AGEMA_signal_1831), .Z(new_AGEMA_signal_2072) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[45]), .ZN(MCInst_MCR2_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1949), .Z(new_AGEMA_signal_2026) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_0_n1), 
        .B(ShiftRowsOutput[16]), .ZN(MCOutput[0]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1974), .B(
        new_AGEMA_signal_1781), .Z(new_AGEMA_signal_2027) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[32]), 
        .ZN(MCInst_MCR3_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1892), .Z(new_AGEMA_signal_1974) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_1_n1), 
        .B(ShiftRowsOutput[17]), .ZN(MCOutput[1]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2028), .B(
        new_AGEMA_signal_1832), .Z(new_AGEMA_signal_2073) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[33]), 
        .ZN(MCInst_MCR3_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1954), .Z(new_AGEMA_signal_2028) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_0_n1), 
        .B(ShiftRowsOutput[20]), .ZN(MCOutput[4]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1976), .B(
        new_AGEMA_signal_1783), .Z(new_AGEMA_signal_2029) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[36]), 
        .ZN(MCInst_MCR3_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1894), .Z(new_AGEMA_signal_1976) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_1_n1), 
        .B(ShiftRowsOutput[21]), .ZN(MCOutput[5]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2030), .B(
        new_AGEMA_signal_1879), .Z(new_AGEMA_signal_2074) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[37]), 
        .ZN(MCInst_MCR3_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1955), .Z(new_AGEMA_signal_2030) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_0_n1), 
        .B(ShiftRowsOutput[24]), .ZN(MCOutput[8]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1978), .B(
        new_AGEMA_signal_1777), .Z(new_AGEMA_signal_2031) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[40]), 
        .ZN(MCInst_MCR3_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1896), .Z(new_AGEMA_signal_1978) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_1_n1), 
        .B(ShiftRowsOutput[25]), .ZN(MCOutput[9]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2032), .B(
        new_AGEMA_signal_1830), .Z(new_AGEMA_signal_2075) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[41]), 
        .ZN(MCInst_MCR3_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1956), .Z(new_AGEMA_signal_2032) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_0_n1), 
        .B(ShiftRowsOutput[28]), .ZN(MCOutput[12]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2076), .B(
        new_AGEMA_signal_1779), .Z(new_AGEMA_signal_2108) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[44]), 
        .ZN(MCInst_MCR3_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2009), .Z(new_AGEMA_signal_2076) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_1_n1), 
        .B(ShiftRowsOutput[29]), .ZN(MCOutput[13]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2109), .B(
        new_AGEMA_signal_1831), .Z(new_AGEMA_signal_2118) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[45]), 
        .ZN(MCInst_MCR3_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2062), .Z(new_AGEMA_signal_2109) );
  DFF_X1 new_AGEMA_reg_buffer_1455_s_current_state_reg ( .D(
        new_AGEMA_signal_2643), .CK(clk), .Q(new_AGEMA_signal_2644), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1459_s_current_state_reg ( .D(
        new_AGEMA_signal_2647), .CK(clk), .Q(new_AGEMA_signal_2648), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1463_s_current_state_reg ( .D(
        new_AGEMA_signal_2651), .CK(clk), .Q(new_AGEMA_signal_2652), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1467_s_current_state_reg ( .D(
        new_AGEMA_signal_2655), .CK(clk), .Q(new_AGEMA_signal_2656), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1471_s_current_state_reg ( .D(
        new_AGEMA_signal_2659), .CK(clk), .Q(new_AGEMA_signal_2660), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1475_s_current_state_reg ( .D(
        new_AGEMA_signal_2663), .CK(clk), .Q(new_AGEMA_signal_2664), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1479_s_current_state_reg ( .D(
        new_AGEMA_signal_2667), .CK(clk), .Q(new_AGEMA_signal_2668), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1483_s_current_state_reg ( .D(
        new_AGEMA_signal_2671), .CK(clk), .Q(new_AGEMA_signal_2672), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1487_s_current_state_reg ( .D(
        new_AGEMA_signal_2675), .CK(clk), .Q(new_AGEMA_signal_2676), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1491_s_current_state_reg ( .D(
        new_AGEMA_signal_2679), .CK(clk), .Q(new_AGEMA_signal_2680), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1495_s_current_state_reg ( .D(
        new_AGEMA_signal_2683), .CK(clk), .Q(new_AGEMA_signal_2684), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1499_s_current_state_reg ( .D(
        new_AGEMA_signal_2687), .CK(clk), .Q(new_AGEMA_signal_2688), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1503_s_current_state_reg ( .D(
        new_AGEMA_signal_2691), .CK(clk), .Q(new_AGEMA_signal_2692), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1507_s_current_state_reg ( .D(
        new_AGEMA_signal_2695), .CK(clk), .Q(new_AGEMA_signal_2696), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1511_s_current_state_reg ( .D(
        new_AGEMA_signal_2699), .CK(clk), .Q(new_AGEMA_signal_2700), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1515_s_current_state_reg ( .D(
        new_AGEMA_signal_2703), .CK(clk), .Q(new_AGEMA_signal_2704), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1519_s_current_state_reg ( .D(
        new_AGEMA_signal_2707), .CK(clk), .Q(new_AGEMA_signal_2708), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1523_s_current_state_reg ( .D(
        new_AGEMA_signal_2711), .CK(clk), .Q(new_AGEMA_signal_2712), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1527_s_current_state_reg ( .D(
        new_AGEMA_signal_2715), .CK(clk), .Q(new_AGEMA_signal_2716), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1531_s_current_state_reg ( .D(
        new_AGEMA_signal_2719), .CK(clk), .Q(new_AGEMA_signal_2720), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1535_s_current_state_reg ( .D(
        new_AGEMA_signal_2723), .CK(clk), .Q(new_AGEMA_signal_2724), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1539_s_current_state_reg ( .D(
        new_AGEMA_signal_2727), .CK(clk), .Q(new_AGEMA_signal_2728), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1543_s_current_state_reg ( .D(
        new_AGEMA_signal_2731), .CK(clk), .Q(new_AGEMA_signal_2732), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1547_s_current_state_reg ( .D(
        new_AGEMA_signal_2735), .CK(clk), .Q(new_AGEMA_signal_2736), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1551_s_current_state_reg ( .D(
        new_AGEMA_signal_2739), .CK(clk), .Q(new_AGEMA_signal_2740), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1555_s_current_state_reg ( .D(
        new_AGEMA_signal_2743), .CK(clk), .Q(new_AGEMA_signal_2744), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1559_s_current_state_reg ( .D(
        new_AGEMA_signal_2747), .CK(clk), .Q(new_AGEMA_signal_2748), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1563_s_current_state_reg ( .D(
        new_AGEMA_signal_2751), .CK(clk), .Q(new_AGEMA_signal_2752), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1567_s_current_state_reg ( .D(
        new_AGEMA_signal_2755), .CK(clk), .Q(new_AGEMA_signal_2756), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1571_s_current_state_reg ( .D(
        new_AGEMA_signal_2759), .CK(clk), .Q(new_AGEMA_signal_2760), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1575_s_current_state_reg ( .D(
        new_AGEMA_signal_2763), .CK(clk), .Q(new_AGEMA_signal_2764), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1579_s_current_state_reg ( .D(
        new_AGEMA_signal_2767), .CK(clk), .Q(new_AGEMA_signal_2768), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1583_s_current_state_reg ( .D(
        new_AGEMA_signal_2771), .CK(clk), .Q(new_AGEMA_signal_2772), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1587_s_current_state_reg ( .D(
        new_AGEMA_signal_2775), .CK(clk), .Q(new_AGEMA_signal_2776), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1591_s_current_state_reg ( .D(
        new_AGEMA_signal_2779), .CK(clk), .Q(new_AGEMA_signal_2780), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1595_s_current_state_reg ( .D(
        new_AGEMA_signal_2783), .CK(clk), .Q(new_AGEMA_signal_2784), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1599_s_current_state_reg ( .D(
        new_AGEMA_signal_2787), .CK(clk), .Q(new_AGEMA_signal_2788), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1603_s_current_state_reg ( .D(
        new_AGEMA_signal_2791), .CK(clk), .Q(new_AGEMA_signal_2792), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1607_s_current_state_reg ( .D(
        new_AGEMA_signal_2795), .CK(clk), .Q(new_AGEMA_signal_2796), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1611_s_current_state_reg ( .D(
        new_AGEMA_signal_2799), .CK(clk), .Q(new_AGEMA_signal_2800), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1615_s_current_state_reg ( .D(
        new_AGEMA_signal_2803), .CK(clk), .Q(new_AGEMA_signal_2804), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1619_s_current_state_reg ( .D(
        new_AGEMA_signal_2807), .CK(clk), .Q(new_AGEMA_signal_2808), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1623_s_current_state_reg ( .D(
        new_AGEMA_signal_2811), .CK(clk), .Q(new_AGEMA_signal_2812), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1627_s_current_state_reg ( .D(
        new_AGEMA_signal_2815), .CK(clk), .Q(new_AGEMA_signal_2816), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1631_s_current_state_reg ( .D(
        new_AGEMA_signal_2819), .CK(clk), .Q(new_AGEMA_signal_2820), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1635_s_current_state_reg ( .D(
        new_AGEMA_signal_2823), .CK(clk), .Q(new_AGEMA_signal_2824), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1639_s_current_state_reg ( .D(
        new_AGEMA_signal_2827), .CK(clk), .Q(new_AGEMA_signal_2828), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1643_s_current_state_reg ( .D(
        new_AGEMA_signal_2831), .CK(clk), .Q(new_AGEMA_signal_2832), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1647_s_current_state_reg ( .D(
        new_AGEMA_signal_2835), .CK(clk), .Q(new_AGEMA_signal_2836), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1651_s_current_state_reg ( .D(
        new_AGEMA_signal_2839), .CK(clk), .Q(new_AGEMA_signal_2840), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1655_s_current_state_reg ( .D(
        new_AGEMA_signal_2843), .CK(clk), .Q(new_AGEMA_signal_2844), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1659_s_current_state_reg ( .D(
        new_AGEMA_signal_2847), .CK(clk), .Q(new_AGEMA_signal_2848), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1663_s_current_state_reg ( .D(
        new_AGEMA_signal_2851), .CK(clk), .Q(new_AGEMA_signal_2852), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1667_s_current_state_reg ( .D(
        new_AGEMA_signal_2855), .CK(clk), .Q(new_AGEMA_signal_2856), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1671_s_current_state_reg ( .D(
        new_AGEMA_signal_2859), .CK(clk), .Q(new_AGEMA_signal_2860), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1675_s_current_state_reg ( .D(
        new_AGEMA_signal_2863), .CK(clk), .Q(new_AGEMA_signal_2864), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1679_s_current_state_reg ( .D(
        new_AGEMA_signal_2867), .CK(clk), .Q(new_AGEMA_signal_2868), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1683_s_current_state_reg ( .D(
        new_AGEMA_signal_2871), .CK(clk), .Q(new_AGEMA_signal_2872), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1687_s_current_state_reg ( .D(
        new_AGEMA_signal_2875), .CK(clk), .Q(new_AGEMA_signal_2876), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1691_s_current_state_reg ( .D(
        new_AGEMA_signal_2879), .CK(clk), .Q(new_AGEMA_signal_2880), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1695_s_current_state_reg ( .D(
        new_AGEMA_signal_2883), .CK(clk), .Q(new_AGEMA_signal_2884), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1699_s_current_state_reg ( .D(
        new_AGEMA_signal_2887), .CK(clk), .Q(new_AGEMA_signal_2888), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1703_s_current_state_reg ( .D(
        new_AGEMA_signal_2891), .CK(clk), .Q(new_AGEMA_signal_2892), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1707_s_current_state_reg ( .D(
        new_AGEMA_signal_2895), .CK(clk), .Q(new_AGEMA_signal_2896), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1711_s_current_state_reg ( .D(
        new_AGEMA_signal_2899), .CK(clk), .Q(new_AGEMA_signal_2900), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1717_s_current_state_reg ( .D(
        new_AGEMA_signal_2905), .CK(clk), .Q(new_AGEMA_signal_2906), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1719_s_current_state_reg ( .D(
        new_AGEMA_signal_2907), .CK(clk), .Q(new_AGEMA_signal_2908), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1727_s_current_state_reg ( .D(
        new_AGEMA_signal_2915), .CK(clk), .Q(new_AGEMA_signal_2916), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1731_s_current_state_reg ( .D(
        new_AGEMA_signal_2919), .CK(clk), .Q(new_AGEMA_signal_2920), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1733_s_current_state_reg ( .D(
        new_AGEMA_signal_2921), .CK(clk), .Q(new_AGEMA_signal_2922), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1735_s_current_state_reg ( .D(
        new_AGEMA_signal_2923), .CK(clk), .Q(new_AGEMA_signal_2924), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1741_s_current_state_reg ( .D(
        new_AGEMA_signal_2929), .CK(clk), .Q(new_AGEMA_signal_2930), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1743_s_current_state_reg ( .D(
        new_AGEMA_signal_2931), .CK(clk), .Q(new_AGEMA_signal_2932), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1751_s_current_state_reg ( .D(
        new_AGEMA_signal_2939), .CK(clk), .Q(new_AGEMA_signal_2940), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1755_s_current_state_reg ( .D(
        new_AGEMA_signal_2943), .CK(clk), .Q(new_AGEMA_signal_2944), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1757_s_current_state_reg ( .D(
        new_AGEMA_signal_2945), .CK(clk), .Q(new_AGEMA_signal_2946), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1759_s_current_state_reg ( .D(
        new_AGEMA_signal_2947), .CK(clk), .Q(new_AGEMA_signal_2948), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1765_s_current_state_reg ( .D(
        new_AGEMA_signal_2953), .CK(clk), .Q(new_AGEMA_signal_2954), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1767_s_current_state_reg ( .D(
        new_AGEMA_signal_2955), .CK(clk), .Q(new_AGEMA_signal_2956), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1775_s_current_state_reg ( .D(
        new_AGEMA_signal_2963), .CK(clk), .Q(new_AGEMA_signal_2964), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1779_s_current_state_reg ( .D(
        new_AGEMA_signal_2967), .CK(clk), .Q(new_AGEMA_signal_2968), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1781_s_current_state_reg ( .D(
        new_AGEMA_signal_2969), .CK(clk), .Q(new_AGEMA_signal_2970), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1783_s_current_state_reg ( .D(
        new_AGEMA_signal_2971), .CK(clk), .Q(new_AGEMA_signal_2972), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1789_s_current_state_reg ( .D(
        new_AGEMA_signal_2977), .CK(clk), .Q(new_AGEMA_signal_2978), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1791_s_current_state_reg ( .D(
        new_AGEMA_signal_2979), .CK(clk), .Q(new_AGEMA_signal_2980), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1799_s_current_state_reg ( .D(
        new_AGEMA_signal_2987), .CK(clk), .Q(new_AGEMA_signal_2988), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1803_s_current_state_reg ( .D(
        new_AGEMA_signal_2991), .CK(clk), .Q(new_AGEMA_signal_2992), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1805_s_current_state_reg ( .D(
        new_AGEMA_signal_2993), .CK(clk), .Q(new_AGEMA_signal_2994), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1807_s_current_state_reg ( .D(
        new_AGEMA_signal_2995), .CK(clk), .Q(new_AGEMA_signal_2996), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1813_s_current_state_reg ( .D(
        new_AGEMA_signal_3001), .CK(clk), .Q(new_AGEMA_signal_3002), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1815_s_current_state_reg ( .D(
        new_AGEMA_signal_3003), .CK(clk), .Q(new_AGEMA_signal_3004), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1823_s_current_state_reg ( .D(
        new_AGEMA_signal_3011), .CK(clk), .Q(new_AGEMA_signal_3012), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1827_s_current_state_reg ( .D(
        new_AGEMA_signal_3015), .CK(clk), .Q(new_AGEMA_signal_3016), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1829_s_current_state_reg ( .D(
        new_AGEMA_signal_3017), .CK(clk), .Q(new_AGEMA_signal_3018), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1831_s_current_state_reg ( .D(
        new_AGEMA_signal_3019), .CK(clk), .Q(new_AGEMA_signal_3020), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1837_s_current_state_reg ( .D(
        new_AGEMA_signal_3025), .CK(clk), .Q(new_AGEMA_signal_3026), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1839_s_current_state_reg ( .D(
        new_AGEMA_signal_3027), .CK(clk), .Q(new_AGEMA_signal_3028), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1847_s_current_state_reg ( .D(
        new_AGEMA_signal_3035), .CK(clk), .Q(new_AGEMA_signal_3036), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1851_s_current_state_reg ( .D(
        new_AGEMA_signal_3039), .CK(clk), .Q(new_AGEMA_signal_3040), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1853_s_current_state_reg ( .D(
        new_AGEMA_signal_3041), .CK(clk), .Q(new_AGEMA_signal_3042), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1855_s_current_state_reg ( .D(
        new_AGEMA_signal_3043), .CK(clk), .Q(new_AGEMA_signal_3044), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1861_s_current_state_reg ( .D(
        new_AGEMA_signal_3049), .CK(clk), .Q(new_AGEMA_signal_3050), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1863_s_current_state_reg ( .D(
        new_AGEMA_signal_3051), .CK(clk), .Q(new_AGEMA_signal_3052), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1871_s_current_state_reg ( .D(
        new_AGEMA_signal_3059), .CK(clk), .Q(new_AGEMA_signal_3060), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1875_s_current_state_reg ( .D(
        new_AGEMA_signal_3063), .CK(clk), .Q(new_AGEMA_signal_3064), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1877_s_current_state_reg ( .D(
        new_AGEMA_signal_3065), .CK(clk), .Q(new_AGEMA_signal_3066), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1879_s_current_state_reg ( .D(
        new_AGEMA_signal_3067), .CK(clk), .Q(new_AGEMA_signal_3068), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1885_s_current_state_reg ( .D(
        new_AGEMA_signal_3073), .CK(clk), .Q(new_AGEMA_signal_3074), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1887_s_current_state_reg ( .D(
        new_AGEMA_signal_3075), .CK(clk), .Q(new_AGEMA_signal_3076), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1895_s_current_state_reg ( .D(
        new_AGEMA_signal_3083), .CK(clk), .Q(new_AGEMA_signal_3084), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1899_s_current_state_reg ( .D(
        new_AGEMA_signal_3087), .CK(clk), .Q(new_AGEMA_signal_3088), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1901_s_current_state_reg ( .D(
        new_AGEMA_signal_3089), .CK(clk), .Q(new_AGEMA_signal_3090), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1903_s_current_state_reg ( .D(
        new_AGEMA_signal_3091), .CK(clk), .Q(new_AGEMA_signal_3092), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1909_s_current_state_reg ( .D(
        new_AGEMA_signal_3097), .CK(clk), .Q(new_AGEMA_signal_3098), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1911_s_current_state_reg ( .D(
        new_AGEMA_signal_3099), .CK(clk), .Q(new_AGEMA_signal_3100), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1919_s_current_state_reg ( .D(
        new_AGEMA_signal_3107), .CK(clk), .Q(new_AGEMA_signal_3108), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1923_s_current_state_reg ( .D(
        new_AGEMA_signal_3111), .CK(clk), .Q(new_AGEMA_signal_3112), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1925_s_current_state_reg ( .D(
        new_AGEMA_signal_3113), .CK(clk), .Q(new_AGEMA_signal_3114), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1927_s_current_state_reg ( .D(
        new_AGEMA_signal_3115), .CK(clk), .Q(new_AGEMA_signal_3116), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1933_s_current_state_reg ( .D(
        new_AGEMA_signal_3121), .CK(clk), .Q(new_AGEMA_signal_3122), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1935_s_current_state_reg ( .D(
        new_AGEMA_signal_3123), .CK(clk), .Q(new_AGEMA_signal_3124), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1943_s_current_state_reg ( .D(
        new_AGEMA_signal_3131), .CK(clk), .Q(new_AGEMA_signal_3132), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1947_s_current_state_reg ( .D(
        new_AGEMA_signal_3135), .CK(clk), .Q(new_AGEMA_signal_3136), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1949_s_current_state_reg ( .D(
        new_AGEMA_signal_3137), .CK(clk), .Q(new_AGEMA_signal_3138), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1951_s_current_state_reg ( .D(
        new_AGEMA_signal_3139), .CK(clk), .Q(new_AGEMA_signal_3140), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1957_s_current_state_reg ( .D(
        new_AGEMA_signal_3145), .CK(clk), .Q(new_AGEMA_signal_3146), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1959_s_current_state_reg ( .D(
        new_AGEMA_signal_3147), .CK(clk), .Q(new_AGEMA_signal_3148), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1967_s_current_state_reg ( .D(
        new_AGEMA_signal_3155), .CK(clk), .Q(new_AGEMA_signal_3156), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1971_s_current_state_reg ( .D(
        new_AGEMA_signal_3159), .CK(clk), .Q(new_AGEMA_signal_3160), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1973_s_current_state_reg ( .D(
        new_AGEMA_signal_3161), .CK(clk), .Q(new_AGEMA_signal_3162), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1975_s_current_state_reg ( .D(
        new_AGEMA_signal_3163), .CK(clk), .Q(new_AGEMA_signal_3164), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1981_s_current_state_reg ( .D(
        new_AGEMA_signal_3169), .CK(clk), .Q(new_AGEMA_signal_3170), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1983_s_current_state_reg ( .D(
        new_AGEMA_signal_3171), .CK(clk), .Q(new_AGEMA_signal_3172), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1991_s_current_state_reg ( .D(
        new_AGEMA_signal_3179), .CK(clk), .Q(new_AGEMA_signal_3180), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1995_s_current_state_reg ( .D(
        new_AGEMA_signal_3183), .CK(clk), .Q(new_AGEMA_signal_3184), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1997_s_current_state_reg ( .D(
        new_AGEMA_signal_3185), .CK(clk), .Q(new_AGEMA_signal_3186), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1999_s_current_state_reg ( .D(
        new_AGEMA_signal_3187), .CK(clk), .Q(new_AGEMA_signal_3188), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2005_s_current_state_reg ( .D(
        new_AGEMA_signal_3193), .CK(clk), .Q(new_AGEMA_signal_3194), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2007_s_current_state_reg ( .D(
        new_AGEMA_signal_3195), .CK(clk), .Q(new_AGEMA_signal_3196), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2015_s_current_state_reg ( .D(
        new_AGEMA_signal_3203), .CK(clk), .Q(new_AGEMA_signal_3204), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2019_s_current_state_reg ( .D(
        new_AGEMA_signal_3207), .CK(clk), .Q(new_AGEMA_signal_3208), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2021_s_current_state_reg ( .D(
        new_AGEMA_signal_3209), .CK(clk), .Q(new_AGEMA_signal_3210), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2023_s_current_state_reg ( .D(
        new_AGEMA_signal_3211), .CK(clk), .Q(new_AGEMA_signal_3212), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2029_s_current_state_reg ( .D(
        new_AGEMA_signal_3217), .CK(clk), .Q(new_AGEMA_signal_3218), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2031_s_current_state_reg ( .D(
        new_AGEMA_signal_3219), .CK(clk), .Q(new_AGEMA_signal_3220), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2039_s_current_state_reg ( .D(
        new_AGEMA_signal_3227), .CK(clk), .Q(new_AGEMA_signal_3228), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2043_s_current_state_reg ( .D(
        new_AGEMA_signal_3231), .CK(clk), .Q(new_AGEMA_signal_3232), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2045_s_current_state_reg ( .D(
        new_AGEMA_signal_3233), .CK(clk), .Q(new_AGEMA_signal_3234), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2047_s_current_state_reg ( .D(
        new_AGEMA_signal_3235), .CK(clk), .Q(new_AGEMA_signal_3236), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2053_s_current_state_reg ( .D(
        new_AGEMA_signal_3241), .CK(clk), .Q(new_AGEMA_signal_3242), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2055_s_current_state_reg ( .D(
        new_AGEMA_signal_3243), .CK(clk), .Q(new_AGEMA_signal_3244), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2063_s_current_state_reg ( .D(
        new_AGEMA_signal_3251), .CK(clk), .Q(new_AGEMA_signal_3252), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2067_s_current_state_reg ( .D(
        new_AGEMA_signal_3255), .CK(clk), .Q(new_AGEMA_signal_3256), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2069_s_current_state_reg ( .D(
        new_AGEMA_signal_3257), .CK(clk), .Q(new_AGEMA_signal_3258), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2071_s_current_state_reg ( .D(
        new_AGEMA_signal_3259), .CK(clk), .Q(new_AGEMA_signal_3260), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2077_s_current_state_reg ( .D(
        new_AGEMA_signal_3265), .CK(clk), .Q(new_AGEMA_signal_3266), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2079_s_current_state_reg ( .D(
        new_AGEMA_signal_3267), .CK(clk), .Q(new_AGEMA_signal_3268), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2087_s_current_state_reg ( .D(
        new_AGEMA_signal_3275), .CK(clk), .Q(new_AGEMA_signal_3276), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2091_s_current_state_reg ( .D(
        new_AGEMA_signal_3279), .CK(clk), .Q(new_AGEMA_signal_3280), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2093_s_current_state_reg ( .D(
        new_AGEMA_signal_3281), .CK(clk), .Q(new_AGEMA_signal_3282), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2095_s_current_state_reg ( .D(
        new_AGEMA_signal_3283), .CK(clk), .Q(new_AGEMA_signal_3284), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2099_s_current_state_reg ( .D(
        new_AGEMA_signal_3287), .CK(clk), .Q(new_AGEMA_signal_3288), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2103_s_current_state_reg ( .D(
        new_AGEMA_signal_3291), .CK(clk), .Q(new_AGEMA_signal_3292), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2107_s_current_state_reg ( .D(
        new_AGEMA_signal_3295), .CK(clk), .Q(new_AGEMA_signal_3296), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2111_s_current_state_reg ( .D(
        new_AGEMA_signal_3299), .CK(clk), .Q(new_AGEMA_signal_3300), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2115_s_current_state_reg ( .D(
        new_AGEMA_signal_3303), .CK(clk), .Q(new_AGEMA_signal_3304), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2119_s_current_state_reg ( .D(
        new_AGEMA_signal_3307), .CK(clk), .Q(new_AGEMA_signal_3308), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2123_s_current_state_reg ( .D(
        new_AGEMA_signal_3311), .CK(clk), .Q(new_AGEMA_signal_3312), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2127_s_current_state_reg ( .D(
        new_AGEMA_signal_3315), .CK(clk), .Q(new_AGEMA_signal_3316), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2131_s_current_state_reg ( .D(
        new_AGEMA_signal_3319), .CK(clk), .Q(new_AGEMA_signal_3320), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2135_s_current_state_reg ( .D(
        new_AGEMA_signal_3323), .CK(clk), .Q(new_AGEMA_signal_3324), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2139_s_current_state_reg ( .D(
        new_AGEMA_signal_3327), .CK(clk), .Q(new_AGEMA_signal_3328), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2143_s_current_state_reg ( .D(
        new_AGEMA_signal_3331), .CK(clk), .Q(new_AGEMA_signal_3332), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2147_s_current_state_reg ( .D(
        new_AGEMA_signal_3335), .CK(clk), .Q(new_AGEMA_signal_3336), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2151_s_current_state_reg ( .D(
        new_AGEMA_signal_3339), .CK(clk), .Q(new_AGEMA_signal_3340), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2155_s_current_state_reg ( .D(
        new_AGEMA_signal_3343), .CK(clk), .Q(new_AGEMA_signal_3344), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2159_s_current_state_reg ( .D(
        new_AGEMA_signal_3347), .CK(clk), .Q(new_AGEMA_signal_3348), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2163_s_current_state_reg ( .D(
        new_AGEMA_signal_3351), .CK(clk), .Q(new_AGEMA_signal_3352), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2167_s_current_state_reg ( .D(
        new_AGEMA_signal_3355), .CK(clk), .Q(new_AGEMA_signal_3356), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2171_s_current_state_reg ( .D(
        new_AGEMA_signal_3359), .CK(clk), .Q(new_AGEMA_signal_3360), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2175_s_current_state_reg ( .D(
        new_AGEMA_signal_3363), .CK(clk), .Q(new_AGEMA_signal_3364), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2179_s_current_state_reg ( .D(
        new_AGEMA_signal_3367), .CK(clk), .Q(new_AGEMA_signal_3368), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2183_s_current_state_reg ( .D(
        new_AGEMA_signal_3371), .CK(clk), .Q(new_AGEMA_signal_3372), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2187_s_current_state_reg ( .D(
        new_AGEMA_signal_3375), .CK(clk), .Q(new_AGEMA_signal_3376), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2191_s_current_state_reg ( .D(
        new_AGEMA_signal_3379), .CK(clk), .Q(new_AGEMA_signal_3380), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2195_s_current_state_reg ( .D(
        new_AGEMA_signal_3383), .CK(clk), .Q(new_AGEMA_signal_3384), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2199_s_current_state_reg ( .D(
        new_AGEMA_signal_3387), .CK(clk), .Q(new_AGEMA_signal_3388), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2203_s_current_state_reg ( .D(
        new_AGEMA_signal_3391), .CK(clk), .Q(new_AGEMA_signal_3392), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2207_s_current_state_reg ( .D(
        new_AGEMA_signal_3395), .CK(clk), .Q(new_AGEMA_signal_3396), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2211_s_current_state_reg ( .D(
        new_AGEMA_signal_3399), .CK(clk), .Q(new_AGEMA_signal_3400), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2215_s_current_state_reg ( .D(
        new_AGEMA_signal_3403), .CK(clk), .Q(new_AGEMA_signal_3404), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2219_s_current_state_reg ( .D(
        new_AGEMA_signal_3407), .CK(clk), .Q(new_AGEMA_signal_3408), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2223_s_current_state_reg ( .D(
        new_AGEMA_signal_3411), .CK(clk), .Q(new_AGEMA_signal_3412), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2227_s_current_state_reg ( .D(
        new_AGEMA_signal_3415), .CK(clk), .Q(new_AGEMA_signal_3416), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2231_s_current_state_reg ( .D(
        new_AGEMA_signal_3419), .CK(clk), .Q(new_AGEMA_signal_3420), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2235_s_current_state_reg ( .D(
        new_AGEMA_signal_3423), .CK(clk), .Q(new_AGEMA_signal_3424), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2239_s_current_state_reg ( .D(
        new_AGEMA_signal_3427), .CK(clk), .Q(new_AGEMA_signal_3428), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2241_s_current_state_reg ( .D(
        new_AGEMA_signal_3429), .CK(clk), .Q(new_AGEMA_signal_3430), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2243_s_current_state_reg ( .D(
        new_AGEMA_signal_3431), .CK(clk), .Q(new_AGEMA_signal_3432), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2245_s_current_state_reg ( .D(
        new_AGEMA_signal_3433), .CK(clk), .Q(new_AGEMA_signal_3434), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2247_s_current_state_reg ( .D(
        new_AGEMA_signal_3435), .CK(clk), .Q(new_AGEMA_signal_3436), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2249_s_current_state_reg ( .D(
        new_AGEMA_signal_3437), .CK(clk), .Q(new_AGEMA_signal_3438), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2251_s_current_state_reg ( .D(
        new_AGEMA_signal_3439), .CK(clk), .Q(new_AGEMA_signal_3440), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2253_s_current_state_reg ( .D(
        new_AGEMA_signal_3441), .CK(clk), .Q(new_AGEMA_signal_3442), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2255_s_current_state_reg ( .D(
        new_AGEMA_signal_3443), .CK(clk), .Q(new_AGEMA_signal_3444), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2257_s_current_state_reg ( .D(
        new_AGEMA_signal_3445), .CK(clk), .Q(new_AGEMA_signal_3446), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2259_s_current_state_reg ( .D(
        new_AGEMA_signal_3447), .CK(clk), .Q(new_AGEMA_signal_3448), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2261_s_current_state_reg ( .D(
        new_AGEMA_signal_3449), .CK(clk), .Q(new_AGEMA_signal_3450), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2263_s_current_state_reg ( .D(
        new_AGEMA_signal_3451), .CK(clk), .Q(new_AGEMA_signal_3452), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2265_s_current_state_reg ( .D(
        new_AGEMA_signal_3453), .CK(clk), .Q(new_AGEMA_signal_3454), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2267_s_current_state_reg ( .D(
        new_AGEMA_signal_3455), .CK(clk), .Q(new_AGEMA_signal_3456), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2269_s_current_state_reg ( .D(
        new_AGEMA_signal_3457), .CK(clk), .Q(new_AGEMA_signal_3458), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2271_s_current_state_reg ( .D(
        new_AGEMA_signal_3459), .CK(clk), .Q(new_AGEMA_signal_3460), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2273_s_current_state_reg ( .D(
        new_AGEMA_signal_3461), .CK(clk), .Q(new_AGEMA_signal_3462), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2275_s_current_state_reg ( .D(
        new_AGEMA_signal_3463), .CK(clk), .Q(new_AGEMA_signal_3464), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2277_s_current_state_reg ( .D(
        new_AGEMA_signal_3465), .CK(clk), .Q(new_AGEMA_signal_3466), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2279_s_current_state_reg ( .D(
        new_AGEMA_signal_3467), .CK(clk), .Q(new_AGEMA_signal_3468), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2281_s_current_state_reg ( .D(
        new_AGEMA_signal_3469), .CK(clk), .Q(new_AGEMA_signal_3470), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2283_s_current_state_reg ( .D(
        new_AGEMA_signal_3471), .CK(clk), .Q(new_AGEMA_signal_3472), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2285_s_current_state_reg ( .D(
        new_AGEMA_signal_3473), .CK(clk), .Q(new_AGEMA_signal_3474), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2287_s_current_state_reg ( .D(
        new_AGEMA_signal_3475), .CK(clk), .Q(new_AGEMA_signal_3476), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2289_s_current_state_reg ( .D(
        new_AGEMA_signal_3477), .CK(clk), .Q(new_AGEMA_signal_3478), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2291_s_current_state_reg ( .D(
        new_AGEMA_signal_3479), .CK(clk), .Q(new_AGEMA_signal_3480), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2293_s_current_state_reg ( .D(
        new_AGEMA_signal_3481), .CK(clk), .Q(new_AGEMA_signal_3482), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2295_s_current_state_reg ( .D(
        new_AGEMA_signal_3483), .CK(clk), .Q(new_AGEMA_signal_3484), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2297_s_current_state_reg ( .D(
        new_AGEMA_signal_3485), .CK(clk), .Q(new_AGEMA_signal_3486), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2299_s_current_state_reg ( .D(
        new_AGEMA_signal_3487), .CK(clk), .Q(new_AGEMA_signal_3488), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2301_s_current_state_reg ( .D(
        new_AGEMA_signal_3489), .CK(clk), .Q(new_AGEMA_signal_3490), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2303_s_current_state_reg ( .D(
        new_AGEMA_signal_3491), .CK(clk), .Q(new_AGEMA_signal_3492), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2305_s_current_state_reg ( .D(
        new_AGEMA_signal_3493), .CK(clk), .Q(new_AGEMA_signal_3494), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2307_s_current_state_reg ( .D(
        new_AGEMA_signal_3495), .CK(clk), .Q(new_AGEMA_signal_3496), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2309_s_current_state_reg ( .D(
        new_AGEMA_signal_3497), .CK(clk), .Q(new_AGEMA_signal_3498), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2311_s_current_state_reg ( .D(
        new_AGEMA_signal_3499), .CK(clk), .Q(new_AGEMA_signal_3500), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2313_s_current_state_reg ( .D(
        new_AGEMA_signal_3501), .CK(clk), .Q(new_AGEMA_signal_3502), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2315_s_current_state_reg ( .D(
        new_AGEMA_signal_3503), .CK(clk), .Q(new_AGEMA_signal_3504), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2317_s_current_state_reg ( .D(
        new_AGEMA_signal_3505), .CK(clk), .Q(new_AGEMA_signal_3506), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2319_s_current_state_reg ( .D(
        new_AGEMA_signal_3507), .CK(clk), .Q(new_AGEMA_signal_3508), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2321_s_current_state_reg ( .D(
        new_AGEMA_signal_3509), .CK(clk), .Q(new_AGEMA_signal_3510), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2323_s_current_state_reg ( .D(
        new_AGEMA_signal_3511), .CK(clk), .Q(new_AGEMA_signal_3512), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2325_s_current_state_reg ( .D(
        new_AGEMA_signal_3513), .CK(clk), .Q(new_AGEMA_signal_3514), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2327_s_current_state_reg ( .D(
        new_AGEMA_signal_3515), .CK(clk), .Q(new_AGEMA_signal_3516), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2329_s_current_state_reg ( .D(
        new_AGEMA_signal_3517), .CK(clk), .Q(new_AGEMA_signal_3518), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2331_s_current_state_reg ( .D(
        new_AGEMA_signal_3519), .CK(clk), .Q(new_AGEMA_signal_3520), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2333_s_current_state_reg ( .D(
        new_AGEMA_signal_3521), .CK(clk), .Q(new_AGEMA_signal_3522), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2335_s_current_state_reg ( .D(
        new_AGEMA_signal_3523), .CK(clk), .Q(new_AGEMA_signal_3524), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2337_s_current_state_reg ( .D(
        new_AGEMA_signal_3525), .CK(clk), .Q(new_AGEMA_signal_3526), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2339_s_current_state_reg ( .D(
        new_AGEMA_signal_3527), .CK(clk), .Q(new_AGEMA_signal_3528), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2341_s_current_state_reg ( .D(
        new_AGEMA_signal_3529), .CK(clk), .Q(new_AGEMA_signal_3530), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2343_s_current_state_reg ( .D(
        new_AGEMA_signal_3531), .CK(clk), .Q(new_AGEMA_signal_3532), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2345_s_current_state_reg ( .D(
        new_AGEMA_signal_3533), .CK(clk), .Q(new_AGEMA_signal_3534), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2347_s_current_state_reg ( .D(
        new_AGEMA_signal_3535), .CK(clk), .Q(new_AGEMA_signal_3536), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2349_s_current_state_reg ( .D(
        new_AGEMA_signal_3537), .CK(clk), .Q(new_AGEMA_signal_3538), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2351_s_current_state_reg ( .D(
        new_AGEMA_signal_3539), .CK(clk), .Q(new_AGEMA_signal_3540), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2353_s_current_state_reg ( .D(
        new_AGEMA_signal_3541), .CK(clk), .Q(new_AGEMA_signal_3542), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2355_s_current_state_reg ( .D(
        new_AGEMA_signal_3543), .CK(clk), .Q(new_AGEMA_signal_3544), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2357_s_current_state_reg ( .D(
        new_AGEMA_signal_3545), .CK(clk), .Q(new_AGEMA_signal_3546), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2359_s_current_state_reg ( .D(
        new_AGEMA_signal_3547), .CK(clk), .Q(new_AGEMA_signal_3548), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2361_s_current_state_reg ( .D(
        new_AGEMA_signal_3549), .CK(clk), .Q(new_AGEMA_signal_3550), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2363_s_current_state_reg ( .D(
        new_AGEMA_signal_3551), .CK(clk), .Q(new_AGEMA_signal_3552), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2365_s_current_state_reg ( .D(
        new_AGEMA_signal_3553), .CK(clk), .Q(new_AGEMA_signal_3554), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2367_s_current_state_reg ( .D(
        new_AGEMA_signal_3555), .CK(clk), .Q(new_AGEMA_signal_3556), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2371_s_current_state_reg ( .D(
        new_AGEMA_signal_3559), .CK(clk), .Q(new_AGEMA_signal_3560), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2375_s_current_state_reg ( .D(
        new_AGEMA_signal_3563), .CK(clk), .Q(new_AGEMA_signal_3564), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2379_s_current_state_reg ( .D(
        new_AGEMA_signal_3567), .CK(clk), .Q(new_AGEMA_signal_3568), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2383_s_current_state_reg ( .D(
        new_AGEMA_signal_3571), .CK(clk), .Q(new_AGEMA_signal_3572), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2387_s_current_state_reg ( .D(
        new_AGEMA_signal_3575), .CK(clk), .Q(new_AGEMA_signal_3576), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2391_s_current_state_reg ( .D(
        new_AGEMA_signal_3579), .CK(clk), .Q(new_AGEMA_signal_3580), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2395_s_current_state_reg ( .D(
        new_AGEMA_signal_3583), .CK(clk), .Q(new_AGEMA_signal_3584), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2399_s_current_state_reg ( .D(
        new_AGEMA_signal_3587), .CK(clk), .Q(new_AGEMA_signal_3588), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2403_s_current_state_reg ( .D(
        new_AGEMA_signal_3591), .CK(clk), .Q(new_AGEMA_signal_3592), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2407_s_current_state_reg ( .D(
        new_AGEMA_signal_3595), .CK(clk), .Q(new_AGEMA_signal_3596), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2411_s_current_state_reg ( .D(
        new_AGEMA_signal_3599), .CK(clk), .Q(new_AGEMA_signal_3600), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2415_s_current_state_reg ( .D(
        new_AGEMA_signal_3603), .CK(clk), .Q(new_AGEMA_signal_3604), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2419_s_current_state_reg ( .D(
        new_AGEMA_signal_3607), .CK(clk), .Q(new_AGEMA_signal_3608), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2423_s_current_state_reg ( .D(
        new_AGEMA_signal_3611), .CK(clk), .Q(new_AGEMA_signal_3612), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2427_s_current_state_reg ( .D(
        new_AGEMA_signal_3615), .CK(clk), .Q(new_AGEMA_signal_3616), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2431_s_current_state_reg ( .D(
        new_AGEMA_signal_3619), .CK(clk), .Q(new_AGEMA_signal_3620), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2435_s_current_state_reg ( .D(
        new_AGEMA_signal_3623), .CK(clk), .Q(new_AGEMA_signal_3624), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2439_s_current_state_reg ( .D(
        new_AGEMA_signal_3627), .CK(clk), .Q(new_AGEMA_signal_3628), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2443_s_current_state_reg ( .D(
        new_AGEMA_signal_3631), .CK(clk), .Q(new_AGEMA_signal_3632), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2447_s_current_state_reg ( .D(
        new_AGEMA_signal_3635), .CK(clk), .Q(new_AGEMA_signal_3636), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2451_s_current_state_reg ( .D(
        new_AGEMA_signal_3639), .CK(clk), .Q(new_AGEMA_signal_3640), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2455_s_current_state_reg ( .D(
        new_AGEMA_signal_3643), .CK(clk), .Q(new_AGEMA_signal_3644), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2459_s_current_state_reg ( .D(
        new_AGEMA_signal_3647), .CK(clk), .Q(new_AGEMA_signal_3648), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2463_s_current_state_reg ( .D(
        new_AGEMA_signal_3651), .CK(clk), .Q(new_AGEMA_signal_3652), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2467_s_current_state_reg ( .D(
        new_AGEMA_signal_3655), .CK(clk), .Q(new_AGEMA_signal_3656), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2471_s_current_state_reg ( .D(
        new_AGEMA_signal_3659), .CK(clk), .Q(new_AGEMA_signal_3660), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2475_s_current_state_reg ( .D(
        new_AGEMA_signal_3663), .CK(clk), .Q(new_AGEMA_signal_3664), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2479_s_current_state_reg ( .D(
        new_AGEMA_signal_3667), .CK(clk), .Q(new_AGEMA_signal_3668), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2483_s_current_state_reg ( .D(
        new_AGEMA_signal_3671), .CK(clk), .Q(new_AGEMA_signal_3672), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2487_s_current_state_reg ( .D(
        new_AGEMA_signal_3675), .CK(clk), .Q(new_AGEMA_signal_3676), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2491_s_current_state_reg ( .D(
        new_AGEMA_signal_3679), .CK(clk), .Q(new_AGEMA_signal_3680), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2495_s_current_state_reg ( .D(
        new_AGEMA_signal_3683), .CK(clk), .Q(new_AGEMA_signal_3684), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2499_s_current_state_reg ( .D(
        new_AGEMA_signal_3687), .CK(clk), .Q(new_AGEMA_signal_3688), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2503_s_current_state_reg ( .D(
        new_AGEMA_signal_3691), .CK(clk), .Q(new_AGEMA_signal_3692), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2507_s_current_state_reg ( .D(
        new_AGEMA_signal_3695), .CK(clk), .Q(new_AGEMA_signal_3696), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2511_s_current_state_reg ( .D(
        new_AGEMA_signal_3699), .CK(clk), .Q(new_AGEMA_signal_3700), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2515_s_current_state_reg ( .D(
        new_AGEMA_signal_3703), .CK(clk), .Q(new_AGEMA_signal_3704), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2519_s_current_state_reg ( .D(
        new_AGEMA_signal_3707), .CK(clk), .Q(new_AGEMA_signal_3708), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2523_s_current_state_reg ( .D(
        new_AGEMA_signal_3711), .CK(clk), .Q(new_AGEMA_signal_3712), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2527_s_current_state_reg ( .D(
        new_AGEMA_signal_3715), .CK(clk), .Q(new_AGEMA_signal_3716), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2531_s_current_state_reg ( .D(
        new_AGEMA_signal_3719), .CK(clk), .Q(new_AGEMA_signal_3720), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2535_s_current_state_reg ( .D(
        new_AGEMA_signal_3723), .CK(clk), .Q(new_AGEMA_signal_3724), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2539_s_current_state_reg ( .D(
        new_AGEMA_signal_3727), .CK(clk), .Q(new_AGEMA_signal_3728), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2543_s_current_state_reg ( .D(
        new_AGEMA_signal_3731), .CK(clk), .Q(new_AGEMA_signal_3732), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2547_s_current_state_reg ( .D(
        new_AGEMA_signal_3735), .CK(clk), .Q(new_AGEMA_signal_3736), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2551_s_current_state_reg ( .D(
        new_AGEMA_signal_3739), .CK(clk), .Q(new_AGEMA_signal_3740), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2555_s_current_state_reg ( .D(
        new_AGEMA_signal_3743), .CK(clk), .Q(new_AGEMA_signal_3744), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2559_s_current_state_reg ( .D(
        new_AGEMA_signal_3747), .CK(clk), .Q(new_AGEMA_signal_3748), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2563_s_current_state_reg ( .D(
        new_AGEMA_signal_3751), .CK(clk), .Q(new_AGEMA_signal_3752), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2567_s_current_state_reg ( .D(
        new_AGEMA_signal_3755), .CK(clk), .Q(new_AGEMA_signal_3756), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2571_s_current_state_reg ( .D(
        new_AGEMA_signal_3759), .CK(clk), .Q(new_AGEMA_signal_3760), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2575_s_current_state_reg ( .D(
        new_AGEMA_signal_3763), .CK(clk), .Q(new_AGEMA_signal_3764), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2579_s_current_state_reg ( .D(
        new_AGEMA_signal_3767), .CK(clk), .Q(new_AGEMA_signal_3768), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2583_s_current_state_reg ( .D(
        new_AGEMA_signal_3771), .CK(clk), .Q(new_AGEMA_signal_3772), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2587_s_current_state_reg ( .D(
        new_AGEMA_signal_3775), .CK(clk), .Q(new_AGEMA_signal_3776), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2591_s_current_state_reg ( .D(
        new_AGEMA_signal_3779), .CK(clk), .Q(new_AGEMA_signal_3780), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2595_s_current_state_reg ( .D(
        new_AGEMA_signal_3783), .CK(clk), .Q(new_AGEMA_signal_3784), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2599_s_current_state_reg ( .D(
        new_AGEMA_signal_3787), .CK(clk), .Q(new_AGEMA_signal_3788), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2603_s_current_state_reg ( .D(
        new_AGEMA_signal_3791), .CK(clk), .Q(new_AGEMA_signal_3792), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2607_s_current_state_reg ( .D(
        new_AGEMA_signal_3795), .CK(clk), .Q(new_AGEMA_signal_3796), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2611_s_current_state_reg ( .D(
        new_AGEMA_signal_3799), .CK(clk), .Q(new_AGEMA_signal_3800), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2615_s_current_state_reg ( .D(
        new_AGEMA_signal_3803), .CK(clk), .Q(new_AGEMA_signal_3804), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2619_s_current_state_reg ( .D(
        new_AGEMA_signal_3807), .CK(clk), .Q(new_AGEMA_signal_3808), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2623_s_current_state_reg ( .D(
        new_AGEMA_signal_3811), .CK(clk), .Q(new_AGEMA_signal_3812), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2627_s_current_state_reg ( .D(
        new_AGEMA_signal_3815), .CK(clk), .Q(new_AGEMA_signal_3816), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2631_s_current_state_reg ( .D(
        new_AGEMA_signal_3819), .CK(clk), .Q(new_AGEMA_signal_3820), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2635_s_current_state_reg ( .D(
        new_AGEMA_signal_3823), .CK(clk), .Q(new_AGEMA_signal_3824), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2639_s_current_state_reg ( .D(
        new_AGEMA_signal_3827), .CK(clk), .Q(new_AGEMA_signal_3828), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2643_s_current_state_reg ( .D(
        new_AGEMA_signal_3831), .CK(clk), .Q(new_AGEMA_signal_3832), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2647_s_current_state_reg ( .D(
        new_AGEMA_signal_3835), .CK(clk), .Q(new_AGEMA_signal_3836), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2651_s_current_state_reg ( .D(
        new_AGEMA_signal_3839), .CK(clk), .Q(new_AGEMA_signal_3840), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2655_s_current_state_reg ( .D(
        new_AGEMA_signal_3843), .CK(clk), .Q(new_AGEMA_signal_3844), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2659_s_current_state_reg ( .D(
        new_AGEMA_signal_3847), .CK(clk), .Q(new_AGEMA_signal_3848), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2663_s_current_state_reg ( .D(
        new_AGEMA_signal_3851), .CK(clk), .Q(new_AGEMA_signal_3852), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2667_s_current_state_reg ( .D(
        new_AGEMA_signal_3855), .CK(clk), .Q(new_AGEMA_signal_3856), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2671_s_current_state_reg ( .D(
        new_AGEMA_signal_3859), .CK(clk), .Q(new_AGEMA_signal_3860), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2675_s_current_state_reg ( .D(
        new_AGEMA_signal_3863), .CK(clk), .Q(new_AGEMA_signal_3864), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2679_s_current_state_reg ( .D(
        new_AGEMA_signal_3867), .CK(clk), .Q(new_AGEMA_signal_3868), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2683_s_current_state_reg ( .D(
        new_AGEMA_signal_3871), .CK(clk), .Q(new_AGEMA_signal_3872), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2687_s_current_state_reg ( .D(
        new_AGEMA_signal_3875), .CK(clk), .Q(new_AGEMA_signal_3876), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2691_s_current_state_reg ( .D(
        new_AGEMA_signal_3879), .CK(clk), .Q(new_AGEMA_signal_3880), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2695_s_current_state_reg ( .D(
        new_AGEMA_signal_3883), .CK(clk), .Q(new_AGEMA_signal_3884), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2699_s_current_state_reg ( .D(
        new_AGEMA_signal_3887), .CK(clk), .Q(new_AGEMA_signal_3888), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2703_s_current_state_reg ( .D(
        new_AGEMA_signal_3891), .CK(clk), .Q(new_AGEMA_signal_3892), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2707_s_current_state_reg ( .D(
        new_AGEMA_signal_3895), .CK(clk), .Q(new_AGEMA_signal_3896), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2711_s_current_state_reg ( .D(
        new_AGEMA_signal_3899), .CK(clk), .Q(new_AGEMA_signal_3900), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2715_s_current_state_reg ( .D(
        new_AGEMA_signal_3903), .CK(clk), .Q(new_AGEMA_signal_3904), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2719_s_current_state_reg ( .D(
        new_AGEMA_signal_3907), .CK(clk), .Q(new_AGEMA_signal_3908), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2723_s_current_state_reg ( .D(
        new_AGEMA_signal_3911), .CK(clk), .Q(new_AGEMA_signal_3912), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2727_s_current_state_reg ( .D(
        new_AGEMA_signal_3915), .CK(clk), .Q(new_AGEMA_signal_3916), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2731_s_current_state_reg ( .D(
        new_AGEMA_signal_3919), .CK(clk), .Q(new_AGEMA_signal_3920), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2735_s_current_state_reg ( .D(
        new_AGEMA_signal_3923), .CK(clk), .Q(new_AGEMA_signal_3924), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2739_s_current_state_reg ( .D(
        new_AGEMA_signal_3927), .CK(clk), .Q(new_AGEMA_signal_3928), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2743_s_current_state_reg ( .D(
        new_AGEMA_signal_3931), .CK(clk), .Q(new_AGEMA_signal_3932), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2747_s_current_state_reg ( .D(
        new_AGEMA_signal_3935), .CK(clk), .Q(new_AGEMA_signal_3936), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2751_s_current_state_reg ( .D(
        new_AGEMA_signal_3939), .CK(clk), .Q(new_AGEMA_signal_3940), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2755_s_current_state_reg ( .D(
        new_AGEMA_signal_3943), .CK(clk), .Q(new_AGEMA_signal_3944), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2759_s_current_state_reg ( .D(
        new_AGEMA_signal_3947), .CK(clk), .Q(new_AGEMA_signal_3948), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2763_s_current_state_reg ( .D(
        new_AGEMA_signal_3951), .CK(clk), .Q(new_AGEMA_signal_3952), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2767_s_current_state_reg ( .D(
        new_AGEMA_signal_3955), .CK(clk), .Q(new_AGEMA_signal_3956), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2771_s_current_state_reg ( .D(
        new_AGEMA_signal_3959), .CK(clk), .Q(new_AGEMA_signal_3960), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2775_s_current_state_reg ( .D(
        new_AGEMA_signal_3963), .CK(clk), .Q(new_AGEMA_signal_3964), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2779_s_current_state_reg ( .D(
        new_AGEMA_signal_3967), .CK(clk), .Q(new_AGEMA_signal_3968), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2783_s_current_state_reg ( .D(
        new_AGEMA_signal_3971), .CK(clk), .Q(new_AGEMA_signal_3972), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2787_s_current_state_reg ( .D(
        new_AGEMA_signal_3975), .CK(clk), .Q(new_AGEMA_signal_3976), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2791_s_current_state_reg ( .D(
        new_AGEMA_signal_3979), .CK(clk), .Q(new_AGEMA_signal_3980), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2795_s_current_state_reg ( .D(
        new_AGEMA_signal_3983), .CK(clk), .Q(new_AGEMA_signal_3984), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2799_s_current_state_reg ( .D(
        new_AGEMA_signal_3987), .CK(clk), .Q(new_AGEMA_signal_3988), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2803_s_current_state_reg ( .D(
        new_AGEMA_signal_3991), .CK(clk), .Q(new_AGEMA_signal_3992), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2807_s_current_state_reg ( .D(
        new_AGEMA_signal_3995), .CK(clk), .Q(new_AGEMA_signal_3996), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2811_s_current_state_reg ( .D(
        new_AGEMA_signal_3999), .CK(clk), .Q(new_AGEMA_signal_4000), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2815_s_current_state_reg ( .D(
        new_AGEMA_signal_4003), .CK(clk), .Q(new_AGEMA_signal_4004), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2819_s_current_state_reg ( .D(
        new_AGEMA_signal_4007), .CK(clk), .Q(new_AGEMA_signal_4008), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2823_s_current_state_reg ( .D(
        new_AGEMA_signal_4011), .CK(clk), .Q(new_AGEMA_signal_4012), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2827_s_current_state_reg ( .D(
        new_AGEMA_signal_4015), .CK(clk), .Q(new_AGEMA_signal_4016), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2831_s_current_state_reg ( .D(
        new_AGEMA_signal_4019), .CK(clk), .Q(new_AGEMA_signal_4020), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2835_s_current_state_reg ( .D(
        new_AGEMA_signal_4023), .CK(clk), .Q(new_AGEMA_signal_4024), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2839_s_current_state_reg ( .D(
        new_AGEMA_signal_4027), .CK(clk), .Q(new_AGEMA_signal_4028), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2843_s_current_state_reg ( .D(
        new_AGEMA_signal_4031), .CK(clk), .Q(new_AGEMA_signal_4032), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2847_s_current_state_reg ( .D(
        new_AGEMA_signal_4035), .CK(clk), .Q(new_AGEMA_signal_4036), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2851_s_current_state_reg ( .D(
        new_AGEMA_signal_4039), .CK(clk), .Q(new_AGEMA_signal_4040), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2855_s_current_state_reg ( .D(
        new_AGEMA_signal_4043), .CK(clk), .Q(new_AGEMA_signal_4044), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2859_s_current_state_reg ( .D(
        new_AGEMA_signal_4047), .CK(clk), .Q(new_AGEMA_signal_4048), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2863_s_current_state_reg ( .D(
        new_AGEMA_signal_4051), .CK(clk), .Q(new_AGEMA_signal_4052), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2867_s_current_state_reg ( .D(
        new_AGEMA_signal_4055), .CK(clk), .Q(new_AGEMA_signal_4056), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2871_s_current_state_reg ( .D(
        new_AGEMA_signal_4059), .CK(clk), .Q(new_AGEMA_signal_4060), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2875_s_current_state_reg ( .D(
        new_AGEMA_signal_4063), .CK(clk), .Q(new_AGEMA_signal_4064), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2879_s_current_state_reg ( .D(
        new_AGEMA_signal_4067), .CK(clk), .Q(new_AGEMA_signal_4068), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2883_s_current_state_reg ( .D(
        new_AGEMA_signal_4071), .CK(clk), .Q(new_AGEMA_signal_4072), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2887_s_current_state_reg ( .D(
        new_AGEMA_signal_4075), .CK(clk), .Q(new_AGEMA_signal_4076), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2891_s_current_state_reg ( .D(
        new_AGEMA_signal_4079), .CK(clk), .Q(new_AGEMA_signal_4080), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2895_s_current_state_reg ( .D(
        new_AGEMA_signal_4083), .CK(clk), .Q(new_AGEMA_signal_4084), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2899_s_current_state_reg ( .D(
        new_AGEMA_signal_4087), .CK(clk), .Q(new_AGEMA_signal_4088), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2903_s_current_state_reg ( .D(
        new_AGEMA_signal_4091), .CK(clk), .Q(new_AGEMA_signal_4092), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3430), .CK(clk), .Q(Ciphertext_s0[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3432), .CK(clk), .Q(Ciphertext_s1[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3434), .CK(clk), .Q(Ciphertext_s0[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3436), .CK(clk), .Q(Ciphertext_s1[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[61]), .CK(clk), .Q(Ciphertext_s0[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2124), .CK(clk), .Q(Ciphertext_s1[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[60]), .CK(clk), .Q(Ciphertext_s0[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2115), .CK(clk), .Q(Ciphertext_s1[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3438), .CK(clk), .Q(Ciphertext_s0[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3440), .CK(clk), .Q(Ciphertext_s1[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3442), .CK(clk), .Q(Ciphertext_s0[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3444), .CK(clk), .Q(Ciphertext_s1[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[57]), .CK(clk), .Q(Ciphertext_s0[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2101), .CK(clk), .Q(Ciphertext_s1[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[56]), .CK(clk), .Q(Ciphertext_s0[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2058), .CK(clk), .Q(Ciphertext_s1[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3446), .CK(clk), .Q(Ciphertext_s0[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3448), .CK(clk), .Q(Ciphertext_s1[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3450), .CK(clk), .Q(Ciphertext_s0[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3452), .CK(clk), .Q(Ciphertext_s1[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[53]), .CK(clk), .Q(Ciphertext_s0[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2099), .CK(clk), .Q(Ciphertext_s1[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[52]), .CK(clk), .Q(Ciphertext_s0[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2056), .CK(clk), .Q(Ciphertext_s1[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3454), .CK(clk), .Q(Ciphertext_s0[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3456), .CK(clk), .Q(Ciphertext_s1[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3458), .CK(clk), .Q(Ciphertext_s0[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3460), .CK(clk), .Q(Ciphertext_s1[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[49]), .CK(clk), .Q(Ciphertext_s0[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2097), .CK(clk), .Q(Ciphertext_s1[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[48]), .CK(clk), .Q(Ciphertext_s0[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2054), .CK(clk), .Q(Ciphertext_s1[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3462), .CK(clk), .Q(Ciphertext_s0[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3464), .CK(clk), .Q(Ciphertext_s1[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3466), .CK(clk), .Q(Ciphertext_s0[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3468), .CK(clk), .Q(Ciphertext_s1[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[45]), .CK(clk), .Q(Ciphertext_s0[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2095), .CK(clk), .Q(Ciphertext_s1[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[44]), .CK(clk), .Q(Ciphertext_s0[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2052), .CK(clk), .Q(Ciphertext_s1[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3470), .CK(clk), .Q(Ciphertext_s0[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3472), .CK(clk), .Q(Ciphertext_s1[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3474), .CK(clk), .Q(Ciphertext_s0[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3476), .CK(clk), .Q(Ciphertext_s1[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[41]), .CK(clk), .Q(Ciphertext_s0[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1998), .CK(clk), .Q(Ciphertext_s1[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[40]), .CK(clk), .Q(Ciphertext_s0[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1938), .CK(clk), .Q(Ciphertext_s1[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3478), .CK(clk), .Q(Ciphertext_s0[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3480), .CK(clk), .Q(Ciphertext_s1[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3482), .CK(clk), .Q(Ciphertext_s0[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3484), .CK(clk), .Q(Ciphertext_s1[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[37]), .CK(clk), .Q(Ciphertext_s0[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1996), .CK(clk), .Q(Ciphertext_s1[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[36]), .CK(clk), .Q(Ciphertext_s0[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1936), .CK(clk), .Q(Ciphertext_s1[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3486), .CK(clk), .Q(Ciphertext_s0[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3488), .CK(clk), .Q(Ciphertext_s1[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3490), .CK(clk), .Q(Ciphertext_s0[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3492), .CK(clk), .Q(Ciphertext_s1[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[33]), .CK(clk), .Q(Ciphertext_s0[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1994), .CK(clk), .Q(Ciphertext_s1[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[32]), .CK(clk), .Q(Ciphertext_s0[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1934), .CK(clk), .Q(Ciphertext_s1[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3494), .CK(clk), .Q(Ciphertext_s0[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3496), .CK(clk), .Q(Ciphertext_s1[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3498), .CK(clk), .Q(Ciphertext_s0[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3500), .CK(clk), .Q(Ciphertext_s1[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[29]), .CK(clk), .Q(Ciphertext_s0[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2093), .CK(clk), .Q(Ciphertext_s1[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[28]), .CK(clk), .Q(Ciphertext_s0[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2050), .CK(clk), .Q(Ciphertext_s1[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3502), .CK(clk), .Q(Ciphertext_s0[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3504), .CK(clk), .Q(Ciphertext_s1[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3506), .CK(clk), .Q(Ciphertext_s0[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3508), .CK(clk), .Q(Ciphertext_s1[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[25]), .CK(clk), .Q(Ciphertext_s0[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2122), .CK(clk), .Q(Ciphertext_s1[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[24]), .CK(clk), .Q(Ciphertext_s0[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2113), .CK(clk), .Q(Ciphertext_s1[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3510), .CK(clk), .Q(Ciphertext_s0[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3512), .CK(clk), .Q(Ciphertext_s1[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3514), .CK(clk), .Q(Ciphertext_s0[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3516), .CK(clk), .Q(Ciphertext_s1[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[21]), .CK(clk), .Q(Ciphertext_s0[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2089), .CK(clk), .Q(Ciphertext_s1[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[20]), .CK(clk), .Q(Ciphertext_s0[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2046), .CK(clk), .Q(Ciphertext_s1[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3518), .CK(clk), .Q(Ciphertext_s0[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3520), .CK(clk), .Q(Ciphertext_s1[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3522), .CK(clk), .Q(Ciphertext_s0[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3524), .CK(clk), .Q(Ciphertext_s1[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[17]), .CK(clk), .Q(Ciphertext_s0[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2087), .CK(clk), .Q(Ciphertext_s1[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[16]), .CK(clk), .Q(Ciphertext_s0[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2044), .CK(clk), .Q(Ciphertext_s1[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3526), .CK(clk), .Q(Ciphertext_s0[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3528), .CK(clk), .Q(Ciphertext_s1[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3530), .CK(clk), .Q(Ciphertext_s0[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3532), .CK(clk), .Q(Ciphertext_s1[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[13]), .CK(clk), .Q(Ciphertext_s0[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2120), .CK(clk), .Q(Ciphertext_s1[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[12]), .CK(clk), .Q(Ciphertext_s0[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2111), .CK(clk), .Q(Ciphertext_s1[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3534), .CK(clk), .Q(Ciphertext_s0[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3536), .CK(clk), .Q(Ciphertext_s1[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3538), .CK(clk), .Q(Ciphertext_s0[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3540), .CK(clk), .Q(Ciphertext_s1[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[9]), .CK(clk), .Q(Ciphertext_s0[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2083), .CK(clk), .Q(Ciphertext_s1[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[8]), .CK(clk), .Q(Ciphertext_s0[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2040), .CK(clk), .Q(Ciphertext_s1[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3542), .CK(clk), .Q(Ciphertext_s0[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3544), .CK(clk), .Q(Ciphertext_s1[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3546), .CK(clk), .Q(Ciphertext_s0[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3548), .CK(clk), .Q(Ciphertext_s1[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[5]), .CK(clk), .Q(Ciphertext_s0[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2081), .CK(clk), .Q(Ciphertext_s1[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[4]), .CK(clk), .Q(Ciphertext_s0[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2038), .CK(clk), .Q(Ciphertext_s1[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3550), .CK(clk), .Q(Ciphertext_s0[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3552), .CK(clk), .Q(Ciphertext_s1[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3554), .CK(clk), .Q(Ciphertext_s0[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3556), .CK(clk), .Q(Ciphertext_s1[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[1]), .CK(clk), .Q(Ciphertext_s0[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2079), .CK(clk), .Q(Ciphertext_s1[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[0]), .CK(clk), .Q(Ciphertext_s0[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2036), .CK(clk), .Q(Ciphertext_s1[0]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3560), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[31]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3564), .CK(clk), .Q(new_AGEMA_signal_1353), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3568), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[30]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3572), .CK(clk), .Q(new_AGEMA_signal_1350), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3576), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[29]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3580), .CK(clk), .Q(new_AGEMA_signal_1347), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3584), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[28]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3588), .CK(clk), .Q(new_AGEMA_signal_1344), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3592), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[27]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3596), .CK(clk), .Q(new_AGEMA_signal_1341), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3600), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[26]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3604), .CK(clk), .Q(new_AGEMA_signal_1338), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3608), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[25]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3612), .CK(clk), .Q(new_AGEMA_signal_1335), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3616), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[24]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3620), .CK(clk), .Q(new_AGEMA_signal_1332), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3624), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[23]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3628), .CK(clk), .Q(new_AGEMA_signal_1329), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3632), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[22]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3636), .CK(clk), .Q(new_AGEMA_signal_1326), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3640), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[21]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3644), .CK(clk), .Q(new_AGEMA_signal_1323), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3648), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[20]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3652), .CK(clk), .Q(new_AGEMA_signal_1320), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3656), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[19]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3660), .CK(clk), .Q(new_AGEMA_signal_1317), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3664), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[18]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3668), .CK(clk), .Q(new_AGEMA_signal_1314), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3672), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[17]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3676), .CK(clk), .Q(new_AGEMA_signal_1311), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3680), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[16]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3684), .CK(clk), .Q(new_AGEMA_signal_1308), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3688), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[15]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3692), .CK(clk), .Q(new_AGEMA_signal_1305), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3696), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[14]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3700), .CK(clk), .Q(new_AGEMA_signal_1302), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3704), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[13]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3708), .CK(clk), .Q(new_AGEMA_signal_1299), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3712), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[12]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3716), .CK(clk), .Q(new_AGEMA_signal_1296), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3720), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[11]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3724), .CK(clk), .Q(new_AGEMA_signal_1293), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3728), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[10]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3732), .CK(clk), .Q(new_AGEMA_signal_1290), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3736), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[9]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3740), .CK(clk), .Q(new_AGEMA_signal_1287), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3744), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[8]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3748), .CK(clk), .Q(new_AGEMA_signal_1284), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3752), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[7]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3756), .CK(clk), .Q(new_AGEMA_signal_1281), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3760), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[6]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3764), .CK(clk), .Q(new_AGEMA_signal_1278), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3768), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[5]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3772), .CK(clk), .Q(new_AGEMA_signal_1275), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3776), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[4]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3780), .CK(clk), .Q(new_AGEMA_signal_1272), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3784), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[3]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3788), .CK(clk), .Q(new_AGEMA_signal_1269), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3792), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[2]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3796), .CK(clk), .Q(new_AGEMA_signal_1266), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3800), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[1]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3804), .CK(clk), .Q(new_AGEMA_signal_1263), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3808), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[0]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3812), .CK(clk), .Q(new_AGEMA_signal_1260), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3816), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[55]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3820), .CK(clk), .Q(new_AGEMA_signal_1425), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3824), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[54]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3828), .CK(clk), .Q(new_AGEMA_signal_1422), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3832), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[53]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3836), .CK(clk), .Q(new_AGEMA_signal_1419), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3840), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[52]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3844), .CK(clk), .Q(new_AGEMA_signal_1416), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3848), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[63]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3852), .CK(clk), .Q(new_AGEMA_signal_1449), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3856), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[62]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3860), .CK(clk), .Q(new_AGEMA_signal_1446), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3864), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[61]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3868), .CK(clk), .Q(new_AGEMA_signal_1443), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3872), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[60]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3876), .CK(clk), .Q(new_AGEMA_signal_1440), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3880), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[47]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3884), .CK(clk), .Q(new_AGEMA_signal_1401), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3888), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[46]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3892), .CK(clk), .Q(new_AGEMA_signal_1398), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3896), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[45]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3900), .CK(clk), .Q(new_AGEMA_signal_1395), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3904), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[44]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3908), .CK(clk), .Q(new_AGEMA_signal_1392), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3912), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[35]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3916), .CK(clk), .Q(new_AGEMA_signal_1365), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3920), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[34]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3924), .CK(clk), .Q(new_AGEMA_signal_1362), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3928), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[33]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3932), .CK(clk), .Q(new_AGEMA_signal_1359), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3936), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[32]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3940), .CK(clk), .Q(new_AGEMA_signal_1356), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3944), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[39]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3948), .CK(clk), .Q(new_AGEMA_signal_1377), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3952), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[38]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3956), .CK(clk), .Q(new_AGEMA_signal_1374), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3960), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[37]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3964), .CK(clk), .Q(new_AGEMA_signal_1371), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3968), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[36]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3972), .CK(clk), .Q(new_AGEMA_signal_1368), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3976), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[51]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3980), .CK(clk), .Q(new_AGEMA_signal_1413), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3984), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[50]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3988), .CK(clk), .Q(new_AGEMA_signal_1410), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_3992), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[49]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3996), .CK(clk), .Q(new_AGEMA_signal_1407), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_4000), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[48]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4004), .CK(clk), .Q(new_AGEMA_signal_1404), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_4008), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[43]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4012), .CK(clk), .Q(new_AGEMA_signal_1389), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_4016), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[42]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4020), .CK(clk), .Q(new_AGEMA_signal_1386), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_4024), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[41]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4028), .CK(clk), .Q(new_AGEMA_signal_1383), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_4032), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[40]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4036), .CK(clk), .Q(new_AGEMA_signal_1380), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_4040), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[59]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4044), .CK(clk), .Q(new_AGEMA_signal_1437), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_4048), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[58]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4052), .CK(clk), .Q(new_AGEMA_signal_1434), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_4056), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[57]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4060), .CK(clk), .Q(new_AGEMA_signal_1431), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_4064), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[56]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4068), .CK(clk), .Q(new_AGEMA_signal_1428), .QN()
         );
endmodule

