/* modified netlist. Source: module sbox in file Designs/AESSbox/lookup/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 34 time(s)  */

module sbox_HPC1_ClockGating_d1 (SI_s0, clk, SI_s1, Fresh, rst, SO_s0, SO_s1, Synch);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input rst ;
    input [1735:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output Synch ;
    wire N169 ;
    wire N277 ;
    wire N379 ;
    wire N470 ;
    wire N563 ;
    wire N639 ;
    wire N723 ;
    wire N789 ;
    wire n1922 ;
    wire n1923 ;
    wire n1924 ;
    wire n1925 ;
    wire n1926 ;
    wire n1927 ;
    wire n1928 ;
    wire n1929 ;
    wire n1930 ;
    wire n1931 ;
    wire n1932 ;
    wire n1933 ;
    wire n1934 ;
    wire n1935 ;
    wire n1936 ;
    wire n1937 ;
    wire n1938 ;
    wire n1939 ;
    wire n1940 ;
    wire n1941 ;
    wire n1942 ;
    wire n1943 ;
    wire n1944 ;
    wire n1945 ;
    wire n1946 ;
    wire n1947 ;
    wire n1948 ;
    wire n1949 ;
    wire n1950 ;
    wire n1951 ;
    wire n1952 ;
    wire n1953 ;
    wire n1954 ;
    wire n1955 ;
    wire n1956 ;
    wire n1957 ;
    wire n1958 ;
    wire n1959 ;
    wire n1960 ;
    wire n1961 ;
    wire n1962 ;
    wire n1963 ;
    wire n1964 ;
    wire n1965 ;
    wire n1966 ;
    wire n1967 ;
    wire n1968 ;
    wire n1969 ;
    wire n1970 ;
    wire n1971 ;
    wire n1972 ;
    wire n1973 ;
    wire n1974 ;
    wire n1975 ;
    wire n1976 ;
    wire n1977 ;
    wire n1978 ;
    wire n1979 ;
    wire n1980 ;
    wire n1981 ;
    wire n1982 ;
    wire n1983 ;
    wire n1984 ;
    wire n1985 ;
    wire n1986 ;
    wire n1987 ;
    wire n1988 ;
    wire n1989 ;
    wire n1990 ;
    wire n1991 ;
    wire n1992 ;
    wire n1993 ;
    wire n1994 ;
    wire n1995 ;
    wire n1996 ;
    wire n1997 ;
    wire n1998 ;
    wire n1999 ;
    wire n2000 ;
    wire n2001 ;
    wire n2002 ;
    wire n2003 ;
    wire n2004 ;
    wire n2005 ;
    wire n2006 ;
    wire n2007 ;
    wire n2008 ;
    wire n2009 ;
    wire n2010 ;
    wire n2011 ;
    wire n2012 ;
    wire n2013 ;
    wire n2014 ;
    wire n2015 ;
    wire n2016 ;
    wire n2017 ;
    wire n2018 ;
    wire n2019 ;
    wire n2020 ;
    wire n2021 ;
    wire n2022 ;
    wire n2023 ;
    wire n2024 ;
    wire n2025 ;
    wire n2026 ;
    wire n2027 ;
    wire n2028 ;
    wire n2029 ;
    wire n2030 ;
    wire n2031 ;
    wire n2032 ;
    wire n2033 ;
    wire n2034 ;
    wire n2035 ;
    wire n2036 ;
    wire n2037 ;
    wire n2038 ;
    wire n2039 ;
    wire n2040 ;
    wire n2041 ;
    wire n2042 ;
    wire n2043 ;
    wire n2044 ;
    wire n2045 ;
    wire n2046 ;
    wire n2047 ;
    wire n2048 ;
    wire n2049 ;
    wire n2050 ;
    wire n2051 ;
    wire n2052 ;
    wire n2053 ;
    wire n2054 ;
    wire n2055 ;
    wire n2056 ;
    wire n2057 ;
    wire n2058 ;
    wire n2059 ;
    wire n2060 ;
    wire n2061 ;
    wire n2062 ;
    wire n2063 ;
    wire n2064 ;
    wire n2065 ;
    wire n2066 ;
    wire n2067 ;
    wire n2068 ;
    wire n2069 ;
    wire n2070 ;
    wire n2071 ;
    wire n2072 ;
    wire n2073 ;
    wire n2074 ;
    wire n2075 ;
    wire n2076 ;
    wire n2077 ;
    wire n2078 ;
    wire n2079 ;
    wire n2080 ;
    wire n2081 ;
    wire n2082 ;
    wire n2083 ;
    wire n2084 ;
    wire n2085 ;
    wire n2086 ;
    wire n2087 ;
    wire n2088 ;
    wire n2089 ;
    wire n2090 ;
    wire n2091 ;
    wire n2092 ;
    wire n2093 ;
    wire n2094 ;
    wire n2095 ;
    wire n2096 ;
    wire n2097 ;
    wire n2098 ;
    wire n2099 ;
    wire n2100 ;
    wire n2101 ;
    wire n2102 ;
    wire n2103 ;
    wire n2104 ;
    wire n2105 ;
    wire n2106 ;
    wire n2107 ;
    wire n2108 ;
    wire n2109 ;
    wire n2110 ;
    wire n2111 ;
    wire n2112 ;
    wire n2113 ;
    wire n2114 ;
    wire n2115 ;
    wire n2116 ;
    wire n2117 ;
    wire n2118 ;
    wire n2119 ;
    wire n2120 ;
    wire n2121 ;
    wire n2122 ;
    wire n2123 ;
    wire n2124 ;
    wire n2125 ;
    wire n2126 ;
    wire n2127 ;
    wire n2128 ;
    wire n2129 ;
    wire n2130 ;
    wire n2131 ;
    wire n2132 ;
    wire n2133 ;
    wire n2134 ;
    wire n2135 ;
    wire n2136 ;
    wire n2137 ;
    wire n2138 ;
    wire n2139 ;
    wire n2140 ;
    wire n2141 ;
    wire n2142 ;
    wire n2143 ;
    wire n2144 ;
    wire n2145 ;
    wire n2146 ;
    wire n2147 ;
    wire n2148 ;
    wire n2149 ;
    wire n2150 ;
    wire n2151 ;
    wire n2152 ;
    wire n2153 ;
    wire n2154 ;
    wire n2155 ;
    wire n2156 ;
    wire n2157 ;
    wire n2158 ;
    wire n2159 ;
    wire n2160 ;
    wire n2161 ;
    wire n2162 ;
    wire n2163 ;
    wire n2164 ;
    wire n2165 ;
    wire n2166 ;
    wire n2167 ;
    wire n2168 ;
    wire n2169 ;
    wire n2170 ;
    wire n2171 ;
    wire n2172 ;
    wire n2173 ;
    wire n2174 ;
    wire n2175 ;
    wire n2176 ;
    wire n2177 ;
    wire n2178 ;
    wire n2179 ;
    wire n2180 ;
    wire n2181 ;
    wire n2182 ;
    wire n2183 ;
    wire n2184 ;
    wire n2185 ;
    wire n2186 ;
    wire n2187 ;
    wire n2188 ;
    wire n2189 ;
    wire n2190 ;
    wire n2191 ;
    wire n2192 ;
    wire n2193 ;
    wire n2194 ;
    wire n2195 ;
    wire n2196 ;
    wire n2197 ;
    wire n2198 ;
    wire n2199 ;
    wire n2200 ;
    wire n2201 ;
    wire n2202 ;
    wire n2203 ;
    wire n2204 ;
    wire n2205 ;
    wire n2206 ;
    wire n2207 ;
    wire n2208 ;
    wire n2209 ;
    wire n2210 ;
    wire n2211 ;
    wire n2212 ;
    wire n2213 ;
    wire n2214 ;
    wire n2215 ;
    wire n2216 ;
    wire n2217 ;
    wire n2218 ;
    wire n2219 ;
    wire n2220 ;
    wire n2221 ;
    wire n2222 ;
    wire n2223 ;
    wire n2224 ;
    wire n2225 ;
    wire n2226 ;
    wire n2227 ;
    wire n2228 ;
    wire n2229 ;
    wire n2230 ;
    wire n2231 ;
    wire n2232 ;
    wire n2233 ;
    wire n2234 ;
    wire n2235 ;
    wire n2236 ;
    wire n2237 ;
    wire n2238 ;
    wire n2239 ;
    wire n2240 ;
    wire n2241 ;
    wire n2242 ;
    wire n2243 ;
    wire n2244 ;
    wire n2245 ;
    wire n2246 ;
    wire n2247 ;
    wire n2248 ;
    wire n2249 ;
    wire n2250 ;
    wire n2251 ;
    wire n2252 ;
    wire n2253 ;
    wire n2254 ;
    wire n2255 ;
    wire n2256 ;
    wire n2257 ;
    wire n2258 ;
    wire n2259 ;
    wire n2260 ;
    wire n2261 ;
    wire n2262 ;
    wire n2263 ;
    wire n2264 ;
    wire n2265 ;
    wire n2266 ;
    wire n2267 ;
    wire n2268 ;
    wire n2269 ;
    wire n2270 ;
    wire n2271 ;
    wire n2272 ;
    wire n2273 ;
    wire n2274 ;
    wire n2275 ;
    wire n2276 ;
    wire n2277 ;
    wire n2278 ;
    wire n2279 ;
    wire n2280 ;
    wire n2281 ;
    wire n2282 ;
    wire n2283 ;
    wire n2284 ;
    wire n2285 ;
    wire n2286 ;
    wire n2287 ;
    wire n2288 ;
    wire n2289 ;
    wire n2290 ;
    wire n2291 ;
    wire n2292 ;
    wire n2293 ;
    wire n2294 ;
    wire n2295 ;
    wire n2296 ;
    wire n2297 ;
    wire n2298 ;
    wire n2299 ;
    wire n2300 ;
    wire n2301 ;
    wire n2302 ;
    wire n2303 ;
    wire n2304 ;
    wire n2305 ;
    wire n2306 ;
    wire n2307 ;
    wire n2308 ;
    wire n2309 ;
    wire n2310 ;
    wire n2311 ;
    wire n2312 ;
    wire n2313 ;
    wire n2314 ;
    wire n2315 ;
    wire n2316 ;
    wire n2317 ;
    wire n2318 ;
    wire n2319 ;
    wire n2320 ;
    wire n2321 ;
    wire n2322 ;
    wire n2323 ;
    wire n2324 ;
    wire n2325 ;
    wire n2326 ;
    wire n2327 ;
    wire n2328 ;
    wire n2329 ;
    wire n2330 ;
    wire n2331 ;
    wire n2332 ;
    wire n2333 ;
    wire n2334 ;
    wire n2335 ;
    wire n2336 ;
    wire n2337 ;
    wire n2338 ;
    wire n2339 ;
    wire n2340 ;
    wire n2341 ;
    wire n2342 ;
    wire n2343 ;
    wire n2344 ;
    wire n2345 ;
    wire n2346 ;
    wire n2347 ;
    wire n2348 ;
    wire n2349 ;
    wire n2350 ;
    wire n2351 ;
    wire n2352 ;
    wire n2353 ;
    wire n2354 ;
    wire n2355 ;
    wire n2356 ;
    wire n2357 ;
    wire n2358 ;
    wire n2359 ;
    wire n2360 ;
    wire n2361 ;
    wire n2362 ;
    wire n2363 ;
    wire n2364 ;
    wire n2365 ;
    wire n2366 ;
    wire n2367 ;
    wire n2368 ;
    wire n2369 ;
    wire n2370 ;
    wire n2371 ;
    wire n2372 ;
    wire n2373 ;
    wire n2374 ;
    wire n2375 ;
    wire n2376 ;
    wire n2377 ;
    wire n2378 ;
    wire n2379 ;
    wire n2380 ;
    wire n2381 ;
    wire n2382 ;
    wire n2383 ;
    wire n2384 ;
    wire n2385 ;
    wire n2386 ;
    wire n2387 ;
    wire n2388 ;
    wire n2389 ;
    wire n2390 ;
    wire n2391 ;
    wire n2392 ;
    wire n2393 ;
    wire n2394 ;
    wire n2395 ;
    wire n2396 ;
    wire n2397 ;
    wire n2398 ;
    wire n2399 ;
    wire n2400 ;
    wire n2401 ;
    wire n2402 ;
    wire n2403 ;
    wire n2404 ;
    wire n2405 ;
    wire n2406 ;
    wire n2407 ;
    wire n2408 ;
    wire n2409 ;
    wire n2410 ;
    wire n2411 ;
    wire n2412 ;
    wire n2413 ;
    wire n2414 ;
    wire n2415 ;
    wire n2416 ;
    wire n2417 ;
    wire n2418 ;
    wire n2419 ;
    wire n2420 ;
    wire n2421 ;
    wire n2422 ;
    wire n2423 ;
    wire n2424 ;
    wire n2425 ;
    wire n2426 ;
    wire n2427 ;
    wire n2428 ;
    wire n2429 ;
    wire n2430 ;
    wire n2431 ;
    wire n2432 ;
    wire n2433 ;
    wire n2434 ;
    wire n2435 ;
    wire n2436 ;
    wire n2437 ;
    wire n2438 ;
    wire n2439 ;
    wire n2440 ;
    wire n2441 ;
    wire n2442 ;
    wire n2443 ;
    wire n2444 ;
    wire n2445 ;
    wire n2446 ;
    wire n2447 ;
    wire n2448 ;
    wire n2449 ;
    wire n2450 ;
    wire n2451 ;
    wire n2452 ;
    wire n2453 ;
    wire n2454 ;
    wire n2455 ;
    wire n2456 ;
    wire n2457 ;
    wire n2458 ;
    wire n2459 ;
    wire n2460 ;
    wire n2461 ;
    wire n2462 ;
    wire n2463 ;
    wire n2464 ;
    wire n2465 ;
    wire n2466 ;
    wire n2467 ;
    wire n2468 ;
    wire n2469 ;
    wire n2470 ;
    wire n2471 ;
    wire n2472 ;
    wire n2473 ;
    wire n2474 ;
    wire n2475 ;
    wire n2476 ;
    wire n2477 ;
    wire n2478 ;
    wire n2479 ;
    wire n2480 ;
    wire n2481 ;
    wire n2482 ;
    wire n2483 ;
    wire n2484 ;
    wire n2485 ;
    wire n2486 ;
    wire n2487 ;
    wire n2488 ;
    wire n2489 ;
    wire n2490 ;
    wire n2491 ;
    wire n2492 ;
    wire n2493 ;
    wire n2494 ;
    wire n2495 ;
    wire n2496 ;
    wire n2497 ;
    wire n2498 ;
    wire n2499 ;
    wire n2500 ;
    wire n2501 ;
    wire n2502 ;
    wire n2503 ;
    wire n2504 ;
    wire n2505 ;
    wire n2506 ;
    wire n2507 ;
    wire n2508 ;
    wire n2509 ;
    wire n2510 ;
    wire n2511 ;
    wire n2512 ;
    wire n2513 ;
    wire n2514 ;
    wire n2515 ;
    wire n2516 ;
    wire n2517 ;
    wire n2518 ;
    wire n2519 ;
    wire n2520 ;
    wire n2521 ;
    wire n2522 ;
    wire n2523 ;
    wire n2524 ;
    wire n2525 ;
    wire n2526 ;
    wire n2527 ;
    wire n2528 ;
    wire n2529 ;
    wire n2530 ;
    wire n2531 ;
    wire n2532 ;
    wire n2533 ;
    wire n2534 ;
    wire n2535 ;
    wire n2536 ;
    wire n2537 ;
    wire n2538 ;
    wire n2539 ;
    wire n2540 ;
    wire n2541 ;
    wire n2542 ;
    wire n2543 ;
    wire n2544 ;
    wire n2545 ;
    wire n2546 ;
    wire n2547 ;
    wire n2548 ;
    wire n2549 ;
    wire n2550 ;
    wire n2551 ;
    wire n2552 ;
    wire n2553 ;
    wire n2554 ;
    wire n2555 ;
    wire n2556 ;
    wire n2557 ;
    wire n2558 ;
    wire n2559 ;
    wire n2560 ;
    wire n2561 ;
    wire n2562 ;
    wire n2563 ;
    wire n2564 ;
    wire n2565 ;
    wire n2566 ;
    wire n2567 ;
    wire n2568 ;
    wire n2569 ;
    wire n2570 ;
    wire n2571 ;
    wire n2572 ;
    wire n2573 ;
    wire n2574 ;
    wire n2575 ;
    wire n2576 ;
    wire n2577 ;
    wire n2578 ;
    wire n2579 ;
    wire n2580 ;
    wire n2581 ;
    wire n2582 ;
    wire n2583 ;
    wire n2584 ;
    wire n2585 ;
    wire n2586 ;
    wire n2587 ;
    wire n2588 ;
    wire n2589 ;
    wire n2590 ;
    wire n2591 ;
    wire n2592 ;
    wire n2593 ;
    wire n2594 ;
    wire n2595 ;
    wire n2596 ;
    wire n2597 ;
    wire n2598 ;
    wire n2599 ;
    wire n2600 ;
    wire n2601 ;
    wire n2602 ;
    wire n2603 ;
    wire n2604 ;
    wire n2605 ;
    wire n2606 ;
    wire n2607 ;
    wire n2608 ;
    wire n2609 ;
    wire n2610 ;
    wire n2611 ;
    wire n2612 ;
    wire n2613 ;
    wire n2614 ;
    wire n2615 ;
    wire n2616 ;
    wire n2617 ;
    wire n2618 ;
    wire n2619 ;
    wire n2620 ;
    wire n2621 ;
    wire n2622 ;
    wire n2623 ;
    wire n2624 ;
    wire n2625 ;
    wire n2626 ;
    wire n2627 ;
    wire n2628 ;
    wire n2629 ;
    wire n2630 ;
    wire n2631 ;
    wire n2632 ;
    wire n2633 ;
    wire n2634 ;
    wire n2635 ;
    wire n2636 ;
    wire n2637 ;
    wire n2638 ;
    wire n2639 ;
    wire n2640 ;
    wire n2641 ;
    wire n2642 ;
    wire n2643 ;
    wire n2644 ;
    wire n2645 ;
    wire n2646 ;
    wire n2647 ;
    wire n2648 ;
    wire n2649 ;
    wire n2650 ;
    wire n2651 ;
    wire n2652 ;
    wire n2653 ;
    wire n2654 ;
    wire n2655 ;
    wire n2656 ;
    wire n2657 ;
    wire n2658 ;
    wire n2659 ;
    wire n2660 ;
    wire n2661 ;
    wire n2662 ;
    wire n2663 ;
    wire n2664 ;
    wire n2665 ;
    wire n2666 ;
    wire n2667 ;
    wire n2668 ;
    wire n2669 ;
    wire n2670 ;
    wire n2671 ;
    wire n2672 ;
    wire n2673 ;
    wire n2674 ;
    wire n2675 ;
    wire n2676 ;
    wire n2677 ;
    wire n2678 ;
    wire n2679 ;
    wire n2680 ;
    wire n2681 ;
    wire n2682 ;
    wire n2683 ;
    wire n2684 ;
    wire n2685 ;
    wire n2686 ;
    wire n2687 ;
    wire n2688 ;
    wire n2689 ;
    wire n2690 ;
    wire n2691 ;
    wire n2692 ;
    wire n2693 ;
    wire n2694 ;
    wire n2695 ;
    wire n2696 ;
    wire n2697 ;
    wire n2698 ;
    wire n2699 ;
    wire n2700 ;
    wire n2701 ;
    wire n2702 ;
    wire n2703 ;
    wire n2704 ;
    wire n2705 ;
    wire n2706 ;
    wire n2707 ;
    wire n2708 ;
    wire n2709 ;
    wire n2710 ;
    wire n2711 ;
    wire n2712 ;
    wire n2713 ;
    wire n2714 ;
    wire n2715 ;
    wire n2716 ;
    wire n2717 ;
    wire n2718 ;
    wire n2719 ;
    wire n2720 ;
    wire n2721 ;
    wire n2722 ;
    wire n2723 ;
    wire n2724 ;
    wire n2725 ;
    wire n2726 ;
    wire n2727 ;
    wire n2728 ;
    wire n2729 ;
    wire n2730 ;
    wire n2731 ;
    wire n2732 ;
    wire n2733 ;
    wire n2734 ;
    wire n2735 ;
    wire n2736 ;
    wire n2737 ;
    wire n2738 ;
    wire n2739 ;
    wire n2740 ;
    wire n2741 ;
    wire n2742 ;
    wire n2743 ;
    wire n2744 ;
    wire n2745 ;
    wire n2746 ;
    wire n2747 ;
    wire n2748 ;
    wire n2749 ;
    wire n2750 ;
    wire n2751 ;
    wire n2752 ;
    wire n2753 ;
    wire n2754 ;
    wire n2755 ;
    wire n2756 ;
    wire n2757 ;
    wire n2758 ;
    wire n2759 ;
    wire n2760 ;
    wire n2761 ;
    wire n2762 ;
    wire n2763 ;
    wire n2764 ;
    wire n2765 ;
    wire n2766 ;
    wire n2767 ;
    wire n2768 ;
    wire n2769 ;
    wire n2770 ;
    wire n2771 ;
    wire n2772 ;
    wire n2773 ;
    wire n2774 ;
    wire n2775 ;
    wire n2776 ;
    wire n2777 ;
    wire n2778 ;
    wire n2779 ;
    wire n2780 ;
    wire n2781 ;
    wire n2782 ;
    wire n2783 ;
    wire n2784 ;
    wire n2785 ;
    wire n2786 ;
    wire n2787 ;
    wire n2788 ;
    wire n2789 ;
    wire n2790 ;
    wire n2791 ;
    wire n2792 ;
    wire n2793 ;
    wire n2794 ;
    wire n2795 ;
    wire n2796 ;
    wire n2797 ;
    wire n2798 ;
    wire n2799 ;
    wire n2800 ;
    wire n2801 ;
    wire n2802 ;
    wire n2803 ;
    wire n2804 ;
    wire n2805 ;
    wire n2806 ;
    wire n2807 ;
    wire n2808 ;
    wire n2809 ;
    wire n2810 ;
    wire n2811 ;
    wire n2812 ;
    wire n2813 ;
    wire n2814 ;
    wire n2815 ;
    wire n2816 ;
    wire n2817 ;
    wire n2818 ;
    wire n2819 ;
    wire n2820 ;
    wire n2821 ;
    wire n2822 ;
    wire n2823 ;
    wire n2824 ;
    wire n2825 ;
    wire n2826 ;
    wire n2827 ;
    wire n2828 ;
    wire n2829 ;
    wire n2830 ;
    wire n2831 ;
    wire n2832 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire clk_gated ;

    /* cells in depth 0 */
    not_masked #(.security_order(1), .pipeline(0)) U1938 ( .a ({SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_943, n2796}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1939 ( .a ({SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_945, n2810}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1940 ( .a ({SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_947, n2462}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1941 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_949, n2760}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1942 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_951, n2791}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1944 ( .a ({SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_953, n2813}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1945 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_955, n2630}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1946 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_957, n2765}) ) ;
    ClockGatingController #(35) ClockGatingInst ( .clk ( clk ), .rst ( rst ), .GatedClk ( clk_gated ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1937 ( .ina ({new_AGEMA_signal_943, n2796}), .inb ({SI_s1[6], SI_s0[6]}), .clk ( clk ), .rnd ({Fresh[1], Fresh[0]}), .outt ({new_AGEMA_signal_970, n2719}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1943 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_1023, n2672}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1947 ( .ina ({SI_s1[2], SI_s0[2]}), .inb ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[3], Fresh[2]}), .outt ({new_AGEMA_signal_958, n2635}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1948 ( .ina ({new_AGEMA_signal_947, n2462}), .inb ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[5], Fresh[4]}), .outt ({new_AGEMA_signal_971, n2641}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1949 ( .ina ({SI_s1[6], SI_s0[6]}), .inb ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[7], Fresh[6]}), .outt ({new_AGEMA_signal_959, n2790}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1950 ( .ina ({SI_s1[6], SI_s0[6]}), .inb ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[9], Fresh[8]}), .outt ({new_AGEMA_signal_960, n2519}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1951 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_972, n2750}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1952 ( .ina ({new_AGEMA_signal_949, n2760}), .inb ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[11], Fresh[10]}), .outt ({new_AGEMA_signal_973, n2615}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1953 ( .a ({new_AGEMA_signal_973, n2615}), .b ({new_AGEMA_signal_1024, n2640}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1955 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[13], Fresh[12]}), .outt ({new_AGEMA_signal_974, n2699}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1956 ( .a ({new_AGEMA_signal_974, n2699}), .b ({new_AGEMA_signal_1025, n2737}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1957 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .rnd ({Fresh[15], Fresh[14]}), .outt ({new_AGEMA_signal_975, n2816}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1958 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_1026, n2767}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1961 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[17], Fresh[16]}), .outt ({new_AGEMA_signal_976, n2780}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1962 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_1027, n2789}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1963 ( .ina ({SI_s1[6], SI_s0[6]}), .inb ({new_AGEMA_signal_945, n2810}), .clk ( clk ), .rnd ({Fresh[19], Fresh[18]}), .outt ({new_AGEMA_signal_977, n2317}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1965 ( .ina ({new_AGEMA_signal_951, n2791}), .inb ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .rnd ({Fresh[21], Fresh[20]}), .outt ({new_AGEMA_signal_978, n2694}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1966 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_1028, n2769}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1969 ( .ina ({new_AGEMA_signal_949, n2760}), .inb ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[23], Fresh[22]}), .outt ({new_AGEMA_signal_979, n2073}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1970 ( .a ({new_AGEMA_signal_979, n2073}), .b ({new_AGEMA_signal_1029, n2707}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1971 ( .ina ({SI_s1[7], SI_s0[7]}), .inb ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[25], Fresh[24]}), .outt ({new_AGEMA_signal_961, n2315}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1972 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[27], Fresh[26]}), .outt ({new_AGEMA_signal_962, n2682}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1973 ( .a ({new_AGEMA_signal_962, n2682}), .b ({new_AGEMA_signal_980, n2713}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1975 ( .ina ({new_AGEMA_signal_953, n2813}), .inb ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[29], Fresh[28]}), .outt ({new_AGEMA_signal_981, n2723}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1976 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1031, n2688}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1978 ( .ina ({new_AGEMA_signal_945, n2810}), .inb ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[31], Fresh[30]}), .outt ({new_AGEMA_signal_982, n2725}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1979 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1032, n2541}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1984 ( .ina ({new_AGEMA_signal_949, n2760}), .inb ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[33], Fresh[32]}), .outt ({new_AGEMA_signal_983, n2815}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1985 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_1033, n2086}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1987 ( .ina ({new_AGEMA_signal_945, n2810}), .inb ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .rnd ({Fresh[35], Fresh[34]}), .outt ({new_AGEMA_signal_984, n2600}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1990 ( .ina ({new_AGEMA_signal_947, n2462}), .inb ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[37], Fresh[36]}), .outt ({new_AGEMA_signal_985, n2538}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1991 ( .a ({new_AGEMA_signal_985, n2538}), .b ({new_AGEMA_signal_1035, n2786}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1995 ( .ina ({SI_s1[4], SI_s0[4]}), .inb ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[39], Fresh[38]}), .outt ({new_AGEMA_signal_963, n2595}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1996 ( .a ({new_AGEMA_signal_963, n2595}), .b ({new_AGEMA_signal_986, n2742}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1999 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[41], Fresh[40]}), .outt ({new_AGEMA_signal_987, n2753}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2000 ( .a ({new_AGEMA_signal_987, n2753}), .b ({new_AGEMA_signal_1037, n2577}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2004 ( .ina ({new_AGEMA_signal_945, n2810}), .inb ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[43], Fresh[42]}), .outt ({new_AGEMA_signal_988, n2400}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2008 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[45], Fresh[44]}), .outt ({new_AGEMA_signal_989, n2785}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2009 ( .a ({new_AGEMA_signal_989, n2785}), .b ({new_AGEMA_signal_1039, n2792}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2013 ( .ina ({new_AGEMA_signal_953, n2813}), .inb ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[47], Fresh[46]}), .outt ({new_AGEMA_signal_990, n2609}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2014 ( .a ({new_AGEMA_signal_990, n2609}), .b ({new_AGEMA_signal_1040, n2724}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2017 ( .ina ({new_AGEMA_signal_949, n2760}), .inb ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .rnd ({Fresh[49], Fresh[48]}), .outt ({new_AGEMA_signal_991, n2661}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2018 ( .a ({new_AGEMA_signal_991, n2661}), .b ({new_AGEMA_signal_1041, n2174}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2020 ( .ina ({SI_s1[2], SI_s0[2]}), .inb ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[51], Fresh[50]}), .outt ({new_AGEMA_signal_964, n2708}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2021 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_992, n2493}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2025 ( .ina ({new_AGEMA_signal_943, n2796}), .inb ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[53], Fresh[52]}), .outt ({new_AGEMA_signal_993, n2587}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2028 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_1044, n2570}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2029 ( .ina ({SI_s1[5], SI_s0[5]}), .inb ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[55], Fresh[54]}), .outt ({new_AGEMA_signal_965, n2559}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2035 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[57], Fresh[56]}), .outt ({new_AGEMA_signal_994, n2643}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2036 ( .a ({new_AGEMA_signal_994, n2643}), .b ({new_AGEMA_signal_1045, n2442}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2038 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_995, n2739}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2044 ( .ina ({new_AGEMA_signal_947, n2462}), .inb ({new_AGEMA_signal_943, n2796}), .clk ( clk ), .rnd ({Fresh[59], Fresh[58]}), .outt ({new_AGEMA_signal_996, n2437}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2045 ( .ina ({SI_s1[5], SI_s0[5]}), .inb ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[61], Fresh[60]}), .outt ({new_AGEMA_signal_966, n2261}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2046 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_997, n2778}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2052 ( .ina ({SI_s1[7], SI_s0[7]}), .inb ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .rnd ({Fresh[63], Fresh[62]}), .outt ({new_AGEMA_signal_998, n2452}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2055 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_1050, n2766}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2068 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[65], Fresh[64]}), .outt ({new_AGEMA_signal_1000, n2772}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2070 ( .ina ({new_AGEMA_signal_951, n2791}), .inb ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[67], Fresh[66]}), .outt ({new_AGEMA_signal_1001, n2824}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2071 ( .a ({new_AGEMA_signal_1001, n2824}), .b ({new_AGEMA_signal_1053, n2612}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2074 ( .a ({new_AGEMA_signal_988, n2400}), .b ({new_AGEMA_signal_1054, n2313}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2089 ( .ina ({new_AGEMA_signal_945, n2810}), .inb ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .rnd ({Fresh[69], Fresh[68]}), .outt ({new_AGEMA_signal_1002, n2395}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2090 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_1058, n2818}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2094 ( .ina ({SI_s1[6], SI_s0[6]}), .inb ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[71], Fresh[70]}), .outt ({new_AGEMA_signal_967, n2779}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2096 ( .ina ({new_AGEMA_signal_955, n2630}), .inb ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .rnd ({Fresh[73], Fresh[72]}), .outt ({new_AGEMA_signal_1003, n2624}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2097 ( .ina ({SI_s1[4], SI_s0[4]}), .inb ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[75], Fresh[74]}), .outt ({new_AGEMA_signal_968, n2242}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2100 ( .ina ({SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .rnd ({Fresh[77], Fresh[76]}), .outt ({new_AGEMA_signal_1004, n2356}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2119 ( .a ({new_AGEMA_signal_1000, n2772}), .b ({new_AGEMA_signal_1063, n2823}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2122 ( .ina ({new_AGEMA_signal_949, n2760}), .inb ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[79], Fresh[78]}), .outt ({new_AGEMA_signal_1005, n2611}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2131 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_1065, n2828}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2133 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[81], Fresh[80]}), .outt ({new_AGEMA_signal_1006, n2616}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2134 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1066, n2679}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2138 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .rnd ({Fresh[83], Fresh[82]}), .outt ({new_AGEMA_signal_1007, n2563}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2139 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1067, n2809}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2150 ( .a ({new_AGEMA_signal_1005, n2611}), .b ({new_AGEMA_signal_1068, n2709}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2163 ( .ina ({new_AGEMA_signal_943, n2796}), .inb ({new_AGEMA_signal_945, n2810}), .clk ( clk ), .rnd ({Fresh[85], Fresh[84]}), .outt ({new_AGEMA_signal_1008, n2401}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2211 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[87], Fresh[86]}), .outt ({new_AGEMA_signal_1010, n2061}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2232 ( .ina ({new_AGEMA_signal_943, n2796}), .inb ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .rnd ({Fresh[89], Fresh[88]}), .outt ({new_AGEMA_signal_1011, n2721}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2276 ( .ina ({new_AGEMA_signal_951, n2791}), .inb ({new_AGEMA_signal_957, n2765}), .clk ( clk ), .rnd ({Fresh[91], Fresh[90]}), .outt ({new_AGEMA_signal_1012, n2298}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2278 ( .a ({new_AGEMA_signal_1008, n2401}), .b ({new_AGEMA_signal_1080, n2118}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2307 ( .ina ({SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[93], Fresh[92]}), .outt ({new_AGEMA_signal_1013, n2346}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2341 ( .ina ({SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .rnd ({Fresh[95], Fresh[94]}), .outt ({new_AGEMA_signal_1015, n2430}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2383 ( .ina ({SI_s1[5], SI_s0[5]}), .inb ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[97], Fresh[96]}), .outt ({new_AGEMA_signal_969, n2712}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2402 ( .ina ({SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .rnd ({Fresh[99], Fresh[98]}), .outt ({new_AGEMA_signal_1017, n2777}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2615 ( .ina ({SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_947, n2462}), .clk ( clk ), .rnd ({Fresh[101], Fresh[100]}), .outt ({new_AGEMA_signal_1019, n2463}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2627 ( .ina ({new_AGEMA_signal_945, n2810}), .inb ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[103], Fresh[102]}), .outt ({new_AGEMA_signal_1020, n2474}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1954 ( .ina ({new_AGEMA_signal_972, n2750}), .inb ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .rnd ({Fresh[105], Fresh[104]}), .outt ({new_AGEMA_signal_1127, n2575}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1959 ( .ina ({new_AGEMA_signal_1025, n2737}), .inb ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .rnd ({Fresh[107], Fresh[106]}), .outt ({new_AGEMA_signal_1128, n1962}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1964 ( .ina ({new_AGEMA_signal_1027, n2789}), .inb ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .rnd ({Fresh[109], Fresh[108]}), .outt ({new_AGEMA_signal_1129, n1922}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1974 ( .ina ({new_AGEMA_signal_961, n2315}), .inb ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .rnd ({Fresh[111], Fresh[110]}), .outt ({new_AGEMA_signal_1030, n2755}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1977 ( .ina ({new_AGEMA_signal_977, n2317}), .inb ({new_AGEMA_signal_1031, n2688}), .clk ( clk ), .rnd ({Fresh[113], Fresh[112]}), .outt ({new_AGEMA_signal_1130, n1926}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1980 ( .ina ({new_AGEMA_signal_1026, n2767}), .inb ({new_AGEMA_signal_1032, n2541}), .clk ( clk ), .rnd ({Fresh[115], Fresh[114]}), .outt ({new_AGEMA_signal_1131, n1925}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1986 ( .ina ({new_AGEMA_signal_1033, n2086}), .inb ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .rnd ({Fresh[117], Fresh[116]}), .outt ({new_AGEMA_signal_1132, n2151}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1988 ( .ina ({new_AGEMA_signal_971, n2641}), .inb ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .rnd ({Fresh[119], Fresh[118]}), .outt ({new_AGEMA_signal_1034, n2631}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U1989 ( .a ({new_AGEMA_signal_1034, n2631}), .b ({new_AGEMA_signal_1133, n2734}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1992 ( .ina ({new_AGEMA_signal_1029, n2707}), .inb ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .rnd ({Fresh[121], Fresh[120]}), .outt ({new_AGEMA_signal_1134, n2763}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1997 ( .ina ({new_AGEMA_signal_960, n2519}), .inb ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .rnd ({Fresh[123], Fresh[122]}), .outt ({new_AGEMA_signal_1036, n1930}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2005 ( .ina ({new_AGEMA_signal_988, n2400}), .inb ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .rnd ({Fresh[125], Fresh[124]}), .outt ({new_AGEMA_signal_1038, n2492}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2006 ( .a ({new_AGEMA_signal_1038, n2492}), .b ({new_AGEMA_signal_1135, n2732}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2010 ( .ina ({SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .rnd ({Fresh[127], Fresh[126]}), .outt ({new_AGEMA_signal_1136, n1937}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2022 ( .ina ({SI_s1[6], SI_s0[6]}), .inb ({new_AGEMA_signal_992, n2493}), .clk ( clk ), .rnd ({Fresh[129], Fresh[128]}), .outt ({new_AGEMA_signal_1042, n1942}) ) ;
    or_HPC1 #(.security_order(1), .pipeline(0)) U2026 ( .ina ({new_AGEMA_signal_993, n2587}), .inb ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .rnd ({Fresh[131], Fresh[130]}), .outt ({new_AGEMA_signal_1043, n2676}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2030 ( .ina ({new_AGEMA_signal_1027, n2789}), .inb ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .rnd ({Fresh[133], Fresh[132]}), .outt ({new_AGEMA_signal_1139, n1944}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2037 ( .ina ({new_AGEMA_signal_982, n2725}), .inb ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .rnd ({Fresh[135], Fresh[134]}), .outt ({new_AGEMA_signal_1140, n1950}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2039 ( .ina ({SI_s1[7], SI_s0[7]}), .inb ({new_AGEMA_signal_995, n2739}), .clk ( clk ), .rnd ({Fresh[137], Fresh[136]}), .outt ({new_AGEMA_signal_1046, n1949}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2042 ( .ina ({new_AGEMA_signal_972, n2750}), .inb ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .rnd ({Fresh[139], Fresh[138]}), .outt ({new_AGEMA_signal_1047, n2677}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2043 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_1141, n2662}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2047 ( .ina ({new_AGEMA_signal_996, n2437}), .inb ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .rnd ({Fresh[141], Fresh[140]}), .outt ({new_AGEMA_signal_1048, n2627}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2053 ( .ina ({new_AGEMA_signal_975, n2816}), .inb ({new_AGEMA_signal_998, n2452}), .clk ( clk ), .rnd ({Fresh[143], Fresh[142]}), .outt ({new_AGEMA_signal_1049, n1957}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2056 ( .ina ({new_AGEMA_signal_1050, n2766}), .inb ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .rnd ({Fresh[145], Fresh[144]}), .outt ({new_AGEMA_signal_1142, n2088}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2062 ( .ina ({new_AGEMA_signal_960, n2519}), .inb ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .rnd ({Fresh[147], Fresh[146]}), .outt ({new_AGEMA_signal_999, n1964}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2063 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .rnd ({Fresh[149], Fresh[148]}), .outt ({new_AGEMA_signal_1051, n2736}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2069 ( .ina ({new_AGEMA_signal_1000, n2772}), .inb ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[151], Fresh[150]}), .outt ({new_AGEMA_signal_1052, n2673}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2072 ( .ina ({new_AGEMA_signal_1050, n2766}), .inb ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .rnd ({Fresh[153], Fresh[152]}), .outt ({new_AGEMA_signal_1144, n2761}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2073 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1323, n2720}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2075 ( .ina ({new_AGEMA_signal_1054, n2313}), .inb ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .rnd ({Fresh[155], Fresh[154]}), .outt ({new_AGEMA_signal_1145, n2412}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2076 ( .a ({new_AGEMA_signal_1145, n2412}), .b ({new_AGEMA_signal_1324, n2417}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2079 ( .ina ({new_AGEMA_signal_971, n2641}), .inb ({new_AGEMA_signal_966, n2261}), .clk ( clk ), .rnd ({Fresh[157], Fresh[156]}), .outt ({new_AGEMA_signal_1055, n2571}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2080 ( .a ({new_AGEMA_signal_1055, n2571}), .b ({new_AGEMA_signal_1146, n2505}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2081 ( .ina ({new_AGEMA_signal_960, n2519}), .inb ({new_AGEMA_signal_1001, n2824}), .clk ( clk ), .rnd ({Fresh[159], Fresh[158]}), .outt ({new_AGEMA_signal_1056, n2651}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2083 ( .ina ({new_AGEMA_signal_1039, n2792}), .inb ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[161], Fresh[160]}), .outt ({new_AGEMA_signal_1147, n2359}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2086 ( .ina ({new_AGEMA_signal_960, n2519}), .inb ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .rnd ({Fresh[163], Fresh[162]}), .outt ({new_AGEMA_signal_1057, n2101}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2087 ( .a ({new_AGEMA_signal_1057, n2101}), .b ({new_AGEMA_signal_1148, n2625}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2091 ( .ina ({new_AGEMA_signal_970, n2719}), .inb ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .rnd ({Fresh[165], Fresh[164]}), .outt ({new_AGEMA_signal_1059, n2190}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2095 ( .ina ({new_AGEMA_signal_995, n2739}), .inb ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .rnd ({Fresh[167], Fresh[166]}), .outt ({new_AGEMA_signal_1060, n1976}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2098 ( .ina ({new_AGEMA_signal_1023, n2672}), .inb ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .rnd ({Fresh[169], Fresh[168]}), .outt ({new_AGEMA_signal_1150, n2535}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2101 ( .ina ({new_AGEMA_signal_1031, n2688}), .inb ({new_AGEMA_signal_1004, n2356}), .clk ( clk ), .rnd ({Fresh[171], Fresh[170]}), .outt ({new_AGEMA_signal_1151, n1973}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2105 ( .ina ({new_AGEMA_signal_983, n2815}), .inb ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .rnd ({Fresh[173], Fresh[172]}), .outt ({new_AGEMA_signal_1061, n2690}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2111 ( .ina ({new_AGEMA_signal_992, n2493}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[175], Fresh[174]}), .outt ({new_AGEMA_signal_1062, n2817}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2113 ( .ina ({new_AGEMA_signal_1045, n2442}), .inb ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .rnd ({Fresh[177], Fresh[176]}), .outt ({new_AGEMA_signal_1153, n2741}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2118 ( .ina ({new_AGEMA_signal_976, n2780}), .inb ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .rnd ({Fresh[179], Fresh[178]}), .outt ({new_AGEMA_signal_1154, n1992}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2120 ( .ina ({new_AGEMA_signal_1063, n2823}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[181], Fresh[180]}), .outt ({new_AGEMA_signal_1155, n1991}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2123 ( .ina ({new_AGEMA_signal_994, n2643}), .inb ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .rnd ({Fresh[183], Fresh[182]}), .outt ({new_AGEMA_signal_1064, n1993}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2125 ( .ina ({new_AGEMA_signal_1025, n2737}), .inb ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .rnd ({Fresh[185], Fresh[184]}), .outt ({new_AGEMA_signal_1156, n1995}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2132 ( .ina ({new_AGEMA_signal_1058, n2818}), .inb ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .rnd ({Fresh[187], Fresh[186]}), .outt ({new_AGEMA_signal_1157, n2241}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2135 ( .ina ({SI_s1[5], SI_s0[5]}), .inb ({new_AGEMA_signal_1066, n2679}), .clk ( clk ), .rnd ({Fresh[189], Fresh[188]}), .outt ({new_AGEMA_signal_1158, n2003}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2140 ( .ina ({new_AGEMA_signal_1053, n2612}), .inb ({new_AGEMA_signal_1067, n2809}), .clk ( clk ), .rnd ({Fresh[191], Fresh[190]}), .outt ({new_AGEMA_signal_1159, n2008}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2141 ( .ina ({new_AGEMA_signal_1066, n2679}), .inb ({new_AGEMA_signal_1031, n2688}), .clk ( clk ), .rnd ({Fresh[193], Fresh[192]}), .outt ({new_AGEMA_signal_1160, n2572}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2143 ( .ina ({new_AGEMA_signal_1067, n2809}), .inb ({new_AGEMA_signal_1004, n2356}), .clk ( clk ), .rnd ({Fresh[195], Fresh[194]}), .outt ({new_AGEMA_signal_1161, n2004}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2147 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[197], Fresh[196]}), .outt ({new_AGEMA_signal_1162, n2009}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2151 ( .ina ({new_AGEMA_signal_1027, n2789}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[199], Fresh[198]}), .outt ({new_AGEMA_signal_1163, n2533}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2157 ( .ina ({new_AGEMA_signal_970, n2719}), .inb ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .rnd ({Fresh[201], Fresh[200]}), .outt ({new_AGEMA_signal_1069, n2026}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2158 ( .ina ({new_AGEMA_signal_1050, n2766}), .inb ({new_AGEMA_signal_992, n2493}), .clk ( clk ), .rnd ({Fresh[203], Fresh[202]}), .outt ({new_AGEMA_signal_1164, n2022}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2159 ( .ina ({new_AGEMA_signal_947, n2462}), .inb ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .rnd ({Fresh[205], Fresh[204]}), .outt ({new_AGEMA_signal_1070, n2227}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2167 ( .ina ({new_AGEMA_signal_959, n2790}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[207], Fresh[206]}), .outt ({new_AGEMA_signal_1009, n2027}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2171 ( .ina ({new_AGEMA_signal_1058, n2818}), .inb ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .rnd ({Fresh[209], Fresh[208]}), .outt ({new_AGEMA_signal_1167, n2214}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2173 ( .ina ({new_AGEMA_signal_1045, n2442}), .inb ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .rnd ({Fresh[211], Fresh[210]}), .outt ({new_AGEMA_signal_1168, n2290}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2174 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .rnd ({Fresh[213], Fresh[212]}), .outt ({new_AGEMA_signal_1169, n2376}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2178 ( .ina ({new_AGEMA_signal_964, n2708}), .inb ({new_AGEMA_signal_988, n2400}), .clk ( clk ), .rnd ({Fresh[215], Fresh[214]}), .outt ({new_AGEMA_signal_1072, n2034}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2182 ( .ina ({new_AGEMA_signal_1005, n2611}), .inb ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .rnd ({Fresh[217], Fresh[216]}), .outt ({new_AGEMA_signal_1073, n2171}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2183 ( .ina ({new_AGEMA_signal_1065, n2828}), .inb ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .rnd ({Fresh[219], Fresh[218]}), .outt ({new_AGEMA_signal_1170, n2039}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2188 ( .ina ({new_AGEMA_signal_982, n2725}), .inb ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .rnd ({Fresh[221], Fresh[220]}), .outt ({new_AGEMA_signal_1172, n2042}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2191 ( .ina ({new_AGEMA_signal_1029, n2707}), .inb ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .rnd ({Fresh[223], Fresh[222]}), .outt ({new_AGEMA_signal_1173, n2754}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2192 ( .ina ({new_AGEMA_signal_1054, n2313}), .inb ({new_AGEMA_signal_959, n2790}), .clk ( clk ), .rnd ({Fresh[225], Fresh[224]}), .outt ({new_AGEMA_signal_1174, n2044}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2198 ( .ina ({new_AGEMA_signal_1054, n2313}), .inb ({new_AGEMA_signal_971, n2641}), .clk ( clk ), .rnd ({Fresh[227], Fresh[226]}), .outt ({new_AGEMA_signal_1175, n2654}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2202 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1037, n2577}), .clk ( clk ), .rnd ({Fresh[229], Fresh[228]}), .outt ({new_AGEMA_signal_1176, n2055}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2205 ( .ina ({new_AGEMA_signal_1002, n2395}), .inb ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .rnd ({Fresh[231], Fresh[230]}), .outt ({new_AGEMA_signal_1177, n2057}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2208 ( .ina ({new_AGEMA_signal_1066, n2679}), .inb ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .rnd ({Fresh[233], Fresh[232]}), .outt ({new_AGEMA_signal_1178, n2407}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2212 ( .ina ({new_AGEMA_signal_1031, n2688}), .inb ({new_AGEMA_signal_1010, n2061}), .clk ( clk ), .rnd ({Fresh[235], Fresh[234]}), .outt ({new_AGEMA_signal_1179, n2062}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2216 ( .ina ({new_AGEMA_signal_1050, n2766}), .inb ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .rnd ({Fresh[237], Fresh[236]}), .outt ({new_AGEMA_signal_1180, n2731}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2220 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_1181, n2068}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2224 ( .ina ({new_AGEMA_signal_1005, n2611}), .inb ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .rnd ({Fresh[239], Fresh[238]}), .outt ({new_AGEMA_signal_1074, n2642}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2225 ( .ina ({new_AGEMA_signal_982, n2725}), .inb ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .rnd ({Fresh[241], Fresh[240]}), .outt ({new_AGEMA_signal_1182, n2252}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2228 ( .ina ({new_AGEMA_signal_995, n2739}), .inb ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .rnd ({Fresh[243], Fresh[242]}), .outt ({new_AGEMA_signal_1075, n2075}) ) ;
    or_HPC1 #(.security_order(1), .pipeline(0)) U2233 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_981, n2723}), .clk ( clk ), .rnd ({Fresh[245], Fresh[244]}), .outt ({new_AGEMA_signal_1076, n2081}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2234 ( .ina ({new_AGEMA_signal_1039, n2792}), .inb ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .rnd ({Fresh[247], Fresh[246]}), .outt ({new_AGEMA_signal_1183, n2080}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2237 ( .ina ({new_AGEMA_signal_984, n2600}), .inb ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .rnd ({Fresh[249], Fresh[248]}), .outt ({new_AGEMA_signal_1077, n2498}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2238 ( .a ({new_AGEMA_signal_1077, n2498}), .b ({new_AGEMA_signal_1184, n2773}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2239 ( .ina ({new_AGEMA_signal_1026, n2767}), .inb ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .rnd ({Fresh[251], Fresh[250]}), .outt ({new_AGEMA_signal_1185, n2083}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2244 ( .ina ({SI_s1[5], SI_s0[5]}), .inb ({new_AGEMA_signal_1033, n2086}), .clk ( clk ), .rnd ({Fresh[253], Fresh[252]}), .outt ({new_AGEMA_signal_1186, n2562}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2247 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_991, n2661}), .clk ( clk ), .rnd ({Fresh[255], Fresh[254]}), .outt ({new_AGEMA_signal_1078, n2087}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2251 ( .ina ({new_AGEMA_signal_1007, n2563}), .inb ({new_AGEMA_signal_1041, n2174}), .clk ( clk ), .rnd ({Fresh[257], Fresh[256]}), .outt ({new_AGEMA_signal_1187, n2156}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2260 ( .ina ({new_AGEMA_signal_1028, n2769}), .inb ({new_AGEMA_signal_1008, n2401}), .clk ( clk ), .rnd ({Fresh[259], Fresh[258]}), .outt ({new_AGEMA_signal_1188, n2100}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2277 ( .ina ({new_AGEMA_signal_995, n2739}), .inb ({new_AGEMA_signal_1012, n2298}), .clk ( clk ), .rnd ({Fresh[261], Fresh[260]}), .outt ({new_AGEMA_signal_1079, n2544}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2279 ( .ina ({new_AGEMA_signal_1004, n2356}), .inb ({new_AGEMA_signal_1080, n2118}), .clk ( clk ), .rnd ({Fresh[263], Fresh[262]}), .outt ({new_AGEMA_signal_1191, n2121}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2284 ( .ina ({new_AGEMA_signal_1029, n2707}), .inb ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .rnd ({Fresh[265], Fresh[264]}), .outt ({new_AGEMA_signal_1193, n2122}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2286 ( .ina ({new_AGEMA_signal_1039, n2792}), .inb ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .rnd ({Fresh[267], Fresh[266]}), .outt ({new_AGEMA_signal_1194, n2811}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2294 ( .ina ({new_AGEMA_signal_996, n2437}), .inb ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .rnd ({Fresh[269], Fresh[268]}), .outt ({new_AGEMA_signal_1081, n2647}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2297 ( .ina ({new_AGEMA_signal_986, n2742}), .inb ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .rnd ({Fresh[271], Fresh[270]}), .outt ({new_AGEMA_signal_1082, n2132}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2304 ( .ina ({new_AGEMA_signal_1006, n2616}), .inb ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .rnd ({Fresh[273], Fresh[272]}), .outt ({new_AGEMA_signal_1199, n2220}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2305 ( .ina ({SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .rnd ({Fresh[275], Fresh[274]}), .outt ({new_AGEMA_signal_1200, n2138}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2312 ( .ina ({new_AGEMA_signal_1053, n2612}), .inb ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .rnd ({Fresh[277], Fresh[276]}), .outt ({new_AGEMA_signal_1201, n2555}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2322 ( .ina ({new_AGEMA_signal_1053, n2612}), .inb ({new_AGEMA_signal_943, n2796}), .clk ( clk ), .rnd ({Fresh[279], Fresh[278]}), .outt ({new_AGEMA_signal_1202, n2429}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2328 ( .ina ({new_AGEMA_signal_996, n2437}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[281], Fresh[280]}), .outt ({new_AGEMA_signal_1083, n2162}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2337 ( .ina ({new_AGEMA_signal_961, n2315}), .inb ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .rnd ({Fresh[283], Fresh[282]}), .outt ({new_AGEMA_signal_1014, n2545}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2340 ( .ina ({new_AGEMA_signal_965, n2559}), .inb ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .rnd ({Fresh[285], Fresh[284]}), .outt ({new_AGEMA_signal_1085, n2178}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2342 ( .ina ({new_AGEMA_signal_1015, n2430}), .inb ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .rnd ({Fresh[287], Fresh[286]}), .outt ({new_AGEMA_signal_1204, n2176}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2343 ( .ina ({new_AGEMA_signal_1041, n2174}), .inb ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[289], Fresh[288]}), .outt ({new_AGEMA_signal_1205, n2175}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2348 ( .ina ({new_AGEMA_signal_966, n2261}), .inb ({new_AGEMA_signal_943, n2796}), .clk ( clk ), .rnd ({Fresh[291], Fresh[290]}), .outt ({new_AGEMA_signal_1016, n2182}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2353 ( .ina ({new_AGEMA_signal_1035, n2786}), .inb ({new_AGEMA_signal_1015, n2430}), .clk ( clk ), .rnd ({Fresh[293], Fresh[292]}), .outt ({new_AGEMA_signal_1206, n2188}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2355 ( .ina ({new_AGEMA_signal_1039, n2792}), .inb ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .rnd ({Fresh[295], Fresh[294]}), .outt ({new_AGEMA_signal_1207, n2189}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2357 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .rnd ({Fresh[297], Fresh[296]}), .outt ({new_AGEMA_signal_1208, n2446}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2362 ( .ina ({new_AGEMA_signal_972, n2750}), .inb ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .rnd ({Fresh[299], Fresh[298]}), .outt ({new_AGEMA_signal_1087, n2576}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2363 ( .ina ({new_AGEMA_signal_990, n2609}), .inb ({new_AGEMA_signal_957, n2765}), .clk ( clk ), .rnd ({Fresh[301], Fresh[300]}), .outt ({new_AGEMA_signal_1088, n2748}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) U2368 ( .a ({new_AGEMA_signal_1175, n2654}), .b ({new_AGEMA_signal_1375, n2674}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2378 ( .ina ({new_AGEMA_signal_983, n2815}), .inb ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .rnd ({Fresh[303], Fresh[302]}), .outt ({new_AGEMA_signal_1089, n2213}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2380 ( .ina ({new_AGEMA_signal_975, n2816}), .inb ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[305], Fresh[304]}), .outt ({new_AGEMA_signal_1090, n2215}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2384 ( .ina ({new_AGEMA_signal_969, n2712}), .inb ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .rnd ({Fresh[307], Fresh[306]}), .outt ({new_AGEMA_signal_1211, n2218}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2386 ( .ina ({new_AGEMA_signal_1012, n2298}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[309], Fresh[308]}), .outt ({new_AGEMA_signal_1212, n2219}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2405 ( .ina ({new_AGEMA_signal_1029, n2707}), .inb ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .rnd ({Fresh[311], Fresh[310]}), .outt ({new_AGEMA_signal_1217, n2240}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2407 ( .ina ({new_AGEMA_signal_1068, n2709}), .inb ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .rnd ({Fresh[313], Fresh[312]}), .outt ({new_AGEMA_signal_1218, n2561}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2408 ( .ina ({SI_s1[5], SI_s0[5]}), .inb ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .rnd ({Fresh[315], Fresh[314]}), .outt ({new_AGEMA_signal_1219, n2243}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2411 ( .ina ({new_AGEMA_signal_973, n2615}), .inb ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .rnd ({Fresh[317], Fresh[316]}), .outt ({new_AGEMA_signal_1220, n2245}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2422 ( .ina ({new_AGEMA_signal_1023, n2672}), .inb ({new_AGEMA_signal_1015, n2430}), .clk ( clk ), .rnd ({Fresh[319], Fresh[318]}), .outt ({new_AGEMA_signal_1221, n2540}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2423 ( .ina ({new_AGEMA_signal_966, n2261}), .inb ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .rnd ({Fresh[321], Fresh[320]}), .outt ({new_AGEMA_signal_1222, n2259}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2426 ( .ina ({new_AGEMA_signal_966, n2261}), .inb ({new_AGEMA_signal_991, n2661}), .clk ( clk ), .rnd ({Fresh[323], Fresh[322]}), .outt ({new_AGEMA_signal_1091, n2262}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2431 ( .ina ({new_AGEMA_signal_961, n2315}), .inb ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .rnd ({Fresh[325], Fresh[324]}), .outt ({new_AGEMA_signal_1092, n2266}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2432 ( .ina ({new_AGEMA_signal_1000, n2772}), .inb ({new_AGEMA_signal_943, n2796}), .clk ( clk ), .rnd ({Fresh[327], Fresh[326]}), .outt ({new_AGEMA_signal_1093, n2645}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2436 ( .ina ({SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .rnd ({Fresh[329], Fresh[328]}), .outt ({new_AGEMA_signal_1094, n2268}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2443 ( .ina ({new_AGEMA_signal_975, n2816}), .inb ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .rnd ({Fresh[331], Fresh[330]}), .outt ({new_AGEMA_signal_1225, n2278}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2448 ( .ina ({new_AGEMA_signal_951, n2791}), .inb ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .rnd ({Fresh[333], Fresh[332]}), .outt ({new_AGEMA_signal_1095, n2383}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2455 ( .ina ({new_AGEMA_signal_997, n2778}), .inb ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .rnd ({Fresh[335], Fresh[334]}), .outt ({new_AGEMA_signal_1228, n2774}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2458 ( .ina ({new_AGEMA_signal_1063, n2823}), .inb ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .rnd ({Fresh[337], Fresh[336]}), .outt ({new_AGEMA_signal_1229, n2287}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2470 ( .ina ({new_AGEMA_signal_960, n2519}), .inb ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .rnd ({Fresh[339], Fresh[338]}), .outt ({new_AGEMA_signal_1231, n2438}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2471 ( .ina ({new_AGEMA_signal_1012, n2298}), .inb ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .rnd ({Fresh[341], Fresh[340]}), .outt ({new_AGEMA_signal_1096, n2299}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2481 ( .ina ({new_AGEMA_signal_1050, n2766}), .inb ({new_AGEMA_signal_1054, n2313}), .clk ( clk ), .rnd ({Fresh[343], Fresh[342]}), .outt ({new_AGEMA_signal_1232, n2371}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2484 ( .ina ({new_AGEMA_signal_961, n2315}), .inb ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .rnd ({Fresh[345], Fresh[344]}), .outt ({new_AGEMA_signal_1018, n2316}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2486 ( .ina ({new_AGEMA_signal_1003, n2624}), .inb ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .rnd ({Fresh[347], Fresh[346]}), .outt ({new_AGEMA_signal_1098, n2318}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2492 ( .ina ({new_AGEMA_signal_964, n2708}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[349], Fresh[348]}), .outt ({new_AGEMA_signal_1235, n2325}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2494 ( .ina ({new_AGEMA_signal_964, n2708}), .inb ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .rnd ({Fresh[351], Fresh[350]}), .outt ({new_AGEMA_signal_1236, n2328}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2495 ( .ina ({new_AGEMA_signal_986, n2742}), .inb ({new_AGEMA_signal_981, n2723}), .clk ( clk ), .rnd ({Fresh[353], Fresh[352]}), .outt ({new_AGEMA_signal_1099, n2327}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2505 ( .ina ({new_AGEMA_signal_1025, n2737}), .inb ({new_AGEMA_signal_978, n2694}), .clk ( clk ), .rnd ({Fresh[355], Fresh[354]}), .outt ({new_AGEMA_signal_1237, n2343}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2510 ( .ina ({new_AGEMA_signal_1007, n2563}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[357], Fresh[356]}), .outt ({new_AGEMA_signal_1239, n2344}) ) ;
    and_HPC1 #(.security_order(1), .pipeline(0)) U2512 ( .ina ({new_AGEMA_signal_1002, n2395}), .inb ({new_AGEMA_signal_1013, n2346}), .clk ( clk ), .rnd ({Fresh[359], Fresh[358]}), .outt ({new_AGEMA_signal_1100, n2348}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2513 ( .ina ({new_AGEMA_signal_986, n2742}), .inb ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .rnd ({Fresh[361], Fresh[360]}), .outt ({new_AGEMA_signal_1101, n2347}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2520 ( .ina ({new_AGEMA_signal_978, n2694}), .inb ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .rnd ({Fresh[363], Fresh[362]}), .outt ({new_AGEMA_signal_1102, n2363}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2521 ( .ina ({new_AGEMA_signal_1067, n2809}), .inb ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[365], Fresh[364]}), .outt ({new_AGEMA_signal_1243, n2353}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2524 ( .ina ({new_AGEMA_signal_1058, n2818}), .inb ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .rnd ({Fresh[367], Fresh[366]}), .outt ({new_AGEMA_signal_1244, n2355}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2530 ( .ina ({new_AGEMA_signal_969, n2712}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[369], Fresh[368]}), .outt ({new_AGEMA_signal_1245, n2364}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2543 ( .ina ({SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1008, n2401}), .clk ( clk ), .rnd ({Fresh[371], Fresh[370]}), .outt ({new_AGEMA_signal_1103, n2415}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2558 ( .ina ({new_AGEMA_signal_1002, n2395}), .inb ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .rnd ({Fresh[373], Fresh[372]}), .outt ({new_AGEMA_signal_1104, n2700}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2563 ( .ina ({SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_988, n2400}), .clk ( clk ), .rnd ({Fresh[375], Fresh[374]}), .outt ({new_AGEMA_signal_1105, n2594}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2564 ( .ina ({new_AGEMA_signal_1008, n2401}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[377], Fresh[376]}), .outt ({new_AGEMA_signal_1106, n2402}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2585 ( .ina ({new_AGEMA_signal_969, n2712}), .inb ({new_AGEMA_signal_1063, n2823}), .clk ( clk ), .rnd ({Fresh[379], Fresh[378]}), .outt ({new_AGEMA_signal_1255, n2428}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2588 ( .ina ({new_AGEMA_signal_1015, n2430}), .inb ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .rnd ({Fresh[381], Fresh[380]}), .outt ({new_AGEMA_signal_1256, n2431}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2594 ( .ina ({new_AGEMA_signal_996, n2437}), .inb ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .rnd ({Fresh[383], Fresh[382]}), .outt ({new_AGEMA_signal_1107, n2483}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2599 ( .ina ({new_AGEMA_signal_1045, n2442}), .inb ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .rnd ({Fresh[385], Fresh[384]}), .outt ({new_AGEMA_signal_1258, n2443}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2606 ( .ina ({new_AGEMA_signal_1050, n2766}), .inb ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .rnd ({Fresh[387], Fresh[386]}), .outt ({new_AGEMA_signal_1259, n2693}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2608 ( .ina ({new_AGEMA_signal_998, n2452}), .inb ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .rnd ({Fresh[389], Fresh[388]}), .outt ({new_AGEMA_signal_1108, n2453}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2616 ( .ina ({new_AGEMA_signal_959, n2790}), .inb ({new_AGEMA_signal_1019, n2463}), .clk ( clk ), .rnd ({Fresh[391], Fresh[390]}), .outt ({new_AGEMA_signal_1109, n2464}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2620 ( .ina ({new_AGEMA_signal_982, n2725}), .inb ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .rnd ({Fresh[393], Fresh[392]}), .outt ({new_AGEMA_signal_1110, n2468}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2624 ( .ina ({new_AGEMA_signal_997, n2778}), .inb ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[395], Fresh[394]}), .outt ({new_AGEMA_signal_1111, n2473}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2625 ( .ina ({new_AGEMA_signal_983, n2815}), .inb ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .rnd ({Fresh[397], Fresh[396]}), .outt ({new_AGEMA_signal_1112, n2472}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2628 ( .ina ({new_AGEMA_signal_991, n2661}), .inb ({new_AGEMA_signal_1020, n2474}), .clk ( clk ), .rnd ({Fresh[399], Fresh[398]}), .outt ({new_AGEMA_signal_1113, n2475}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2632 ( .ina ({new_AGEMA_signal_945, n2810}), .inb ({new_AGEMA_signal_1065, n2828}), .clk ( clk ), .rnd ({Fresh[401], Fresh[400]}), .outt ({new_AGEMA_signal_1263, n2480}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2638 ( .ina ({new_AGEMA_signal_1037, n2577}), .inb ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .rnd ({Fresh[403], Fresh[402]}), .outt ({new_AGEMA_signal_1264, n2487}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2641 ( .ina ({new_AGEMA_signal_1006, n2616}), .inb ({new_AGEMA_signal_1001, n2824}), .clk ( clk ), .rnd ({Fresh[405], Fresh[404]}), .outt ({new_AGEMA_signal_1114, n2488}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2665 ( .ina ({new_AGEMA_signal_1035, n2786}), .inb ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .rnd ({Fresh[407], Fresh[406]}), .outt ({new_AGEMA_signal_1270, n2520}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2667 ( .ina ({new_AGEMA_signal_980, n2713}), .inb ({new_AGEMA_signal_993, n2587}), .clk ( clk ), .rnd ({Fresh[409], Fresh[408]}), .outt ({new_AGEMA_signal_1115, n2521}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2674 ( .ina ({new_AGEMA_signal_1025, n2737}), .inb ({new_AGEMA_signal_963, n2595}), .clk ( clk ), .rnd ({Fresh[411], Fresh[410]}), .outt ({new_AGEMA_signal_1271, n2531}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2689 ( .ina ({new_AGEMA_signal_1001, n2824}), .inb ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .rnd ({Fresh[413], Fresh[412]}), .outt ({new_AGEMA_signal_1273, n2553}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2691 ( .ina ({new_AGEMA_signal_978, n2694}), .inb ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .rnd ({Fresh[415], Fresh[414]}), .outt ({new_AGEMA_signal_1274, n2554}) ) ;
    and_HPC1 #(.security_order(1), .pipeline(0)) U2695 ( .ina ({new_AGEMA_signal_965, n2559}), .inb ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .rnd ({Fresh[417], Fresh[416]}), .outt ({new_AGEMA_signal_1116, n2560}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2698 ( .ina ({new_AGEMA_signal_1040, n2724}), .inb ({new_AGEMA_signal_1007, n2563}), .clk ( clk ), .rnd ({Fresh[419], Fresh[418]}), .outt ({new_AGEMA_signal_1275, n2564}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2714 ( .ina ({new_AGEMA_signal_1031, n2688}), .inb ({new_AGEMA_signal_978, n2694}), .clk ( clk ), .rnd ({Fresh[421], Fresh[420]}), .outt ({new_AGEMA_signal_1278, n2586}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2720 ( .ina ({new_AGEMA_signal_963, n2595}), .inb ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .rnd ({Fresh[423], Fresh[422]}), .outt ({new_AGEMA_signal_1117, n2597}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2721 ( .ina ({new_AGEMA_signal_1024, n2640}), .inb ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .rnd ({Fresh[425], Fresh[424]}), .outt ({new_AGEMA_signal_1280, n2596}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2723 ( .ina ({new_AGEMA_signal_1040, n2724}), .inb ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .rnd ({Fresh[427], Fresh[426]}), .outt ({new_AGEMA_signal_1281, n2598}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2725 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[429], Fresh[428]}), .outt ({new_AGEMA_signal_1021, n2599}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2732 ( .ina ({new_AGEMA_signal_1029, n2707}), .inb ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .rnd ({Fresh[431], Fresh[430]}), .outt ({new_AGEMA_signal_1283, n2610}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2734 ( .ina ({new_AGEMA_signal_1026, n2767}), .inb ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .rnd ({Fresh[433], Fresh[432]}), .outt ({new_AGEMA_signal_1284, n2614}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2735 ( .ina ({new_AGEMA_signal_1053, n2612}), .inb ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .rnd ({Fresh[435], Fresh[434]}), .outt ({new_AGEMA_signal_1285, n2613}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2737 ( .ina ({new_AGEMA_signal_1006, n2616}), .inb ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .rnd ({Fresh[437], Fresh[436]}), .outt ({new_AGEMA_signal_1119, n2617}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2742 ( .ina ({new_AGEMA_signal_1003, n2624}), .inb ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .rnd ({Fresh[439], Fresh[438]}), .outt ({new_AGEMA_signal_1120, n2629}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2751 ( .ina ({new_AGEMA_signal_971, n2641}), .inb ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .rnd ({Fresh[441], Fresh[440]}), .outt ({new_AGEMA_signal_1287, n2784}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2757 ( .ina ({new_AGEMA_signal_989, n2785}), .inb ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .rnd ({Fresh[443], Fresh[442]}), .outt ({new_AGEMA_signal_1121, n2650}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2775 ( .ina ({new_AGEMA_signal_949, n2760}), .inb ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .rnd ({Fresh[445], Fresh[444]}), .outt ({new_AGEMA_signal_1022, n2683}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2789 ( .ina ({new_AGEMA_signal_981, n2723}), .inb ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .rnd ({Fresh[447], Fresh[446]}), .outt ({new_AGEMA_signal_1294, n2711}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2790 ( .ina ({new_AGEMA_signal_1068, n2709}), .inb ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .rnd ({Fresh[449], Fresh[448]}), .outt ({new_AGEMA_signal_1295, n2710}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2792 ( .ina ({new_AGEMA_signal_980, n2713}), .inb ({new_AGEMA_signal_969, n2712}), .clk ( clk ), .rnd ({Fresh[451], Fresh[450]}), .outt ({new_AGEMA_signal_1122, n2714}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2797 ( .ina ({new_AGEMA_signal_959, n2790}), .inb ({new_AGEMA_signal_1011, n2721}), .clk ( clk ), .rnd ({Fresh[453], Fresh[452]}), .outt ({new_AGEMA_signal_1123, n2722}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2799 ( .ina ({new_AGEMA_signal_982, n2725}), .inb ({new_AGEMA_signal_1040, n2724}), .clk ( clk ), .rnd ({Fresh[455], Fresh[454]}), .outt ({new_AGEMA_signal_1297, n2726}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2806 ( .ina ({new_AGEMA_signal_1025, n2737}), .inb ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .rnd ({Fresh[457], Fresh[456]}), .outt ({new_AGEMA_signal_1298, n2738}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2822 ( .ina ({new_AGEMA_signal_1026, n2767}), .inb ({new_AGEMA_signal_1050, n2766}), .clk ( clk ), .rnd ({Fresh[459], Fresh[458]}), .outt ({new_AGEMA_signal_1301, n2768}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2828 ( .ina ({new_AGEMA_signal_997, n2778}), .inb ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .rnd ({Fresh[461], Fresh[460]}), .outt ({new_AGEMA_signal_1124, n2782}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2829 ( .ina ({new_AGEMA_signal_976, n2780}), .inb ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .rnd ({Fresh[463], Fresh[462]}), .outt ({new_AGEMA_signal_1125, n2781}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2832 ( .ina ({new_AGEMA_signal_1035, n2786}), .inb ({new_AGEMA_signal_989, n2785}), .clk ( clk ), .rnd ({Fresh[465], Fresh[464]}), .outt ({new_AGEMA_signal_1303, n2787}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2834 ( .ina ({new_AGEMA_signal_959, n2790}), .inb ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .rnd ({Fresh[467], Fresh[466]}), .outt ({new_AGEMA_signal_1304, n2794}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2835 ( .ina ({new_AGEMA_signal_1039, n2792}), .inb ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .rnd ({Fresh[469], Fresh[468]}), .outt ({new_AGEMA_signal_1305, n2793}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2844 ( .ina ({new_AGEMA_signal_945, n2810}), .inb ({new_AGEMA_signal_1067, n2809}), .clk ( clk ), .rnd ({Fresh[471], Fresh[470]}), .outt ({new_AGEMA_signal_1306, n2812}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2847 ( .ina ({new_AGEMA_signal_975, n2816}), .inb ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .rnd ({Fresh[473], Fresh[472]}), .outt ({new_AGEMA_signal_1126, n2820}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2851 ( .ina ({new_AGEMA_signal_1001, n2824}), .inb ({new_AGEMA_signal_1063, n2823}), .clk ( clk ), .rnd ({Fresh[475], Fresh[474]}), .outt ({new_AGEMA_signal_1308, n2825}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1960 ( .ina ({new_AGEMA_signal_1127, n2575}), .inb ({new_AGEMA_signal_1128, n1962}), .clk ( clk ), .rnd ({Fresh[477], Fresh[476]}), .outt ({new_AGEMA_signal_1309, n1924}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1967 ( .ina ({new_AGEMA_signal_1129, n1922}), .inb ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .rnd ({Fresh[479], Fresh[478]}), .outt ({new_AGEMA_signal_1310, n1923}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1981 ( .ina ({new_AGEMA_signal_1130, n1926}), .inb ({new_AGEMA_signal_1131, n1925}), .clk ( clk ), .rnd ({Fresh[481], Fresh[480]}), .outt ({new_AGEMA_signal_1311, n1927}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1993 ( .ina ({new_AGEMA_signal_1133, n2734}), .inb ({new_AGEMA_signal_1134, n2763}), .clk ( clk ), .rnd ({Fresh[483], Fresh[482]}), .outt ({new_AGEMA_signal_1312, n1929}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2007 ( .ina ({SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .rnd ({Fresh[485], Fresh[484]}), .outt ({new_AGEMA_signal_1313, n2665}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2011 ( .ina ({SI_s1[6], SI_s0[6]}), .inb ({new_AGEMA_signal_1136, n1937}), .clk ( clk ), .rnd ({Fresh[487], Fresh[486]}), .outt ({new_AGEMA_signal_1314, n1938}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2019 ( .ina ({new_AGEMA_signal_1041, n2174}), .inb ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .rnd ({Fresh[489], Fresh[488]}), .outt ({new_AGEMA_signal_1315, n2235}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2023 ( .ina ({SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1042, n1942}), .clk ( clk ), .rnd ({Fresh[491], Fresh[490]}), .outt ({new_AGEMA_signal_1137, n1943}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2027 ( .ina ({new_AGEMA_signal_1043, n2676}), .inb ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[493], Fresh[492]}), .outt ({new_AGEMA_signal_1138, n1946}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2031 ( .ina ({new_AGEMA_signal_1044, n2570}), .inb ({new_AGEMA_signal_1139, n1944}), .clk ( clk ), .rnd ({Fresh[495], Fresh[494]}), .outt ({new_AGEMA_signal_1316, n1945}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2034 ( .ina ({new_AGEMA_signal_1039, n2792}), .inb ({new_AGEMA_signal_1133, n2734}), .clk ( clk ), .rnd ({Fresh[497], Fresh[496]}), .outt ({new_AGEMA_signal_1317, n1956}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2040 ( .ina ({new_AGEMA_signal_1140, n1950}), .inb ({new_AGEMA_signal_1046, n1949}), .clk ( clk ), .rnd ({Fresh[499], Fresh[498]}), .outt ({new_AGEMA_signal_1318, n1951}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2048 ( .ina ({new_AGEMA_signal_1141, n2662}), .inb ({new_AGEMA_signal_1048, n2627}), .clk ( clk ), .rnd ({Fresh[501], Fresh[500]}), .outt ({new_AGEMA_signal_1319, n1952}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2057 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1142, n2088}), .clk ( clk ), .rnd ({Fresh[503], Fresh[502]}), .outt ({new_AGEMA_signal_1320, n2687}) ) ;
    or_HPC1 #(.security_order(1), .pipeline(0)) U2061 ( .ina ({new_AGEMA_signal_1128, n1962}), .inb ({new_AGEMA_signal_993, n2587}), .clk ( clk ), .rnd ({Fresh[505], Fresh[504]}), .outt ({new_AGEMA_signal_1321, n1966}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2064 ( .ina ({new_AGEMA_signal_1051, n2736}), .inb ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .rnd ({Fresh[507], Fresh[506]}), .outt ({new_AGEMA_signal_1143, n1963}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2077 ( .ina ({new_AGEMA_signal_1323, n2720}), .inb ({new_AGEMA_signal_1324, n2417}), .clk ( clk ), .rnd ({Fresh[509], Fresh[508]}), .outt ({new_AGEMA_signal_1480, n1968}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2082 ( .ina ({new_AGEMA_signal_1146, n2505}), .inb ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .rnd ({Fresh[511], Fresh[510]}), .outt ({new_AGEMA_signal_1325, n2684}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2088 ( .ina ({new_AGEMA_signal_964, n2708}), .inb ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .rnd ({Fresh[513], Fresh[512]}), .outt ({new_AGEMA_signal_1326, n1972}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2092 ( .ina ({new_AGEMA_signal_1058, n2818}), .inb ({new_AGEMA_signal_1059, n2190}), .clk ( clk ), .rnd ({Fresh[515], Fresh[514]}), .outt ({new_AGEMA_signal_1149, n1971}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2099 ( .ina ({new_AGEMA_signal_959, n2790}), .inb ({new_AGEMA_signal_1150, n2535}), .clk ( clk ), .rnd ({Fresh[517], Fresh[516]}), .outt ({new_AGEMA_signal_1327, n1974}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2106 ( .ina ({new_AGEMA_signal_1135, n2732}), .inb ({new_AGEMA_signal_958, n2635}), .clk ( clk ), .rnd ({Fresh[519], Fresh[518]}), .outt ({new_AGEMA_signal_1328, n1979}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2112 ( .ina ({new_AGEMA_signal_1035, n2786}), .inb ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .rnd ({Fresh[521], Fresh[520]}), .outt ({new_AGEMA_signal_1152, n1985}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2121 ( .ina ({new_AGEMA_signal_1154, n1992}), .inb ({new_AGEMA_signal_1155, n1991}), .clk ( clk ), .rnd ({Fresh[523], Fresh[522]}), .outt ({new_AGEMA_signal_1330, n1994}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2126 ( .ina ({new_AGEMA_signal_988, n2400}), .inb ({new_AGEMA_signal_1156, n1995}), .clk ( clk ), .rnd ({Fresh[525], Fresh[524]}), .outt ({new_AGEMA_signal_1331, n1996}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2136 ( .ina ({SI_s1[1], SI_s0[1]}), .inb ({new_AGEMA_signal_1158, n2003}), .clk ( clk ), .rnd ({Fresh[527], Fresh[526]}), .outt ({new_AGEMA_signal_1332, n2137}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2142 ( .ina ({new_AGEMA_signal_983, n2815}), .inb ({new_AGEMA_signal_1160, n2572}), .clk ( clk ), .rnd ({Fresh[529], Fresh[528]}), .outt ({new_AGEMA_signal_1333, n2006}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2144 ( .ina ({new_AGEMA_signal_981, n2723}), .inb ({new_AGEMA_signal_1161, n2004}), .clk ( clk ), .rnd ({Fresh[531], Fresh[530]}), .outt ({new_AGEMA_signal_1334, n2005}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2152 ( .ina ({new_AGEMA_signal_1068, n2709}), .inb ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .rnd ({Fresh[533], Fresh[532]}), .outt ({new_AGEMA_signal_1335, n2013}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2160 ( .ina ({new_AGEMA_signal_987, n2753}), .inb ({new_AGEMA_signal_1070, n2227}), .clk ( clk ), .rnd ({Fresh[535], Fresh[534]}), .outt ({new_AGEMA_signal_1165, n2020}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2164 ( .ina ({new_AGEMA_signal_1062, n2817}), .inb ({new_AGEMA_signal_1008, n2401}), .clk ( clk ), .rnd ({Fresh[537], Fresh[536]}), .outt ({new_AGEMA_signal_1166, n2023}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2168 ( .ina ({new_AGEMA_signal_1009, n2027}), .inb ({new_AGEMA_signal_957, n2765}), .clk ( clk ), .rnd ({Fresh[539], Fresh[538]}), .outt ({new_AGEMA_signal_1071, n2028}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2172 ( .ina ({new_AGEMA_signal_1167, n2214}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[541], Fresh[540]}), .outt ({new_AGEMA_signal_1337, n2033}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2175 ( .ina ({new_AGEMA_signal_1169, n2376}), .inb ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .rnd ({Fresh[543], Fresh[542]}), .outt ({new_AGEMA_signal_1338, n2031}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2184 ( .ina ({new_AGEMA_signal_1048, n2627}), .inb ({new_AGEMA_signal_1170, n2039}), .clk ( clk ), .rnd ({Fresh[545], Fresh[544]}), .outt ({new_AGEMA_signal_1339, n2040}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2187 ( .ina ({new_AGEMA_signal_994, n2643}), .inb ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .rnd ({Fresh[547], Fresh[546]}), .outt ({new_AGEMA_signal_1171, n2050}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2193 ( .ina ({new_AGEMA_signal_1007, n2563}), .inb ({new_AGEMA_signal_1174, n2044}), .clk ( clk ), .rnd ({Fresh[549], Fresh[548]}), .outt ({new_AGEMA_signal_1340, n2045}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2199 ( .ina ({new_AGEMA_signal_1175, n2654}), .inb ({new_AGEMA_signal_958, n2635}), .clk ( clk ), .rnd ({Fresh[551], Fresh[550]}), .outt ({new_AGEMA_signal_1341, n2051}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2203 ( .ina ({new_AGEMA_signal_1053, n2612}), .inb ({new_AGEMA_signal_1176, n2055}), .clk ( clk ), .rnd ({Fresh[553], Fresh[552]}), .outt ({new_AGEMA_signal_1342, n2056}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2209 ( .ina ({new_AGEMA_signal_1178, n2407}), .inb ({new_AGEMA_signal_1001, n2824}), .clk ( clk ), .rnd ({Fresh[555], Fresh[554]}), .outt ({new_AGEMA_signal_1343, n2060}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2215 ( .ina ({new_AGEMA_signal_975, n2816}), .inb ({new_AGEMA_signal_1175, n2654}), .clk ( clk ), .rnd ({Fresh[557], Fresh[556]}), .outt ({new_AGEMA_signal_1344, n2066}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2217 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .rnd ({Fresh[559], Fresh[558]}), .outt ({new_AGEMA_signal_1345, n2065}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2221 ( .ina ({new_AGEMA_signal_1181, n2068}), .inb ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .rnd ({Fresh[561], Fresh[560]}), .outt ({new_AGEMA_signal_1346, n2069}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2226 ( .ina ({new_AGEMA_signal_979, n2073}), .inb ({new_AGEMA_signal_1182, n2252}), .clk ( clk ), .rnd ({Fresh[563], Fresh[562]}), .outt ({new_AGEMA_signal_1347, n2074}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2235 ( .ina ({new_AGEMA_signal_1076, n2081}), .inb ({new_AGEMA_signal_1183, n2080}), .clk ( clk ), .rnd ({Fresh[565], Fresh[564]}), .outt ({new_AGEMA_signal_1348, n2082}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2240 ( .ina ({new_AGEMA_signal_981, n2723}), .inb ({new_AGEMA_signal_1185, n2083}), .clk ( clk ), .rnd ({Fresh[567], Fresh[566]}), .outt ({new_AGEMA_signal_1349, n2084}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2242 ( .ina ({new_AGEMA_signal_1163, n2533}), .inb ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[569], Fresh[568]}), .outt ({new_AGEMA_signal_1350, n2085}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2245 ( .ina ({new_AGEMA_signal_960, n2519}), .inb ({new_AGEMA_signal_1186, n2562}), .clk ( clk ), .rnd ({Fresh[571], Fresh[570]}), .outt ({new_AGEMA_signal_1351, n2131}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2248 ( .ina ({new_AGEMA_signal_1142, n2088}), .inb ({new_AGEMA_signal_1078, n2087}), .clk ( clk ), .rnd ({Fresh[573], Fresh[572]}), .outt ({new_AGEMA_signal_1352, n2089}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2252 ( .ina ({new_AGEMA_signal_955, n2630}), .inb ({new_AGEMA_signal_1187, n2156}), .clk ( clk ), .rnd ({Fresh[575], Fresh[574]}), .outt ({new_AGEMA_signal_1353, n2330}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2254 ( .ina ({new_AGEMA_signal_1006, n2616}), .inb ({new_AGEMA_signal_1132, n2151}), .clk ( clk ), .rnd ({Fresh[577], Fresh[576]}), .outt ({new_AGEMA_signal_1354, n2092}) ) ;
    or_HPC1 #(.security_order(1), .pipeline(0)) U2256 ( .ina ({new_AGEMA_signal_1144, n2761}), .inb ({new_AGEMA_signal_1147, n2359}), .clk ( clk ), .rnd ({Fresh[579], Fresh[578]}), .outt ({new_AGEMA_signal_1355, n2094}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2261 ( .ina ({new_AGEMA_signal_1057, n2101}), .inb ({new_AGEMA_signal_1188, n2100}), .clk ( clk ), .rnd ({Fresh[581], Fresh[580]}), .outt ({new_AGEMA_signal_1356, n2160}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2265 ( .ina ({new_AGEMA_signal_1038, n2492}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[583], Fresh[582]}), .outt ({new_AGEMA_signal_1189, n2504}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2271 ( .ina ({new_AGEMA_signal_1324, n2417}), .inb ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .rnd ({Fresh[585], Fresh[584]}), .outt ({new_AGEMA_signal_1504, n2114}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2273 ( .ina ({new_AGEMA_signal_1047, n2677}), .inb ({new_AGEMA_signal_981, n2723}), .clk ( clk ), .rnd ({Fresh[587], Fresh[586]}), .outt ({new_AGEMA_signal_1190, n2115}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2280 ( .ina ({new_AGEMA_signal_951, n2791}), .inb ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .rnd ({Fresh[589], Fresh[588]}), .outt ({new_AGEMA_signal_1358, n2291}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2281 ( .ina ({SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .rnd ({Fresh[591], Fresh[590]}), .outt ({new_AGEMA_signal_1192, n2119}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2291 ( .ina ({new_AGEMA_signal_976, n2780}), .inb ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .rnd ({Fresh[593], Fresh[592]}), .outt ({new_AGEMA_signal_1195, n2130}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2292 ( .ina ({new_AGEMA_signal_1062, n2817}), .inb ({new_AGEMA_signal_1034, n2631}), .clk ( clk ), .rnd ({Fresh[595], Fresh[594]}), .outt ({new_AGEMA_signal_1196, n2129}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2295 ( .ina ({new_AGEMA_signal_1081, n2647}), .inb ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .rnd ({Fresh[597], Fresh[596]}), .outt ({new_AGEMA_signal_1197, n2150}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2298 ( .ina ({new_AGEMA_signal_1038, n2492}), .inb ({new_AGEMA_signal_1082, n2132}), .clk ( clk ), .rnd ({Fresh[599], Fresh[598]}), .outt ({new_AGEMA_signal_1198, n2133}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2302 ( .ina ({new_AGEMA_signal_1163, n2533}), .inb ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .rnd ({Fresh[601], Fresh[600]}), .outt ({new_AGEMA_signal_1361, n2136}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2306 ( .ina ({new_AGEMA_signal_1160, n2572}), .inb ({new_AGEMA_signal_1200, n2138}), .clk ( clk ), .rnd ({Fresh[603], Fresh[602]}), .outt ({new_AGEMA_signal_1362, n2139}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2313 ( .ina ({new_AGEMA_signal_1040, n2724}), .inb ({new_AGEMA_signal_1201, n2555}), .clk ( clk ), .rnd ({Fresh[605], Fresh[604]}), .outt ({new_AGEMA_signal_1363, n2144}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2318 ( .ina ({new_AGEMA_signal_1132, n2151}), .inb ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .rnd ({Fresh[607], Fresh[606]}), .outt ({new_AGEMA_signal_1364, n2152}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2321 ( .ina ({new_AGEMA_signal_1048, n2627}), .inb ({new_AGEMA_signal_1187, n2156}), .clk ( clk ), .rnd ({Fresh[609], Fresh[608]}), .outt ({new_AGEMA_signal_1365, n2170}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2323 ( .ina ({new_AGEMA_signal_1202, n2429}), .inb ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .rnd ({Fresh[611], Fresh[610]}), .outt ({new_AGEMA_signal_1366, n2157}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2329 ( .ina ({new_AGEMA_signal_977, n2317}), .inb ({new_AGEMA_signal_1083, n2162}), .clk ( clk ), .rnd ({Fresh[613], Fresh[612]}), .outt ({new_AGEMA_signal_1203, n2163}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2335 ( .ina ({new_AGEMA_signal_1073, n2171}), .inb ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .rnd ({Fresh[615], Fresh[614]}), .outt ({new_AGEMA_signal_1368, n2172}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2338 ( .ina ({SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1014, n2545}), .clk ( clk ), .rnd ({Fresh[617], Fresh[616]}), .outt ({new_AGEMA_signal_1084, n2186}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2339 ( .ina ({new_AGEMA_signal_959, n2790}), .inb ({new_AGEMA_signal_1168, n2290}), .clk ( clk ), .rnd ({Fresh[619], Fresh[618]}), .outt ({new_AGEMA_signal_1369, n2181}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2344 ( .ina ({new_AGEMA_signal_1204, n2176}), .inb ({new_AGEMA_signal_1205, n2175}), .clk ( clk ), .rnd ({Fresh[621], Fresh[620]}), .outt ({new_AGEMA_signal_1370, n2177}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2349 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1016, n2182}), .clk ( clk ), .rnd ({Fresh[623], Fresh[622]}), .outt ({new_AGEMA_signal_1086, n2183}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2354 ( .ina ({new_AGEMA_signal_1031, n2688}), .inb ({new_AGEMA_signal_1206, n2188}), .clk ( clk ), .rnd ({Fresh[625], Fresh[624]}), .outt ({new_AGEMA_signal_1371, n2195}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2356 ( .ina ({new_AGEMA_signal_1059, n2190}), .inb ({new_AGEMA_signal_1207, n2189}), .clk ( clk ), .rnd ({Fresh[627], Fresh[626]}), .outt ({new_AGEMA_signal_1372, n2193}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2358 ( .ina ({new_AGEMA_signal_990, n2609}), .inb ({new_AGEMA_signal_1208, n2446}), .clk ( clk ), .rnd ({Fresh[629], Fresh[628]}), .outt ({new_AGEMA_signal_1373, n2191}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2364 ( .ina ({new_AGEMA_signal_1087, n2576}), .inb ({new_AGEMA_signal_1088, n2748}), .clk ( clk ), .rnd ({Fresh[631], Fresh[630]}), .outt ({new_AGEMA_signal_1209, n2196}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2367 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1146, n2505}), .clk ( clk ), .rnd ({Fresh[633], Fresh[632]}), .outt ({new_AGEMA_signal_1374, n2201}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2369 ( .ina ({new_AGEMA_signal_1375, n2674}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[635], Fresh[634]}), .outt ({new_AGEMA_signal_1515, n2200}) ) ;
    mux2_HPC1 #(.security_order(1), .pipeline(0)) U2371 ( .ins ({new_AGEMA_signal_953, n2813}), .inb ({new_AGEMA_signal_1133, n2734}), .ina ({new_AGEMA_signal_1324, n2417}), .clk ( clk ), .rnd ({Fresh[637], Fresh[636]}), .outt ({new_AGEMA_signal_1516, n2202}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2379 ( .ina ({new_AGEMA_signal_1167, n2214}), .inb ({new_AGEMA_signal_1089, n2213}), .clk ( clk ), .rnd ({Fresh[639], Fresh[638]}), .outt ({new_AGEMA_signal_1376, n2217}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2381 ( .ina ({new_AGEMA_signal_1024, n2640}), .inb ({new_AGEMA_signal_1090, n2215}), .clk ( clk ), .rnd ({Fresh[641], Fresh[640]}), .outt ({new_AGEMA_signal_1210, n2216}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2385 ( .ina ({new_AGEMA_signal_1211, n2218}), .inb ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .rnd ({Fresh[643], Fresh[642]}), .outt ({new_AGEMA_signal_1377, n2222}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2387 ( .ina ({new_AGEMA_signal_1199, n2220}), .inb ({new_AGEMA_signal_1212, n2219}), .clk ( clk ), .rnd ({Fresh[645], Fresh[644]}), .outt ({new_AGEMA_signal_1378, n2221}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2391 ( .ina ({new_AGEMA_signal_1048, n2627}), .inb ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .rnd ({Fresh[647], Fresh[646]}), .outt ({new_AGEMA_signal_1213, n2226}) ) ;
    mux2_HPC1 #(.security_order(1), .pipeline(0)) U2393 ( .ins ({new_AGEMA_signal_953, n2813}), .inb ({new_AGEMA_signal_1056, n2651}), .ina ({new_AGEMA_signal_1070, n2227}), .clk ( clk ), .rnd ({Fresh[649], Fresh[648]}), .outt ({new_AGEMA_signal_1214, n2228}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2397 ( .ina ({new_AGEMA_signal_987, n2753}), .inb ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .rnd ({Fresh[651], Fresh[650]}), .outt ({new_AGEMA_signal_1215, n2237}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2398 ( .ina ({new_AGEMA_signal_1324, n2417}), .inb ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .rnd ({Fresh[653], Fresh[652]}), .outt ({new_AGEMA_signal_1520, n2233}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2403 ( .ina ({new_AGEMA_signal_1017, n2777}), .inb ({new_AGEMA_signal_1034, n2631}), .clk ( clk ), .rnd ({Fresh[655], Fresh[654]}), .outt ({new_AGEMA_signal_1216, n2238}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2406 ( .ina ({new_AGEMA_signal_1157, n2241}), .inb ({new_AGEMA_signal_1217, n2240}), .clk ( clk ), .rnd ({Fresh[657], Fresh[656]}), .outt ({new_AGEMA_signal_1380, n2248}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2409 ( .ina ({new_AGEMA_signal_1218, n2561}), .inb ({new_AGEMA_signal_1219, n2243}), .clk ( clk ), .rnd ({Fresh[659], Fresh[658]}), .outt ({new_AGEMA_signal_1381, n2244}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2414 ( .ina ({new_AGEMA_signal_1169, n2376}), .inb ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .rnd ({Fresh[661], Fresh[660]}), .outt ({new_AGEMA_signal_1382, n2249}) ) ;
    mux2_HPC1 #(.security_order(1), .pipeline(0)) U2417 ( .ins ({new_AGEMA_signal_953, n2813}), .inb ({new_AGEMA_signal_1182, n2252}), .ina ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .rnd ({Fresh[663], Fresh[662]}), .outt ({new_AGEMA_signal_1383, n2253}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2424 ( .ina ({new_AGEMA_signal_1163, n2533}), .inb ({new_AGEMA_signal_1222, n2259}), .clk ( clk ), .rnd ({Fresh[665], Fresh[664]}), .outt ({new_AGEMA_signal_1384, n2260}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2429 ( .ina ({new_AGEMA_signal_1324, n2417}), .inb ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .rnd ({Fresh[667], Fresh[666]}), .outt ({new_AGEMA_signal_1524, n2273}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2430 ( .ina ({new_AGEMA_signal_991, n2661}), .inb ({new_AGEMA_signal_1323, n2720}), .clk ( clk ), .rnd ({Fresh[669], Fresh[668]}), .outt ({new_AGEMA_signal_1525, n2752}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2433 ( .ina ({new_AGEMA_signal_1093, n2645}), .inb ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .rnd ({Fresh[671], Fresh[670]}), .outt ({new_AGEMA_signal_1223, n2265}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2437 ( .ina ({new_AGEMA_signal_947, n2462}), .inb ({new_AGEMA_signal_1094, n2268}), .clk ( clk ), .rnd ({Fresh[673], Fresh[672]}), .outt ({new_AGEMA_signal_1224, n2269}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2444 ( .ina ({new_AGEMA_signal_982, n2725}), .inb ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .rnd ({Fresh[675], Fresh[674]}), .outt ({new_AGEMA_signal_1226, n2277}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2449 ( .ina ({new_AGEMA_signal_978, n2694}), .inb ({new_AGEMA_signal_1095, n2383}), .clk ( clk ), .rnd ({Fresh[677], Fresh[676]}), .outt ({new_AGEMA_signal_1227, n2282}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2452 ( .ina ({new_AGEMA_signal_1051, n2736}), .inb ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .rnd ({Fresh[679], Fresh[678]}), .outt ({new_AGEMA_signal_1389, n2284}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2456 ( .ina ({new_AGEMA_signal_1228, n2774}), .inb ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .rnd ({Fresh[681], Fresh[680]}), .outt ({new_AGEMA_signal_1390, n2459}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2459 ( .ina ({SI_s1[6], SI_s0[6]}), .inb ({new_AGEMA_signal_1229, n2287}), .clk ( clk ), .rnd ({Fresh[683], Fresh[682]}), .outt ({new_AGEMA_signal_1391, n2288}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2462 ( .ina ({SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1144, n2761}), .clk ( clk ), .rnd ({Fresh[685], Fresh[684]}), .outt ({new_AGEMA_signal_1392, n2458}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2464 ( .ina ({new_AGEMA_signal_977, n2317}), .inb ({new_AGEMA_signal_1168, n2290}), .clk ( clk ), .rnd ({Fresh[687], Fresh[686]}), .outt ({new_AGEMA_signal_1393, n2293}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2467 ( .ina ({new_AGEMA_signal_1006, n2616}), .inb ({new_AGEMA_signal_1074, n2642}), .clk ( clk ), .rnd ({Fresh[689], Fresh[688]}), .outt ({new_AGEMA_signal_1230, n2294}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2472 ( .ina ({new_AGEMA_signal_1231, n2438}), .inb ({new_AGEMA_signal_1096, n2299}), .clk ( clk ), .rnd ({Fresh[691], Fresh[690]}), .outt ({new_AGEMA_signal_1394, n2300}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2480 ( .ina ({new_AGEMA_signal_1133, n2734}), .inb ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .rnd ({Fresh[693], Fresh[692]}), .outt ({new_AGEMA_signal_1395, n2323}) ) ;
    and_HPC1 #(.security_order(1), .pipeline(0)) U2482 ( .ina ({new_AGEMA_signal_1055, n2571}), .inb ({new_AGEMA_signal_1232, n2371}), .clk ( clk ), .rnd ({Fresh[695], Fresh[694]}), .outt ({new_AGEMA_signal_1396, n2314}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2485 ( .ina ({new_AGEMA_signal_1018, n2316}), .inb ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .rnd ({Fresh[697], Fresh[696]}), .outt ({new_AGEMA_signal_1097, n2319}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2491 ( .ina ({new_AGEMA_signal_1074, n2642}), .inb ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .rnd ({Fresh[699], Fresh[698]}), .outt ({new_AGEMA_signal_1234, n2326}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2496 ( .ina ({new_AGEMA_signal_1236, n2328}), .inb ({new_AGEMA_signal_1099, n2327}), .clk ( clk ), .rnd ({Fresh[701], Fresh[700]}), .outt ({new_AGEMA_signal_1398, n2329}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2501 ( .ina ({new_AGEMA_signal_1324, n2417}), .inb ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .rnd ({Fresh[703], Fresh[702]}), .outt ({new_AGEMA_signal_1537, n2335}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2506 ( .ina ({new_AGEMA_signal_1068, n2709}), .inb ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .rnd ({Fresh[705], Fresh[704]}), .outt ({new_AGEMA_signal_1399, n2341}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2507 ( .ina ({new_AGEMA_signal_945, n2810}), .inb ({new_AGEMA_signal_1051, n2736}), .clk ( clk ), .rnd ({Fresh[707], Fresh[706]}), .outt ({new_AGEMA_signal_1238, n2340}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2514 ( .ina ({new_AGEMA_signal_1100, n2348}), .inb ({new_AGEMA_signal_1101, n2347}), .clk ( clk ), .rnd ({Fresh[709], Fresh[708]}), .outt ({new_AGEMA_signal_1240, n2349}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2517 ( .ina ({new_AGEMA_signal_1003, n2624}), .inb ({new_AGEMA_signal_1061, n2690}), .clk ( clk ), .rnd ({Fresh[711], Fresh[710]}), .outt ({new_AGEMA_signal_1241, n2375}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2518 ( .ina ({new_AGEMA_signal_1040, n2724}), .inb ({new_AGEMA_signal_1051, n2736}), .clk ( clk ), .rnd ({Fresh[713], Fresh[712]}), .outt ({new_AGEMA_signal_1242, n2352}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2522 ( .ina ({new_AGEMA_signal_1243, n2353}), .inb ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .rnd ({Fresh[715], Fresh[714]}), .outt ({new_AGEMA_signal_1401, n2354}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2525 ( .ina ({new_AGEMA_signal_1004, n2356}), .inb ({new_AGEMA_signal_1244, n2355}), .clk ( clk ), .rnd ({Fresh[717], Fresh[716]}), .outt ({new_AGEMA_signal_1402, n2357}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2527 ( .ina ({new_AGEMA_signal_1147, n2359}), .inb ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .rnd ({Fresh[719], Fresh[718]}), .outt ({new_AGEMA_signal_1403, n2360}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2534 ( .ina ({SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .rnd ({Fresh[721], Fresh[720]}), .outt ({new_AGEMA_signal_1540, n2369}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2536 ( .ina ({new_AGEMA_signal_1232, n2371}), .inb ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .rnd ({Fresh[723], Fresh[722]}), .outt ({new_AGEMA_signal_1404, n2372}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2539 ( .ina ({new_AGEMA_signal_1087, n2576}), .inb ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .rnd ({Fresh[725], Fresh[724]}), .outt ({new_AGEMA_signal_1405, n2377}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2544 ( .ina ({new_AGEMA_signal_990, n2609}), .inb ({new_AGEMA_signal_1103, n2415}), .clk ( clk ), .rnd ({Fresh[727], Fresh[726]}), .outt ({new_AGEMA_signal_1246, n2467}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2545 ( .ina ({new_AGEMA_signal_1050, n2766}), .inb ({new_AGEMA_signal_1095, n2383}), .clk ( clk ), .rnd ({Fresh[729], Fresh[728]}), .outt ({new_AGEMA_signal_1247, n2385}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2546 ( .ina ({new_AGEMA_signal_1056, n2651}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[731], Fresh[730]}), .outt ({new_AGEMA_signal_1248, n2384}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2548 ( .ina ({new_AGEMA_signal_981, n2723}), .inb ({new_AGEMA_signal_1202, n2429}), .clk ( clk ), .rnd ({Fresh[733], Fresh[732]}), .outt ({new_AGEMA_signal_1407, n2386}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2552 ( .ina ({new_AGEMA_signal_1031, n2688}), .inb ({new_AGEMA_signal_1081, n2647}), .clk ( clk ), .rnd ({Fresh[735], Fresh[734]}), .outt ({new_AGEMA_signal_1249, n2394}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2553 ( .ina ({new_AGEMA_signal_1056, n2651}), .inb ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .rnd ({Fresh[737], Fresh[736]}), .outt ({new_AGEMA_signal_1250, n2391}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2554 ( .ina ({new_AGEMA_signal_1146, n2505}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[739], Fresh[738]}), .outt ({new_AGEMA_signal_1408, n2390}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2559 ( .ina ({new_AGEMA_signal_1006, n2616}), .inb ({new_AGEMA_signal_1104, n2700}), .clk ( clk ), .rnd ({Fresh[741], Fresh[740]}), .outt ({new_AGEMA_signal_1251, n2396}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2562 ( .ina ({new_AGEMA_signal_1026, n2767}), .inb ({new_AGEMA_signal_1231, n2438}), .clk ( clk ), .rnd ({Fresh[743], Fresh[742]}), .outt ({new_AGEMA_signal_1409, n2406}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2565 ( .ina ({new_AGEMA_signal_1105, n2594}), .inb ({new_AGEMA_signal_1106, n2402}), .clk ( clk ), .rnd ({Fresh[745], Fresh[744]}), .outt ({new_AGEMA_signal_1252, n2403}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2569 ( .ina ({new_AGEMA_signal_1178, n2407}), .inb ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .rnd ({Fresh[747], Fresh[746]}), .outt ({new_AGEMA_signal_1411, n2408}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2573 ( .ina ({new_AGEMA_signal_1145, n2412}), .inb ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .rnd ({Fresh[749], Fresh[748]}), .outt ({new_AGEMA_signal_1412, n2574}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2574 ( .ina ({new_AGEMA_signal_1077, n2498}), .inb ({new_AGEMA_signal_1007, n2563}), .clk ( clk ), .rnd ({Fresh[751], Fresh[750]}), .outt ({new_AGEMA_signal_1253, n2413}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2577 ( .ina ({new_AGEMA_signal_1103, n2415}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[753], Fresh[752]}), .outt ({new_AGEMA_signal_1254, n2416}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2586 ( .ina ({new_AGEMA_signal_1255, n2428}), .inb ({new_AGEMA_signal_971, n2641}), .clk ( clk ), .rnd ({Fresh[755], Fresh[754]}), .outt ({new_AGEMA_signal_1414, n2433}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2587 ( .ina ({SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1202, n2429}), .clk ( clk ), .rnd ({Fresh[757], Fresh[756]}), .outt ({new_AGEMA_signal_1415, n2689}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2591 ( .ina ({new_AGEMA_signal_1081, n2647}), .inb ({new_AGEMA_signal_1038, n2492}), .clk ( clk ), .rnd ({Fresh[759], Fresh[758]}), .outt ({new_AGEMA_signal_1257, n2434}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2595 ( .ina ({new_AGEMA_signal_1231, n2438}), .inb ({new_AGEMA_signal_1107, n2483}), .clk ( clk ), .rnd ({Fresh[761], Fresh[760]}), .outt ({new_AGEMA_signal_1417, n2439}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2598 ( .ina ({new_AGEMA_signal_1050, n2766}), .inb ({new_AGEMA_signal_1221, n2540}), .clk ( clk ), .rnd ({Fresh[763], Fresh[762]}), .outt ({new_AGEMA_signal_1418, n2445}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2600 ( .ina ({new_AGEMA_signal_1061, n2690}), .inb ({new_AGEMA_signal_1258, n2443}), .clk ( clk ), .rnd ({Fresh[765], Fresh[764]}), .outt ({new_AGEMA_signal_1419, n2444}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2602 ( .ina ({new_AGEMA_signal_959, n2790}), .inb ({new_AGEMA_signal_1208, n2446}), .clk ( clk ), .rnd ({Fresh[767], Fresh[766]}), .outt ({new_AGEMA_signal_1420, n2447}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2607 ( .ina ({new_AGEMA_signal_1144, n2761}), .inb ({new_AGEMA_signal_1259, n2693}), .clk ( clk ), .rnd ({Fresh[769], Fresh[768]}), .outt ({new_AGEMA_signal_1421, n2454}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2617 ( .ina ({new_AGEMA_signal_951, n2791}), .inb ({new_AGEMA_signal_1109, n2464}), .clk ( clk ), .rnd ({Fresh[771], Fresh[770]}), .outt ({new_AGEMA_signal_1260, n2465}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2622 ( .ina ({new_AGEMA_signal_953, n2813}), .inb ({new_AGEMA_signal_1087, n2576}), .clk ( clk ), .rnd ({Fresh[773], Fresh[772]}), .outt ({new_AGEMA_signal_1261, n2470}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2626 ( .ina ({new_AGEMA_signal_1111, n2473}), .inb ({new_AGEMA_signal_1112, n2472}), .clk ( clk ), .rnd ({Fresh[775], Fresh[774]}), .outt ({new_AGEMA_signal_1262, n2476}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2633 ( .ina ({new_AGEMA_signal_970, n2719}), .inb ({new_AGEMA_signal_1263, n2480}), .clk ( clk ), .rnd ({Fresh[777], Fresh[776]}), .outt ({new_AGEMA_signal_1424, n2481}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2639 ( .ina ({new_AGEMA_signal_1029, n2707}), .inb ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .rnd ({Fresh[779], Fresh[778]}), .outt ({new_AGEMA_signal_1265, n2486}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2642 ( .ina ({new_AGEMA_signal_991, n2661}), .inb ({new_AGEMA_signal_1114, n2488}), .clk ( clk ), .rnd ({Fresh[781], Fresh[780]}), .outt ({new_AGEMA_signal_1266, n2489}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2645 ( .ina ({new_AGEMA_signal_992, n2493}), .inb ({new_AGEMA_signal_1038, n2492}), .clk ( clk ), .rnd ({Fresh[783], Fresh[782]}), .outt ({new_AGEMA_signal_1267, n2497}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2646 ( .ina ({new_AGEMA_signal_1037, n2577}), .inb ({new_AGEMA_signal_1104, n2700}), .clk ( clk ), .rnd ({Fresh[785], Fresh[784]}), .outt ({new_AGEMA_signal_1268, n2495}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2647 ( .ina ({new_AGEMA_signal_976, n2780}), .inb ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .rnd ({Fresh[787], Fresh[786]}), .outt ({new_AGEMA_signal_1426, n2494}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2650 ( .ina ({new_AGEMA_signal_1077, n2498}), .inb ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[789], Fresh[788]}), .outt ({new_AGEMA_signal_1269, n2499}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2653 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .rnd ({Fresh[791], Fresh[790]}), .outt ({new_AGEMA_signal_1557, n2503}) ) ;
    mux2_HPC1 #(.security_order(1), .pipeline(0)) U2655 ( .ins ({new_AGEMA_signal_953, n2813}), .inb ({new_AGEMA_signal_1146, n2505}), .ina ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .rnd ({Fresh[793], Fresh[792]}), .outt ({new_AGEMA_signal_1427, n2506}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2662 ( .ina ({new_AGEMA_signal_1141, n2662}), .inb ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[795], Fresh[794]}), .outt ({new_AGEMA_signal_1428, n2518}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2663 ( .ina ({new_AGEMA_signal_1323, n2720}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[797], Fresh[796]}), .outt ({new_AGEMA_signal_1558, n2517}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2666 ( .ina ({new_AGEMA_signal_1270, n2520}), .inb ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .rnd ({Fresh[799], Fresh[798]}), .outt ({new_AGEMA_signal_1429, n2523}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2668 ( .ina ({new_AGEMA_signal_1228, n2774}), .inb ({new_AGEMA_signal_1115, n2521}), .clk ( clk ), .rnd ({Fresh[801], Fresh[800]}), .outt ({new_AGEMA_signal_1430, n2522}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2675 ( .ina ({SI_s1[1], SI_s0[1]}), .inb ({new_AGEMA_signal_1271, n2531}), .clk ( clk ), .rnd ({Fresh[803], Fresh[802]}), .outt ({new_AGEMA_signal_1431, n2532}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2677 ( .ina ({new_AGEMA_signal_1028, n2769}), .inb ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .rnd ({Fresh[805], Fresh[804]}), .outt ({new_AGEMA_signal_1432, n2534}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2681 ( .ina ({new_AGEMA_signal_1032, n2541}), .inb ({new_AGEMA_signal_1221, n2540}), .clk ( clk ), .rnd ({Fresh[807], Fresh[806]}), .outt ({new_AGEMA_signal_1433, n2542}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2683 ( .ina ({new_AGEMA_signal_1014, n2545}), .inb ({new_AGEMA_signal_1079, n2544}), .clk ( clk ), .rnd ({Fresh[809], Fresh[808]}), .outt ({new_AGEMA_signal_1272, n2546}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2687 ( .ina ({new_AGEMA_signal_1052, n2673}), .inb ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .rnd ({Fresh[811], Fresh[810]}), .outt ({new_AGEMA_signal_1435, n2551}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2690 ( .ina ({new_AGEMA_signal_1273, n2553}), .inb ({new_AGEMA_signal_1066, n2679}), .clk ( clk ), .rnd ({Fresh[813], Fresh[812]}), .outt ({new_AGEMA_signal_1436, n2558}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2692 ( .ina ({new_AGEMA_signal_1201, n2555}), .inb ({new_AGEMA_signal_1274, n2554}), .clk ( clk ), .rnd ({Fresh[815], Fresh[814]}), .outt ({new_AGEMA_signal_1437, n2556}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2696 ( .ina ({new_AGEMA_signal_1218, n2561}), .inb ({new_AGEMA_signal_1116, n2560}), .clk ( clk ), .rnd ({Fresh[817], Fresh[816]}), .outt ({new_AGEMA_signal_1438, n2566}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2697 ( .ina ({new_AGEMA_signal_974, n2699}), .inb ({new_AGEMA_signal_1186, n2562}), .clk ( clk ), .rnd ({Fresh[819], Fresh[818]}), .outt ({new_AGEMA_signal_1439, n2715}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2703 ( .ina ({new_AGEMA_signal_1160, n2572}), .inb ({new_AGEMA_signal_1055, n2571}), .clk ( clk ), .rnd ({Fresh[821], Fresh[820]}), .outt ({new_AGEMA_signal_1440, n2573}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2705 ( .ina ({new_AGEMA_signal_1026, n2767}), .inb ({new_AGEMA_signal_1173, n2754}), .clk ( clk ), .rnd ({Fresh[823], Fresh[822]}), .outt ({new_AGEMA_signal_1441, n2585}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2706 ( .ina ({new_AGEMA_signal_1027, n2789}), .inb ({new_AGEMA_signal_1048, n2627}), .clk ( clk ), .rnd ({Fresh[825], Fresh[824]}), .outt ({new_AGEMA_signal_1276, n2581}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2707 ( .ina ({new_AGEMA_signal_1127, n2575}), .inb ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .rnd ({Fresh[827], Fresh[826]}), .outt ({new_AGEMA_signal_1442, n2579}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2708 ( .ina ({new_AGEMA_signal_1037, n2577}), .inb ({new_AGEMA_signal_1087, n2576}), .clk ( clk ), .rnd ({Fresh[829], Fresh[828]}), .outt ({new_AGEMA_signal_1277, n2578}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2711 ( .ina ({new_AGEMA_signal_1148, n2625}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[831], Fresh[830]}), .outt ({new_AGEMA_signal_1443, n2582}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2715 ( .ina ({new_AGEMA_signal_993, n2587}), .inb ({new_AGEMA_signal_1278, n2586}), .clk ( clk ), .rnd ({Fresh[833], Fresh[832]}), .outt ({new_AGEMA_signal_1444, n2588}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2719 ( .ina ({new_AGEMA_signal_1105, n2594}), .inb ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .rnd ({Fresh[835], Fresh[834]}), .outt ({new_AGEMA_signal_1279, n2607}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2722 ( .ina ({new_AGEMA_signal_1117, n2597}), .inb ({new_AGEMA_signal_1280, n2596}), .clk ( clk ), .rnd ({Fresh[837], Fresh[836]}), .outt ({new_AGEMA_signal_1445, n2605}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2724 ( .ina ({new_AGEMA_signal_1281, n2598}), .inb ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .rnd ({Fresh[839], Fresh[838]}), .outt ({new_AGEMA_signal_1446, n2603}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2726 ( .ina ({new_AGEMA_signal_1021, n2599}), .inb ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .rnd ({Fresh[841], Fresh[840]}), .outt ({new_AGEMA_signal_1118, n2601}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2733 ( .ina ({new_AGEMA_signal_1283, n2610}), .inb ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .rnd ({Fresh[843], Fresh[842]}), .outt ({new_AGEMA_signal_1447, n2620}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2736 ( .ina ({new_AGEMA_signal_1284, n2614}), .inb ({new_AGEMA_signal_1285, n2613}), .clk ( clk ), .rnd ({Fresh[845], Fresh[844]}), .outt ({new_AGEMA_signal_1448, n2618}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2743 ( .ina ({new_AGEMA_signal_953, n2813}), .inb ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .rnd ({Fresh[847], Fresh[846]}), .outt ({new_AGEMA_signal_1449, n2626}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2746 ( .ina ({new_AGEMA_signal_1034, n2631}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[849], Fresh[848]}), .outt ({new_AGEMA_signal_1286, n2632}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2752 ( .ina ({new_AGEMA_signal_1287, n2784}), .inb ({new_AGEMA_signal_1074, n2642}), .clk ( clk ), .rnd ({Fresh[851], Fresh[850]}), .outt ({new_AGEMA_signal_1450, n2644}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2754 ( .ina ({SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1093, n2645}), .clk ( clk ), .rnd ({Fresh[853], Fresh[852]}), .outt ({new_AGEMA_signal_1288, n2646}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2758 ( .ina ({new_AGEMA_signal_1056, n2651}), .inb ({new_AGEMA_signal_1121, n2650}), .clk ( clk ), .rnd ({Fresh[855], Fresh[854]}), .outt ({new_AGEMA_signal_1289, n2653}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2760 ( .ina ({new_AGEMA_signal_1017, n2777}), .inb ({new_AGEMA_signal_1175, n2654}), .clk ( clk ), .rnd ({Fresh[857], Fresh[856]}), .outt ({new_AGEMA_signal_1452, n2655}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2764 ( .ina ({new_AGEMA_signal_1141, n2662}), .inb ({new_AGEMA_signal_991, n2661}), .clk ( clk ), .rnd ({Fresh[859], Fresh[858]}), .outt ({new_AGEMA_signal_1453, n2663}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2770 ( .ina ({new_AGEMA_signal_1052, n2673}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[861], Fresh[860]}), .outt ({new_AGEMA_signal_1290, n2675}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2772 ( .ina ({new_AGEMA_signal_1047, n2677}), .inb ({new_AGEMA_signal_1043, n2676}), .clk ( clk ), .rnd ({Fresh[863], Fresh[862]}), .outt ({new_AGEMA_signal_1291, n2678}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2780 ( .ina ({new_AGEMA_signal_1061, n2690}), .inb ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .rnd ({Fresh[865], Fresh[864]}), .outt ({new_AGEMA_signal_1292, n2691}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2782 ( .ina ({new_AGEMA_signal_978, n2694}), .inb ({new_AGEMA_signal_1259, n2693}), .clk ( clk ), .rnd ({Fresh[867], Fresh[866]}), .outt ({new_AGEMA_signal_1455, n2695}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2785 ( .ina ({new_AGEMA_signal_1104, n2700}), .inb ({new_AGEMA_signal_974, n2699}), .clk ( clk ), .rnd ({Fresh[869], Fresh[868]}), .outt ({new_AGEMA_signal_1293, n2701}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2791 ( .ina ({new_AGEMA_signal_1294, n2711}), .inb ({new_AGEMA_signal_1295, n2710}), .clk ( clk ), .rnd ({Fresh[871], Fresh[870]}), .outt ({new_AGEMA_signal_1456, n2717}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2796 ( .ina ({new_AGEMA_signal_1323, n2720}), .inb ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .rnd ({Fresh[873], Fresh[872]}), .outt ({new_AGEMA_signal_1576, n2729}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2798 ( .ina ({new_AGEMA_signal_981, n2723}), .inb ({new_AGEMA_signal_1123, n2722}), .clk ( clk ), .rnd ({Fresh[875], Fresh[874]}), .outt ({new_AGEMA_signal_1296, n2727}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2803 ( .ina ({new_AGEMA_signal_1135, n2732}), .inb ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .rnd ({Fresh[877], Fresh[876]}), .outt ({new_AGEMA_signal_1458, n2733}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2807 ( .ina ({new_AGEMA_signal_995, n2739}), .inb ({new_AGEMA_signal_1298, n2738}), .clk ( clk ), .rnd ({Fresh[879], Fresh[878]}), .outt ({new_AGEMA_signal_1459, n2740}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2812 ( .ina ({new_AGEMA_signal_1088, n2748}), .inb ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .rnd ({Fresh[881], Fresh[880]}), .outt ({new_AGEMA_signal_1299, n2749}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2815 ( .ina ({new_AGEMA_signal_1173, n2754}), .inb ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .rnd ({Fresh[883], Fresh[882]}), .outt ({new_AGEMA_signal_1461, n2757}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2816 ( .ina ({new_AGEMA_signal_1030, n2755}), .inb ({new_AGEMA_signal_1000, n2772}), .clk ( clk ), .rnd ({Fresh[885], Fresh[884]}), .outt ({new_AGEMA_signal_1300, n2756}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2819 ( .ina ({new_AGEMA_signal_1144, n2761}), .inb ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .rnd ({Fresh[887], Fresh[886]}), .outt ({new_AGEMA_signal_1462, n2762}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2823 ( .ina ({new_AGEMA_signal_1028, n2769}), .inb ({new_AGEMA_signal_1301, n2768}), .clk ( clk ), .rnd ({Fresh[889], Fresh[888]}), .outt ({new_AGEMA_signal_1463, n2770}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2825 ( .ina ({new_AGEMA_signal_1184, n2773}), .inb ({new_AGEMA_signal_1000, n2772}), .clk ( clk ), .rnd ({Fresh[891], Fresh[890]}), .outt ({new_AGEMA_signal_1464, n2776}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2826 ( .ina ({new_AGEMA_signal_1228, n2774}), .inb ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[893], Fresh[892]}), .outt ({new_AGEMA_signal_1465, n2775}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2830 ( .ina ({new_AGEMA_signal_1124, n2782}), .inb ({new_AGEMA_signal_1125, n2781}), .clk ( clk ), .rnd ({Fresh[895], Fresh[894]}), .outt ({new_AGEMA_signal_1302, n2783}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2836 ( .ina ({new_AGEMA_signal_1304, n2794}), .inb ({new_AGEMA_signal_1305, n2793}), .clk ( clk ), .rnd ({Fresh[897], Fresh[896]}), .outt ({new_AGEMA_signal_1467, n2795}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2845 ( .ina ({new_AGEMA_signal_1306, n2812}), .inb ({new_AGEMA_signal_1194, n2811}), .clk ( clk ), .rnd ({Fresh[899], Fresh[898]}), .outt ({new_AGEMA_signal_1468, n2814}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2848 ( .ina ({new_AGEMA_signal_1058, n2818}), .inb ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .rnd ({Fresh[901], Fresh[900]}), .outt ({new_AGEMA_signal_1307, n2819}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1968 ( .ina ({new_AGEMA_signal_1309, n1924}), .inb ({new_AGEMA_signal_1310, n1923}), .clk ( clk ), .rnd ({Fresh[903], Fresh[902]}), .outt ({new_AGEMA_signal_1470, n1936}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1982 ( .ina ({new_AGEMA_signal_1030, n2755}), .inb ({new_AGEMA_signal_1311, n1927}), .clk ( clk ), .rnd ({Fresh[905], Fresh[904]}), .outt ({new_AGEMA_signal_1471, n1928}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U1994 ( .ina ({new_AGEMA_signal_1132, n2151}), .inb ({new_AGEMA_signal_1312, n1929}), .clk ( clk ), .rnd ({Fresh[907], Fresh[906]}), .outt ({new_AGEMA_signal_1472, n1931}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2012 ( .ina ({new_AGEMA_signal_1313, n2665}), .inb ({new_AGEMA_signal_1314, n1938}), .clk ( clk ), .rnd ({Fresh[909], Fresh[908]}), .outt ({new_AGEMA_signal_1473, n1939}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2024 ( .ina ({new_AGEMA_signal_1315, n2235}), .inb ({new_AGEMA_signal_1137, n1943}), .clk ( clk ), .rnd ({Fresh[911], Fresh[910]}), .outt ({new_AGEMA_signal_1474, n1948}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2032 ( .ina ({new_AGEMA_signal_1138, n1946}), .inb ({new_AGEMA_signal_1316, n1945}), .clk ( clk ), .rnd ({Fresh[913], Fresh[912]}), .outt ({new_AGEMA_signal_1475, n1947}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2041 ( .ina ({new_AGEMA_signal_1045, n2442}), .inb ({new_AGEMA_signal_1318, n1951}), .clk ( clk ), .rnd ({Fresh[915], Fresh[914]}), .outt ({new_AGEMA_signal_1476, n1954}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2049 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1319, n1952}), .clk ( clk ), .rnd ({Fresh[917], Fresh[916]}), .outt ({new_AGEMA_signal_1477, n1953}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2058 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1320, n2687}), .clk ( clk ), .rnd ({Fresh[919], Fresh[918]}), .outt ({new_AGEMA_signal_1478, n2658}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2065 ( .ina ({new_AGEMA_signal_999, n1964}), .inb ({new_AGEMA_signal_1143, n1963}), .clk ( clk ), .rnd ({Fresh[921], Fresh[920]}), .outt ({new_AGEMA_signal_1322, n1965}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2078 ( .ina ({new_AGEMA_signal_1052, n2673}), .inb ({new_AGEMA_signal_1480, n1968}), .clk ( clk ), .rnd ({Fresh[923], Fresh[922]}), .outt ({new_AGEMA_signal_1591, n1970}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2084 ( .ina ({new_AGEMA_signal_1325, n2684}), .inb ({new_AGEMA_signal_1147, n2359}), .clk ( clk ), .rnd ({Fresh[925], Fresh[924]}), .outt ({new_AGEMA_signal_1481, n1969}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2093 ( .ina ({new_AGEMA_signal_1326, n1972}), .inb ({new_AGEMA_signal_1149, n1971}), .clk ( clk ), .rnd ({Fresh[927], Fresh[926]}), .outt ({new_AGEMA_signal_1482, n1978}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2102 ( .ina ({new_AGEMA_signal_1327, n1974}), .inb ({new_AGEMA_signal_1151, n1973}), .clk ( clk ), .rnd ({Fresh[929], Fresh[928]}), .outt ({new_AGEMA_signal_1483, n1975}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2107 ( .ina ({new_AGEMA_signal_1061, n2690}), .inb ({new_AGEMA_signal_1328, n1979}), .clk ( clk ), .rnd ({Fresh[931], Fresh[930]}), .outt ({new_AGEMA_signal_1484, n1980}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2114 ( .ina ({new_AGEMA_signal_1152, n1985}), .inb ({new_AGEMA_signal_1153, n2741}), .clk ( clk ), .rnd ({Fresh[933], Fresh[932]}), .outt ({new_AGEMA_signal_1329, n1986}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2124 ( .ina ({new_AGEMA_signal_1330, n1994}), .inb ({new_AGEMA_signal_1064, n1993}), .clk ( clk ), .rnd ({Fresh[935], Fresh[934]}), .outt ({new_AGEMA_signal_1486, n1997}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2137 ( .ina ({new_AGEMA_signal_1157, n2241}), .inb ({new_AGEMA_signal_1332, n2137}), .clk ( clk ), .rnd ({Fresh[937], Fresh[936]}), .outt ({new_AGEMA_signal_1487, n2012}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2145 ( .ina ({new_AGEMA_signal_1333, n2006}), .inb ({new_AGEMA_signal_1334, n2005}), .clk ( clk ), .rnd ({Fresh[939], Fresh[938]}), .outt ({new_AGEMA_signal_1488, n2007}) ) ;
    mux2_HPC1 #(.security_order(1), .pipeline(0)) U2161 ( .ins ({new_AGEMA_signal_953, n2813}), .inb ({new_AGEMA_signal_1165, n2020}), .ina ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .rnd ({Fresh[941], Fresh[940]}), .outt ({new_AGEMA_signal_1336, n2021}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2176 ( .ina ({new_AGEMA_signal_1168, n2290}), .inb ({new_AGEMA_signal_1338, n2031}), .clk ( clk ), .rnd ({Fresh[943], Fresh[942]}), .outt ({new_AGEMA_signal_1490, n2032}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2185 ( .ina ({new_AGEMA_signal_1073, n2171}), .inb ({new_AGEMA_signal_1339, n2040}), .clk ( clk ), .rnd ({Fresh[945], Fresh[944]}), .outt ({new_AGEMA_signal_1491, n2041}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2189 ( .ina ({new_AGEMA_signal_1313, n2665}), .inb ({new_AGEMA_signal_1172, n2042}), .clk ( clk ), .rnd ({Fresh[947], Fresh[946]}), .outt ({new_AGEMA_signal_1492, n2043}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2194 ( .ina ({new_AGEMA_signal_1173, n2754}), .inb ({new_AGEMA_signal_1340, n2045}), .clk ( clk ), .rnd ({Fresh[949], Fresh[948]}), .outt ({new_AGEMA_signal_1493, n2046}) ) ;
    mux2_HPC1 #(.security_order(1), .pipeline(0)) U2204 ( .ins ({new_AGEMA_signal_953, n2813}), .inb ({new_AGEMA_signal_1342, n2056}), .ina ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .rnd ({Fresh[951], Fresh[950]}), .outt ({new_AGEMA_signal_1494, n2058}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2210 ( .ina ({new_AGEMA_signal_1150, n2535}), .inb ({new_AGEMA_signal_1343, n2060}), .clk ( clk ), .rnd ({Fresh[953], Fresh[952]}), .outt ({new_AGEMA_signal_1495, n2063}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2218 ( .ina ({new_AGEMA_signal_1344, n2066}), .inb ({new_AGEMA_signal_1345, n2065}), .clk ( clk ), .rnd ({Fresh[955], Fresh[954]}), .outt ({new_AGEMA_signal_1496, n2652}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2227 ( .ina ({new_AGEMA_signal_1074, n2642}), .inb ({new_AGEMA_signal_1347, n2074}), .clk ( clk ), .rnd ({Fresh[957], Fresh[956]}), .outt ({new_AGEMA_signal_1497, n2076}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2236 ( .ina ({new_AGEMA_signal_1011, n2721}), .inb ({new_AGEMA_signal_1348, n2082}), .clk ( clk ), .rnd ({Fresh[959], Fresh[958]}), .outt ({new_AGEMA_signal_1498, n2105}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2241 ( .ina ({new_AGEMA_signal_1184, n2773}), .inb ({new_AGEMA_signal_1349, n2084}), .clk ( clk ), .rnd ({Fresh[961], Fresh[960]}), .outt ({new_AGEMA_signal_1499, n2099}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2243 ( .ina ({new_AGEMA_signal_1350, n2085}), .inb ({new_AGEMA_signal_1048, n2627}), .clk ( clk ), .rnd ({Fresh[963], Fresh[962]}), .outt ({new_AGEMA_signal_1500, n2091}) ) ;
    and_HPC1 #(.security_order(1), .pipeline(0)) U2246 ( .ina ({new_AGEMA_signal_987, n2753}), .inb ({new_AGEMA_signal_1351, n2131}), .clk ( clk ), .rnd ({Fresh[965], Fresh[964]}), .outt ({new_AGEMA_signal_1501, n2090}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2253 ( .ina ({new_AGEMA_signal_1034, n2631}), .inb ({new_AGEMA_signal_1353, n2330}), .clk ( clk ), .rnd ({Fresh[967], Fresh[966]}), .outt ({new_AGEMA_signal_1502, n2093}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2262 ( .ina ({new_AGEMA_signal_1169, n2376}), .inb ({new_AGEMA_signal_1356, n2160}), .clk ( clk ), .rnd ({Fresh[969], Fresh[968]}), .outt ({new_AGEMA_signal_1503, n2102}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2266 ( .ina ({new_AGEMA_signal_1189, n2504}), .inb ({new_AGEMA_signal_1063, n2823}), .clk ( clk ), .rnd ({Fresh[971], Fresh[970]}), .outt ({new_AGEMA_signal_1357, n2106}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2272 ( .ina ({new_AGEMA_signal_980, n2713}), .inb ({new_AGEMA_signal_1504, n2114}), .clk ( clk ), .rnd ({Fresh[973], Fresh[972]}), .outt ({new_AGEMA_signal_1606, n2116}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2282 ( .ina ({new_AGEMA_signal_1358, n2291}), .inb ({new_AGEMA_signal_1192, n2119}), .clk ( clk ), .rnd ({Fresh[975], Fresh[974]}), .outt ({new_AGEMA_signal_1505, n2120}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2293 ( .ina ({new_AGEMA_signal_1195, n2130}), .inb ({new_AGEMA_signal_1196, n2129}), .clk ( clk ), .rnd ({Fresh[977], Fresh[976]}), .outt ({new_AGEMA_signal_1359, n2155}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2296 ( .ina ({new_AGEMA_signal_994, n2643}), .inb ({new_AGEMA_signal_1351, n2131}), .clk ( clk ), .rnd ({Fresh[979], Fresh[978]}), .outt ({new_AGEMA_signal_1506, n2543}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2299 ( .ina ({new_AGEMA_signal_1198, n2133}), .inb ({new_AGEMA_signal_975, n2816}), .clk ( clk ), .rnd ({Fresh[981], Fresh[980]}), .outt ({new_AGEMA_signal_1360, n2134}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2303 ( .ina ({new_AGEMA_signal_1332, n2137}), .inb ({new_AGEMA_signal_1361, n2136}), .clk ( clk ), .rnd ({Fresh[983], Fresh[982]}), .outt ({new_AGEMA_signal_1508, n2143}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2308 ( .ina ({new_AGEMA_signal_1362, n2139}), .inb ({new_AGEMA_signal_1013, n2346}), .clk ( clk ), .rnd ({Fresh[985], Fresh[984]}), .outt ({new_AGEMA_signal_1509, n2140}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2324 ( .ina ({new_AGEMA_signal_1366, n2157}), .inb ({new_AGEMA_signal_1066, n2679}), .clk ( clk ), .rnd ({Fresh[987], Fresh[986]}), .outt ({new_AGEMA_signal_1510, n2159}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2326 ( .ina ({new_AGEMA_signal_1356, n2160}), .inb ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .rnd ({Fresh[989], Fresh[988]}), .outt ({new_AGEMA_signal_1511, n2161}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2330 ( .ina ({new_AGEMA_signal_1045, n2442}), .inb ({new_AGEMA_signal_1203, n2163}), .clk ( clk ), .rnd ({Fresh[991], Fresh[990]}), .outt ({new_AGEMA_signal_1367, n2164}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2345 ( .ina ({new_AGEMA_signal_1085, n2178}), .inb ({new_AGEMA_signal_1370, n2177}), .clk ( clk ), .rnd ({Fresh[993], Fresh[992]}), .outt ({new_AGEMA_signal_1513, n2179}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2359 ( .ina ({new_AGEMA_signal_961, n2315}), .inb ({new_AGEMA_signal_1373, n2191}), .clk ( clk ), .rnd ({Fresh[995], Fresh[994]}), .outt ({new_AGEMA_signal_1514, n2192}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2370 ( .ina ({new_AGEMA_signal_1374, n2201}), .inb ({new_AGEMA_signal_1515, n2200}), .clk ( clk ), .rnd ({Fresh[997], Fresh[996]}), .outt ({new_AGEMA_signal_1613, n2203}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2382 ( .ina ({new_AGEMA_signal_1376, n2217}), .inb ({new_AGEMA_signal_1210, n2216}), .clk ( clk ), .rnd ({Fresh[999], Fresh[998]}), .outt ({new_AGEMA_signal_1517, n2224}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2388 ( .ina ({new_AGEMA_signal_1377, n2222}), .inb ({new_AGEMA_signal_1378, n2221}), .clk ( clk ), .rnd ({Fresh[1001], Fresh[1000]}), .outt ({new_AGEMA_signal_1518, n2223}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2392 ( .ina ({new_AGEMA_signal_1189, n2504}), .inb ({new_AGEMA_signal_1213, n2226}), .clk ( clk ), .rnd ({Fresh[1003], Fresh[1002]}), .outt ({new_AGEMA_signal_1379, n2229}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2399 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1520, n2233}), .clk ( clk ), .rnd ({Fresh[1005], Fresh[1004]}), .outt ({new_AGEMA_signal_1616, n2234}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2410 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1381, n2244}), .clk ( clk ), .rnd ({Fresh[1007], Fresh[1006]}), .outt ({new_AGEMA_signal_1521, n2246}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2418 ( .ina ({new_AGEMA_signal_1146, n2505}), .inb ({new_AGEMA_signal_1383, n2253}), .clk ( clk ), .rnd ({Fresh[1009], Fresh[1008]}), .outt ({new_AGEMA_signal_1522, n2254}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2425 ( .ina ({new_AGEMA_signal_1221, n2540}), .inb ({new_AGEMA_signal_1384, n2260}), .clk ( clk ), .rnd ({Fresh[1011], Fresh[1010]}), .outt ({new_AGEMA_signal_1523, n2263}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2434 ( .ina ({new_AGEMA_signal_1092, n2266}), .inb ({new_AGEMA_signal_1223, n2265}), .clk ( clk ), .rnd ({Fresh[1013], Fresh[1012]}), .outt ({new_AGEMA_signal_1385, n2267}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2438 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1224, n2269}), .clk ( clk ), .rnd ({Fresh[1015], Fresh[1014]}), .outt ({new_AGEMA_signal_1386, n2270}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2445 ( .ina ({new_AGEMA_signal_1225, n2278}), .inb ({new_AGEMA_signal_1226, n2277}), .clk ( clk ), .rnd ({Fresh[1017], Fresh[1016]}), .outt ({new_AGEMA_signal_1387, n2279}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2450 ( .ina ({new_AGEMA_signal_967, n2779}), .inb ({new_AGEMA_signal_1227, n2282}), .clk ( clk ), .rnd ({Fresh[1019], Fresh[1018]}), .outt ({new_AGEMA_signal_1388, n2283}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2453 ( .ina ({new_AGEMA_signal_1184, n2773}), .inb ({new_AGEMA_signal_1389, n2284}), .clk ( clk ), .rnd ({Fresh[1021], Fresh[1020]}), .outt ({new_AGEMA_signal_1528, n2285}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2457 ( .ina ({new_AGEMA_signal_1045, n2442}), .inb ({new_AGEMA_signal_1390, n2459}), .clk ( clk ), .rnd ({Fresh[1023], Fresh[1022]}), .outt ({new_AGEMA_signal_1529, n2686}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2460 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1391, n2288}), .clk ( clk ), .rnd ({Fresh[1025], Fresh[1024]}), .outt ({new_AGEMA_signal_1530, n2289}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2463 ( .ina ({new_AGEMA_signal_1392, n2458}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[1027], Fresh[1026]}), .outt ({new_AGEMA_signal_1531, n2297}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2465 ( .ina ({new_AGEMA_signal_1003, n2624}), .inb ({new_AGEMA_signal_1358, n2291}), .clk ( clk ), .rnd ({Fresh[1029], Fresh[1028]}), .outt ({new_AGEMA_signal_1532, n2292}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2473 ( .ina ({new_AGEMA_signal_981, n2723}), .inb ({new_AGEMA_signal_1394, n2300}), .clk ( clk ), .rnd ({Fresh[1031], Fresh[1030]}), .outt ({new_AGEMA_signal_1533, n2301}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2483 ( .ina ({SI_s1[1], SI_s0[1]}), .inb ({new_AGEMA_signal_1396, n2314}), .clk ( clk ), .rnd ({Fresh[1033], Fresh[1032]}), .outt ({new_AGEMA_signal_1534, n2321}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2487 ( .ina ({new_AGEMA_signal_1097, n2319}), .inb ({new_AGEMA_signal_1098, n2318}), .clk ( clk ), .rnd ({Fresh[1035], Fresh[1034]}), .outt ({new_AGEMA_signal_1233, n2320}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2493 ( .ina ({new_AGEMA_signal_1234, n2326}), .inb ({new_AGEMA_signal_1235, n2325}), .clk ( clk ), .rnd ({Fresh[1037], Fresh[1036]}), .outt ({new_AGEMA_signal_1397, n2334}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2497 ( .ina ({new_AGEMA_signal_1398, n2329}), .inb ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .rnd ({Fresh[1039], Fresh[1038]}), .outt ({new_AGEMA_signal_1535, n2332}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2498 ( .ina ({new_AGEMA_signal_1047, n2677}), .inb ({new_AGEMA_signal_1353, n2330}), .clk ( clk ), .rnd ({Fresh[1041], Fresh[1040]}), .outt ({new_AGEMA_signal_1536, n2331}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2502 ( .ina ({new_AGEMA_signal_1037, n2577}), .inb ({new_AGEMA_signal_1537, n2335}), .clk ( clk ), .rnd ({Fresh[1043], Fresh[1042]}), .outt ({new_AGEMA_signal_1626, n2336}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2508 ( .ina ({new_AGEMA_signal_1399, n2341}), .inb ({new_AGEMA_signal_1238, n2340}), .clk ( clk ), .rnd ({Fresh[1045], Fresh[1044]}), .outt ({new_AGEMA_signal_1538, n2342}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2519 ( .ina ({new_AGEMA_signal_1242, n2352}), .inb ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .rnd ({Fresh[1047], Fresh[1046]}), .outt ({new_AGEMA_signal_1400, n2367}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2523 ( .ina ({new_AGEMA_signal_1401, n2354}), .inb ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .rnd ({Fresh[1049], Fresh[1048]}), .outt ({new_AGEMA_signal_1539, n2358}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2547 ( .ina ({new_AGEMA_signal_1247, n2385}), .inb ({new_AGEMA_signal_1248, n2384}), .clk ( clk ), .rnd ({Fresh[1051], Fresh[1050]}), .outt ({new_AGEMA_signal_1406, n2387}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2555 ( .ina ({new_AGEMA_signal_1250, n2391}), .inb ({new_AGEMA_signal_1408, n2390}), .clk ( clk ), .rnd ({Fresh[1053], Fresh[1052]}), .outt ({new_AGEMA_signal_1542, n2392}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2566 ( .ina ({new_AGEMA_signal_1252, n2403}), .inb ({SI_s1[6], SI_s0[6]}), .clk ( clk ), .rnd ({Fresh[1055], Fresh[1054]}), .outt ({new_AGEMA_signal_1410, n2404}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2570 ( .ina ({new_AGEMA_signal_1150, n2535}), .inb ({new_AGEMA_signal_1411, n2408}), .clk ( clk ), .rnd ({Fresh[1057], Fresh[1056]}), .outt ({new_AGEMA_signal_1544, n2409}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2575 ( .ina ({new_AGEMA_signal_1412, n2574}), .inb ({new_AGEMA_signal_1253, n2413}), .clk ( clk ), .rnd ({Fresh[1059], Fresh[1058]}), .outt ({new_AGEMA_signal_1545, n2414}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2578 ( .ina ({new_AGEMA_signal_1148, n2625}), .inb ({new_AGEMA_signal_1254, n2416}), .clk ( clk ), .rnd ({Fresh[1061], Fresh[1060]}), .outt ({new_AGEMA_signal_1413, n2418}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2589 ( .ina ({new_AGEMA_signal_1415, n2689}), .inb ({new_AGEMA_signal_1256, n2431}), .clk ( clk ), .rnd ({Fresh[1063], Fresh[1062]}), .outt ({new_AGEMA_signal_1547, n2432}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2592 ( .ina ({SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_1257, n2434}), .clk ( clk ), .rnd ({Fresh[1065], Fresh[1064]}), .outt ({new_AGEMA_signal_1416, n2435}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2601 ( .ina ({new_AGEMA_signal_1418, n2445}), .inb ({new_AGEMA_signal_1419, n2444}), .clk ( clk ), .rnd ({Fresh[1067], Fresh[1066]}), .outt ({new_AGEMA_signal_1548, n2449}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2603 ( .ina ({SI_s1[1], SI_s0[1]}), .inb ({new_AGEMA_signal_1420, n2447}), .clk ( clk ), .rnd ({Fresh[1069], Fresh[1068]}), .outt ({new_AGEMA_signal_1549, n2448}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2609 ( .ina ({new_AGEMA_signal_1421, n2454}), .inb ({new_AGEMA_signal_1108, n2453}), .clk ( clk ), .rnd ({Fresh[1071], Fresh[1070]}), .outt ({new_AGEMA_signal_1550, n2455}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2612 ( .ina ({new_AGEMA_signal_1320, n2687}), .inb ({new_AGEMA_signal_1392, n2458}), .clk ( clk ), .rnd ({Fresh[1073], Fresh[1072]}), .outt ({new_AGEMA_signal_1551, n2460}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2618 ( .ina ({new_AGEMA_signal_1003, n2624}), .inb ({new_AGEMA_signal_1260, n2465}), .clk ( clk ), .rnd ({Fresh[1075], Fresh[1074]}), .outt ({new_AGEMA_signal_1422, n2466}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2629 ( .ina ({new_AGEMA_signal_1262, n2476}), .inb ({new_AGEMA_signal_1113, n2475}), .clk ( clk ), .rnd ({Fresh[1077], Fresh[1076]}), .outt ({new_AGEMA_signal_1423, n2477}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2634 ( .ina ({new_AGEMA_signal_1028, n2769}), .inb ({new_AGEMA_signal_1424, n2481}), .clk ( clk ), .rnd ({Fresh[1079], Fresh[1078]}), .outt ({new_AGEMA_signal_1554, n2482}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2640 ( .ina ({new_AGEMA_signal_1264, n2487}), .inb ({new_AGEMA_signal_1265, n2486}), .clk ( clk ), .rnd ({Fresh[1081], Fresh[1080]}), .outt ({new_AGEMA_signal_1425, n2490}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2648 ( .ina ({new_AGEMA_signal_1268, n2495}), .inb ({new_AGEMA_signal_1426, n2494}), .clk ( clk ), .rnd ({Fresh[1083], Fresh[1082]}), .outt ({new_AGEMA_signal_1556, n2496}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2654 ( .ina ({new_AGEMA_signal_1189, n2504}), .inb ({new_AGEMA_signal_1557, n2503}), .clk ( clk ), .rnd ({Fresh[1085], Fresh[1084]}), .outt ({new_AGEMA_signal_1643, n2507}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2664 ( .ina ({new_AGEMA_signal_1428, n2518}), .inb ({new_AGEMA_signal_1558, n2517}), .clk ( clk ), .rnd ({Fresh[1087], Fresh[1086]}), .outt ({new_AGEMA_signal_1644, n2525}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2669 ( .ina ({new_AGEMA_signal_1429, n2523}), .inb ({new_AGEMA_signal_1430, n2522}), .clk ( clk ), .rnd ({Fresh[1089], Fresh[1088]}), .outt ({new_AGEMA_signal_1559, n2524}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2676 ( .ina ({new_AGEMA_signal_1431, n2532}), .inb ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[1091], Fresh[1090]}), .outt ({new_AGEMA_signal_1560, n2537}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2678 ( .ina ({new_AGEMA_signal_1150, n2535}), .inb ({new_AGEMA_signal_1432, n2534}), .clk ( clk ), .rnd ({Fresh[1093], Fresh[1092]}), .outt ({new_AGEMA_signal_1561, n2536}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2684 ( .ina ({new_AGEMA_signal_1040, n2724}), .inb ({new_AGEMA_signal_1272, n2546}), .clk ( clk ), .rnd ({Fresh[1095], Fresh[1094]}), .outt ({new_AGEMA_signal_1434, n2547}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2693 ( .ina ({new_AGEMA_signal_1031, n2688}), .inb ({new_AGEMA_signal_1437, n2556}), .clk ( clk ), .rnd ({Fresh[1097], Fresh[1096]}), .outt ({new_AGEMA_signal_1562, n2557}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2699 ( .ina ({new_AGEMA_signal_1439, n2715}), .inb ({new_AGEMA_signal_1275, n2564}), .clk ( clk ), .rnd ({Fresh[1099], Fresh[1098]}), .outt ({new_AGEMA_signal_1563, n2565}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2704 ( .ina ({new_AGEMA_signal_1412, n2574}), .inb ({new_AGEMA_signal_1440, n2573}), .clk ( clk ), .rnd ({Fresh[1101], Fresh[1100]}), .outt ({new_AGEMA_signal_1564, n2591}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2709 ( .ina ({new_AGEMA_signal_1442, n2579}), .inb ({new_AGEMA_signal_1277, n2578}), .clk ( clk ), .rnd ({Fresh[1103], Fresh[1102]}), .outt ({new_AGEMA_signal_1565, n2580}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2727 ( .ina ({new_AGEMA_signal_1118, n2601}), .inb ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .rnd ({Fresh[1105], Fresh[1104]}), .outt ({new_AGEMA_signal_1282, n2602}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2738 ( .ina ({new_AGEMA_signal_1448, n2618}), .inb ({new_AGEMA_signal_1119, n2617}), .clk ( clk ), .rnd ({Fresh[1107], Fresh[1106]}), .outt ({new_AGEMA_signal_1567, n2619}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2744 ( .ina ({new_AGEMA_signal_1048, n2627}), .inb ({new_AGEMA_signal_1449, n2626}), .clk ( clk ), .rnd ({Fresh[1109], Fresh[1108]}), .outt ({new_AGEMA_signal_1568, n2628}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2753 ( .ina ({new_AGEMA_signal_1450, n2644}), .inb ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .rnd ({Fresh[1111], Fresh[1110]}), .outt ({new_AGEMA_signal_1569, n2649}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2755 ( .ina ({new_AGEMA_signal_1081, n2647}), .inb ({new_AGEMA_signal_1288, n2646}), .clk ( clk ), .rnd ({Fresh[1113], Fresh[1112]}), .outt ({new_AGEMA_signal_1451, n2648}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2765 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1453, n2663}), .clk ( clk ), .rnd ({Fresh[1115], Fresh[1114]}), .outt ({new_AGEMA_signal_1570, n2664}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2771 ( .ina ({new_AGEMA_signal_1290, n2675}), .inb ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .rnd ({Fresh[1117], Fresh[1116]}), .outt ({new_AGEMA_signal_1571, n2681}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2773 ( .ina ({new_AGEMA_signal_1066, n2679}), .inb ({new_AGEMA_signal_1291, n2678}), .clk ( clk ), .rnd ({Fresh[1119], Fresh[1118]}), .outt ({new_AGEMA_signal_1454, n2680}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2776 ( .ina ({new_AGEMA_signal_1325, n2684}), .inb ({new_AGEMA_signal_1022, n2683}), .clk ( clk ), .rnd ({Fresh[1121], Fresh[1120]}), .outt ({new_AGEMA_signal_1572, n2685}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2778 ( .ina ({new_AGEMA_signal_1320, n2687}), .inb ({new_AGEMA_signal_1040, n2724}), .clk ( clk ), .rnd ({Fresh[1123], Fresh[1122]}), .outt ({new_AGEMA_signal_1573, n2698}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2779 ( .ina ({new_AGEMA_signal_1415, n2689}), .inb ({new_AGEMA_signal_1031, n2688}), .clk ( clk ), .rnd ({Fresh[1125], Fresh[1124]}), .outt ({new_AGEMA_signal_1574, n2692}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2793 ( .ina ({new_AGEMA_signal_1439, n2715}), .inb ({new_AGEMA_signal_1122, n2714}), .clk ( clk ), .rnd ({Fresh[1127], Fresh[1126]}), .outt ({new_AGEMA_signal_1575, n2716}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2800 ( .ina ({new_AGEMA_signal_1296, n2727}), .inb ({new_AGEMA_signal_1297, n2726}), .clk ( clk ), .rnd ({Fresh[1129], Fresh[1128]}), .outt ({new_AGEMA_signal_1457, n2728}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2804 ( .ina ({new_AGEMA_signal_1133, n2734}), .inb ({new_AGEMA_signal_1458, n2733}), .clk ( clk ), .rnd ({Fresh[1131], Fresh[1130]}), .outt ({new_AGEMA_signal_1577, n2735}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2808 ( .ina ({new_AGEMA_signal_1153, n2741}), .inb ({new_AGEMA_signal_1459, n2740}), .clk ( clk ), .rnd ({Fresh[1133], Fresh[1132]}), .outt ({new_AGEMA_signal_1578, n2743}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2813 ( .ina ({new_AGEMA_signal_972, n2750}), .inb ({new_AGEMA_signal_1299, n2749}), .clk ( clk ), .rnd ({Fresh[1135], Fresh[1134]}), .outt ({new_AGEMA_signal_1460, n2751}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2817 ( .ina ({new_AGEMA_signal_1461, n2757}), .inb ({new_AGEMA_signal_1300, n2756}), .clk ( clk ), .rnd ({Fresh[1137], Fresh[1136]}), .outt ({new_AGEMA_signal_1579, n2758}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2820 ( .ina ({new_AGEMA_signal_1134, n2763}), .inb ({new_AGEMA_signal_1462, n2762}), .clk ( clk ), .rnd ({Fresh[1139], Fresh[1138]}), .outt ({new_AGEMA_signal_1580, n2764}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2827 ( .ina ({new_AGEMA_signal_1464, n2776}), .inb ({new_AGEMA_signal_1465, n2775}), .clk ( clk ), .rnd ({Fresh[1141], Fresh[1140]}), .outt ({new_AGEMA_signal_1581, n2800}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2831 ( .ina ({new_AGEMA_signal_1287, n2784}), .inb ({new_AGEMA_signal_1302, n2783}), .clk ( clk ), .rnd ({Fresh[1143], Fresh[1142]}), .outt ({new_AGEMA_signal_1466, n2788}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2837 ( .ina ({new_AGEMA_signal_943, n2796}), .inb ({new_AGEMA_signal_1467, n2795}), .clk ( clk ), .rnd ({Fresh[1145], Fresh[1144]}), .outt ({new_AGEMA_signal_1583, n2797}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2846 ( .ina ({new_AGEMA_signal_1468, n2814}), .inb ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .rnd ({Fresh[1147], Fresh[1146]}), .outt ({new_AGEMA_signal_1584, n2822}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2849 ( .ina ({new_AGEMA_signal_1126, n2820}), .inb ({new_AGEMA_signal_1307, n2819}), .clk ( clk ), .rnd ({Fresh[1149], Fresh[1148]}), .outt ({new_AGEMA_signal_1469, n2821}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1983 ( .ina ({new_AGEMA_signal_1029, n2707}), .inb ({new_AGEMA_signal_1471, n1928}), .clk ( clk ), .rnd ({Fresh[1151], Fresh[1150]}), .outt ({new_AGEMA_signal_1585, n1934}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U1998 ( .ina ({new_AGEMA_signal_1472, n1931}), .inb ({new_AGEMA_signal_1036, n1930}), .clk ( clk ), .rnd ({Fresh[1153], Fresh[1152]}), .outt ({new_AGEMA_signal_1586, n1932}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2015 ( .ina ({new_AGEMA_signal_1473, n1939}), .inb ({new_AGEMA_signal_1040, n2724}), .clk ( clk ), .rnd ({Fresh[1155], Fresh[1154]}), .outt ({new_AGEMA_signal_1587, n1940}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2033 ( .ina ({new_AGEMA_signal_1474, n1948}), .inb ({new_AGEMA_signal_1475, n1947}), .clk ( clk ), .rnd ({Fresh[1157], Fresh[1156]}), .outt ({new_AGEMA_signal_1588, n1961}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2050 ( .ina ({new_AGEMA_signal_1476, n1954}), .inb ({new_AGEMA_signal_1477, n1953}), .clk ( clk ), .rnd ({Fresh[1159], Fresh[1158]}), .outt ({new_AGEMA_signal_1589, n1955}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2066 ( .ina ({new_AGEMA_signal_1321, n1966}), .inb ({new_AGEMA_signal_1322, n1965}), .clk ( clk ), .rnd ({Fresh[1161], Fresh[1160]}), .outt ({new_AGEMA_signal_1479, n1967}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2085 ( .ina ({new_AGEMA_signal_1591, n1970}), .inb ({new_AGEMA_signal_1481, n1969}), .clk ( clk ), .rnd ({Fresh[1163], Fresh[1162]}), .outt ({new_AGEMA_signal_1669, n1984}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2103 ( .ina ({new_AGEMA_signal_1060, n1976}), .inb ({new_AGEMA_signal_1483, n1975}), .clk ( clk ), .rnd ({Fresh[1165], Fresh[1164]}), .outt ({new_AGEMA_signal_1592, n1977}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2108 ( .ina ({SI_s1[1], SI_s0[1]}), .inb ({new_AGEMA_signal_1484, n1980}), .clk ( clk ), .rnd ({Fresh[1167], Fresh[1166]}), .outt ({new_AGEMA_signal_1593, n1981}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2115 ( .ina ({new_AGEMA_signal_983, n2815}), .inb ({new_AGEMA_signal_1329, n1986}), .clk ( clk ), .rnd ({Fresh[1169], Fresh[1168]}), .outt ({new_AGEMA_signal_1485, n1987}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2127 ( .ina ({new_AGEMA_signal_1486, n1997}), .inb ({new_AGEMA_signal_1331, n1996}), .clk ( clk ), .rnd ({Fresh[1171], Fresh[1170]}), .outt ({new_AGEMA_signal_1594, n1998}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2146 ( .ina ({new_AGEMA_signal_1159, n2008}), .inb ({new_AGEMA_signal_1488, n2007}), .clk ( clk ), .rnd ({Fresh[1173], Fresh[1172]}), .outt ({new_AGEMA_signal_1595, n2010}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2162 ( .ina ({new_AGEMA_signal_1164, n2022}), .inb ({new_AGEMA_signal_1336, n2021}), .clk ( clk ), .rnd ({Fresh[1175], Fresh[1174]}), .outt ({new_AGEMA_signal_1489, n2024}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2177 ( .ina ({new_AGEMA_signal_1337, n2033}), .inb ({new_AGEMA_signal_1490, n2032}), .clk ( clk ), .rnd ({Fresh[1177], Fresh[1176]}), .outt ({new_AGEMA_signal_1597, n2035}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2186 ( .ina ({new_AGEMA_signal_1491, n2041}), .inb ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .rnd ({Fresh[1179], Fresh[1178]}), .outt ({new_AGEMA_signal_1598, n2054}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2190 ( .ina ({new_AGEMA_signal_980, n2713}), .inb ({new_AGEMA_signal_1492, n2043}), .clk ( clk ), .rnd ({Fresh[1181], Fresh[1180]}), .outt ({new_AGEMA_signal_1599, n2048}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2195 ( .ina ({new_AGEMA_signal_1493, n2046}), .inb ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .rnd ({Fresh[1183], Fresh[1182]}), .outt ({new_AGEMA_signal_1600, n2047}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2206 ( .ina ({new_AGEMA_signal_1494, n2058}), .inb ({new_AGEMA_signal_1177, n2057}), .clk ( clk ), .rnd ({Fresh[1185], Fresh[1184]}), .outt ({new_AGEMA_signal_1601, n2059}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2213 ( .ina ({new_AGEMA_signal_1495, n2063}), .inb ({new_AGEMA_signal_1179, n2062}), .clk ( clk ), .rnd ({Fresh[1187], Fresh[1186]}), .outt ({new_AGEMA_signal_1602, n2064}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2229 ( .ina ({new_AGEMA_signal_1497, n2076}), .inb ({new_AGEMA_signal_1075, n2075}), .clk ( clk ), .rnd ({Fresh[1189], Fresh[1188]}), .outt ({new_AGEMA_signal_1603, n2077}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2249 ( .ina ({new_AGEMA_signal_1501, n2090}), .inb ({new_AGEMA_signal_1352, n2089}), .clk ( clk ), .rnd ({Fresh[1191], Fresh[1190]}), .outt ({new_AGEMA_signal_1604, n2158}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2255 ( .ina ({new_AGEMA_signal_1502, n2093}), .inb ({new_AGEMA_signal_1354, n2092}), .clk ( clk ), .rnd ({Fresh[1193], Fresh[1192]}), .outt ({new_AGEMA_signal_1605, n2095}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2274 ( .ina ({new_AGEMA_signal_1606, n2116}), .inb ({new_AGEMA_signal_1190, n2115}), .clk ( clk ), .rnd ({Fresh[1195], Fresh[1194]}), .outt ({new_AGEMA_signal_1681, n2117}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2283 ( .ina ({new_AGEMA_signal_1191, n2121}), .inb ({new_AGEMA_signal_1505, n2120}), .clk ( clk ), .rnd ({Fresh[1197], Fresh[1196]}), .outt ({new_AGEMA_signal_1607, n2123}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2300 ( .ina ({new_AGEMA_signal_1320, n2687}), .inb ({new_AGEMA_signal_1360, n2134}), .clk ( clk ), .rnd ({Fresh[1199], Fresh[1198]}), .outt ({new_AGEMA_signal_1507, n2135}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2309 ( .ina ({new_AGEMA_signal_1058, n2818}), .inb ({new_AGEMA_signal_1509, n2140}), .clk ( clk ), .rnd ({Fresh[1201], Fresh[1200]}), .outt ({new_AGEMA_signal_1609, n2141}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2327 ( .ina ({new_AGEMA_signal_1025, n2737}), .inb ({new_AGEMA_signal_1511, n2161}), .clk ( clk ), .rnd ({Fresh[1203], Fresh[1202]}), .outt ({new_AGEMA_signal_1610, n2166}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2331 ( .ina ({new_AGEMA_signal_978, n2694}), .inb ({new_AGEMA_signal_1367, n2164}), .clk ( clk ), .rnd ({Fresh[1205], Fresh[1204]}), .outt ({new_AGEMA_signal_1512, n2165}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2346 ( .ina ({new_AGEMA_signal_1513, n2179}), .inb ({new_AGEMA_signal_1050, n2766}), .clk ( clk ), .rnd ({Fresh[1207], Fresh[1206]}), .outt ({new_AGEMA_signal_1611, n2180}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2360 ( .ina ({new_AGEMA_signal_1372, n2193}), .inb ({new_AGEMA_signal_1514, n2192}), .clk ( clk ), .rnd ({Fresh[1209], Fresh[1208]}), .outt ({new_AGEMA_signal_1612, n2194}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2372 ( .ina ({new_AGEMA_signal_1613, n2203}), .inb ({new_AGEMA_signal_1516, n2202}), .clk ( clk ), .rnd ({Fresh[1211], Fresh[1210]}), .outt ({new_AGEMA_signal_1688, n2204}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2389 ( .ina ({new_AGEMA_signal_1517, n2224}), .inb ({new_AGEMA_signal_1518, n2223}), .clk ( clk ), .rnd ({Fresh[1213], Fresh[1212]}), .outt ({new_AGEMA_signal_1614, n2225}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2394 ( .ina ({new_AGEMA_signal_1379, n2229}), .inb ({new_AGEMA_signal_1214, n2228}), .clk ( clk ), .rnd ({Fresh[1215], Fresh[1214]}), .outt ({new_AGEMA_signal_1519, n2230}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2400 ( .ina ({new_AGEMA_signal_1315, n2235}), .inb ({new_AGEMA_signal_1616, n2234}), .clk ( clk ), .rnd ({Fresh[1217], Fresh[1216]}), .outt ({new_AGEMA_signal_1690, n2236}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2412 ( .ina ({new_AGEMA_signal_1521, n2246}), .inb ({new_AGEMA_signal_1220, n2245}), .clk ( clk ), .rnd ({Fresh[1219], Fresh[1218]}), .outt ({new_AGEMA_signal_1617, n2247}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2419 ( .ina ({new_AGEMA_signal_1522, n2254}), .inb ({new_AGEMA_signal_989, n2785}), .clk ( clk ), .rnd ({Fresh[1221], Fresh[1220]}), .outt ({new_AGEMA_signal_1618, n2255}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2427 ( .ina ({new_AGEMA_signal_1523, n2263}), .inb ({new_AGEMA_signal_1091, n2262}), .clk ( clk ), .rnd ({Fresh[1223], Fresh[1222]}), .outt ({new_AGEMA_signal_1619, n2264}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2435 ( .ina ({new_AGEMA_signal_1525, n2752}), .inb ({new_AGEMA_signal_1385, n2267}), .clk ( clk ), .rnd ({Fresh[1225], Fresh[1224]}), .outt ({new_AGEMA_signal_1620, n2271}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2446 ( .ina ({new_AGEMA_signal_983, n2815}), .inb ({new_AGEMA_signal_1387, n2279}), .clk ( clk ), .rnd ({Fresh[1227], Fresh[1226]}), .outt ({new_AGEMA_signal_1526, n2280}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2451 ( .ina ({SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_1388, n2283}), .clk ( clk ), .rnd ({Fresh[1229], Fresh[1228]}), .outt ({new_AGEMA_signal_1527, n2286}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2461 ( .ina ({new_AGEMA_signal_1529, n2686}), .inb ({new_AGEMA_signal_1530, n2289}), .clk ( clk ), .rnd ({Fresh[1231], Fresh[1230]}), .outt ({new_AGEMA_signal_1622, n2304}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2466 ( .ina ({new_AGEMA_signal_1393, n2293}), .inb ({new_AGEMA_signal_1532, n2292}), .clk ( clk ), .rnd ({Fresh[1233], Fresh[1232]}), .outt ({new_AGEMA_signal_1623, n2295}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2488 ( .ina ({new_AGEMA_signal_1534, n2321}), .inb ({new_AGEMA_signal_1233, n2320}), .clk ( clk ), .rnd ({Fresh[1235], Fresh[1234]}), .outt ({new_AGEMA_signal_1624, n2322}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2499 ( .ina ({new_AGEMA_signal_1535, n2332}), .inb ({new_AGEMA_signal_1536, n2331}), .clk ( clk ), .rnd ({Fresh[1237], Fresh[1236]}), .outt ({new_AGEMA_signal_1625, n2333}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2509 ( .ina ({new_AGEMA_signal_1237, n2343}), .inb ({new_AGEMA_signal_1538, n2342}), .clk ( clk ), .rnd ({Fresh[1239], Fresh[1238]}), .outt ({new_AGEMA_signal_1627, n2345}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2526 ( .ina ({new_AGEMA_signal_1539, n2358}), .inb ({new_AGEMA_signal_1402, n2357}), .clk ( clk ), .rnd ({Fresh[1241], Fresh[1240]}), .outt ({new_AGEMA_signal_1628, n2361}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2549 ( .ina ({new_AGEMA_signal_1406, n2387}), .inb ({new_AGEMA_signal_1407, n2386}), .clk ( clk ), .rnd ({Fresh[1243], Fresh[1242]}), .outt ({new_AGEMA_signal_1541, n2388}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2556 ( .ina ({new_AGEMA_signal_949, n2760}), .inb ({new_AGEMA_signal_1542, n2392}), .clk ( clk ), .rnd ({Fresh[1245], Fresh[1244]}), .outt ({new_AGEMA_signal_1630, n2393}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2567 ( .ina ({new_AGEMA_signal_1027, n2789}), .inb ({new_AGEMA_signal_1410, n2404}), .clk ( clk ), .rnd ({Fresh[1247], Fresh[1246]}), .outt ({new_AGEMA_signal_1543, n2405}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2571 ( .ina ({new_AGEMA_signal_1544, n2409}), .inb ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .rnd ({Fresh[1249], Fresh[1248]}), .outt ({new_AGEMA_signal_1632, n2410}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2576 ( .ina ({new_AGEMA_signal_955, n2630}), .inb ({new_AGEMA_signal_1545, n2414}), .clk ( clk ), .rnd ({Fresh[1251], Fresh[1250]}), .outt ({new_AGEMA_signal_1633, n2421}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2579 ( .ina ({new_AGEMA_signal_1413, n2418}), .inb ({new_AGEMA_signal_1324, n2417}), .clk ( clk ), .rnd ({Fresh[1253], Fresh[1252]}), .outt ({new_AGEMA_signal_1546, n2419}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2590 ( .ina ({new_AGEMA_signal_1414, n2433}), .inb ({new_AGEMA_signal_1547, n2432}), .clk ( clk ), .rnd ({Fresh[1255], Fresh[1254]}), .outt ({new_AGEMA_signal_1635, n2436}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2604 ( .ina ({new_AGEMA_signal_1548, n2449}), .inb ({new_AGEMA_signal_1549, n2448}), .clk ( clk ), .rnd ({Fresh[1257], Fresh[1256]}), .outt ({new_AGEMA_signal_1636, n2450}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2610 ( .ina ({new_AGEMA_signal_1063, n2823}), .inb ({new_AGEMA_signal_1550, n2455}), .clk ( clk ), .rnd ({Fresh[1259], Fresh[1258]}), .outt ({new_AGEMA_signal_1637, n2456}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2613 ( .ina ({new_AGEMA_signal_1551, n2460}), .inb ({new_AGEMA_signal_1390, n2459}), .clk ( clk ), .rnd ({Fresh[1261], Fresh[1260]}), .outt ({new_AGEMA_signal_1638, n2461}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2619 ( .ina ({new_AGEMA_signal_1246, n2467}), .inb ({new_AGEMA_signal_1422, n2466}), .clk ( clk ), .rnd ({Fresh[1263], Fresh[1262]}), .outt ({new_AGEMA_signal_1552, n2469}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2630 ( .ina ({new_AGEMA_signal_970, n2719}), .inb ({new_AGEMA_signal_1423, n2477}), .clk ( clk ), .rnd ({Fresh[1265], Fresh[1264]}), .outt ({new_AGEMA_signal_1553, n2478}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2635 ( .ina ({new_AGEMA_signal_1107, n2483}), .inb ({new_AGEMA_signal_1554, n2482}), .clk ( clk ), .rnd ({Fresh[1267], Fresh[1266]}), .outt ({new_AGEMA_signal_1640, n2484}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2643 ( .ina ({new_AGEMA_signal_1425, n2490}), .inb ({new_AGEMA_signal_1266, n2489}), .clk ( clk ), .rnd ({Fresh[1269], Fresh[1268]}), .outt ({new_AGEMA_signal_1555, n2491}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2649 ( .ina ({new_AGEMA_signal_1267, n2497}), .inb ({new_AGEMA_signal_1556, n2496}), .clk ( clk ), .rnd ({Fresh[1271], Fresh[1270]}), .outt ({new_AGEMA_signal_1642, n2500}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2656 ( .ina ({new_AGEMA_signal_1643, n2507}), .inb ({new_AGEMA_signal_1427, n2506}), .clk ( clk ), .rnd ({Fresh[1273], Fresh[1272]}), .outt ({new_AGEMA_signal_1708, n2508}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2670 ( .ina ({new_AGEMA_signal_1644, n2525}), .inb ({new_AGEMA_signal_1559, n2524}), .clk ( clk ), .rnd ({Fresh[1275], Fresh[1274]}), .outt ({new_AGEMA_signal_1709, n2526}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2679 ( .ina ({new_AGEMA_signal_1560, n2537}), .inb ({new_AGEMA_signal_1561, n2536}), .clk ( clk ), .rnd ({Fresh[1277], Fresh[1276]}), .outt ({new_AGEMA_signal_1645, n2539}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2682 ( .ina ({new_AGEMA_signal_1506, n2543}), .inb ({new_AGEMA_signal_1433, n2542}), .clk ( clk ), .rnd ({Fresh[1279], Fresh[1278]}), .outt ({new_AGEMA_signal_1646, n2548}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2694 ( .ina ({new_AGEMA_signal_1436, n2558}), .inb ({new_AGEMA_signal_1562, n2557}), .clk ( clk ), .rnd ({Fresh[1281], Fresh[1280]}), .outt ({new_AGEMA_signal_1647, n2568}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2700 ( .ina ({new_AGEMA_signal_1438, n2566}), .inb ({new_AGEMA_signal_1563, n2565}), .clk ( clk ), .rnd ({Fresh[1283], Fresh[1282]}), .outt ({new_AGEMA_signal_1648, n2567}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2710 ( .ina ({new_AGEMA_signal_1276, n2581}), .inb ({new_AGEMA_signal_1565, n2580}), .clk ( clk ), .rnd ({Fresh[1285], Fresh[1284]}), .outt ({new_AGEMA_signal_1649, n2583}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2728 ( .ina ({new_AGEMA_signal_1446, n2603}), .inb ({new_AGEMA_signal_1282, n2602}), .clk ( clk ), .rnd ({Fresh[1287], Fresh[1286]}), .outt ({new_AGEMA_signal_1566, n2604}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2739 ( .ina ({new_AGEMA_signal_1447, n2620}), .inb ({new_AGEMA_signal_1567, n2619}), .clk ( clk ), .rnd ({Fresh[1289], Fresh[1288]}), .outt ({new_AGEMA_signal_1651, n2621}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2745 ( .ina ({new_AGEMA_signal_1120, n2629}), .inb ({new_AGEMA_signal_1568, n2628}), .clk ( clk ), .rnd ({Fresh[1291], Fresh[1290]}), .outt ({new_AGEMA_signal_1652, n2633}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2756 ( .ina ({new_AGEMA_signal_1569, n2649}), .inb ({new_AGEMA_signal_1451, n2648}), .clk ( clk ), .rnd ({Fresh[1293], Fresh[1292]}), .outt ({new_AGEMA_signal_1653, n2660}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2759 ( .ina ({new_AGEMA_signal_1289, n2653}), .inb ({new_AGEMA_signal_1496, n2652}), .clk ( clk ), .rnd ({Fresh[1295], Fresh[1294]}), .outt ({new_AGEMA_signal_1654, n2656}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2766 ( .ina ({new_AGEMA_signal_1313, n2665}), .inb ({new_AGEMA_signal_1570, n2664}), .clk ( clk ), .rnd ({Fresh[1297], Fresh[1296]}), .outt ({new_AGEMA_signal_1655, n2666}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2774 ( .ina ({new_AGEMA_signal_1571, n2681}), .inb ({new_AGEMA_signal_1454, n2680}), .clk ( clk ), .rnd ({Fresh[1299], Fresh[1298]}), .outt ({new_AGEMA_signal_1656, n2706}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2777 ( .ina ({new_AGEMA_signal_1529, n2686}), .inb ({new_AGEMA_signal_1572, n2685}), .clk ( clk ), .rnd ({Fresh[1301], Fresh[1300]}), .outt ({new_AGEMA_signal_1657, n2704}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2781 ( .ina ({new_AGEMA_signal_1574, n2692}), .inb ({new_AGEMA_signal_1292, n2691}), .clk ( clk ), .rnd ({Fresh[1303], Fresh[1302]}), .outt ({new_AGEMA_signal_1658, n2696}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2794 ( .ina ({new_AGEMA_signal_1456, n2717}), .inb ({new_AGEMA_signal_1575, n2716}), .clk ( clk ), .rnd ({Fresh[1305], Fresh[1304]}), .outt ({new_AGEMA_signal_1659, n2718}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2801 ( .ina ({new_AGEMA_signal_1576, n2729}), .inb ({new_AGEMA_signal_1457, n2728}), .clk ( clk ), .rnd ({Fresh[1307], Fresh[1306]}), .outt ({new_AGEMA_signal_1660, n2730}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2805 ( .ina ({new_AGEMA_signal_1051, n2736}), .inb ({new_AGEMA_signal_1577, n2735}), .clk ( clk ), .rnd ({Fresh[1309], Fresh[1308]}), .outt ({new_AGEMA_signal_1661, n2745}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2809 ( .ina ({new_AGEMA_signal_1578, n2743}), .inb ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .rnd ({Fresh[1311], Fresh[1310]}), .outt ({new_AGEMA_signal_1662, n2744}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2814 ( .ina ({new_AGEMA_signal_1525, n2752}), .inb ({new_AGEMA_signal_1460, n2751}), .clk ( clk ), .rnd ({Fresh[1313], Fresh[1312]}), .outt ({new_AGEMA_signal_1663, n2759}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2821 ( .ina ({new_AGEMA_signal_957, n2765}), .inb ({new_AGEMA_signal_1580, n2764}), .clk ( clk ), .rnd ({Fresh[1315], Fresh[1314]}), .outt ({new_AGEMA_signal_1664, n2771}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2833 ( .ina ({new_AGEMA_signal_1466, n2788}), .inb ({new_AGEMA_signal_1303, n2787}), .clk ( clk ), .rnd ({Fresh[1317], Fresh[1316]}), .outt ({new_AGEMA_signal_1582, n2798}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2850 ( .ina ({new_AGEMA_signal_1584, n2822}), .inb ({new_AGEMA_signal_1469, n2821}), .clk ( clk ), .rnd ({Fresh[1319], Fresh[1318]}), .outt ({new_AGEMA_signal_1666, n2826}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2001 ( .ina ({new_AGEMA_signal_1586, n1932}), .inb ({new_AGEMA_signal_1037, n2577}), .clk ( clk ), .rnd ({Fresh[1321], Fresh[1320]}), .outt ({new_AGEMA_signal_1667, n1933}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2051 ( .ina ({new_AGEMA_signal_1317, n1956}), .inb ({new_AGEMA_signal_1589, n1955}), .clk ( clk ), .rnd ({Fresh[1323], Fresh[1322]}), .outt ({new_AGEMA_signal_1668, n1958}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2067 ( .ina ({new_AGEMA_signal_1479, n1967}), .inb ({new_AGEMA_signal_963, n2595}), .clk ( clk ), .rnd ({Fresh[1325], Fresh[1324]}), .outt ({new_AGEMA_signal_1590, n1990}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2104 ( .ina ({new_AGEMA_signal_1482, n1978}), .inb ({new_AGEMA_signal_1592, n1977}), .clk ( clk ), .rnd ({Fresh[1327], Fresh[1326]}), .outt ({new_AGEMA_signal_1670, n1982}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2128 ( .ina ({new_AGEMA_signal_996, n2437}), .inb ({new_AGEMA_signal_1594, n1998}), .clk ( clk ), .rnd ({Fresh[1329], Fresh[1328]}), .outt ({new_AGEMA_signal_1671, n1999}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2148 ( .ina ({new_AGEMA_signal_1595, n2010}), .inb ({new_AGEMA_signal_1162, n2009}), .clk ( clk ), .rnd ({Fresh[1331], Fresh[1330]}), .outt ({new_AGEMA_signal_1672, n2011}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2165 ( .ina ({new_AGEMA_signal_1489, n2024}), .inb ({new_AGEMA_signal_1166, n2023}), .clk ( clk ), .rnd ({Fresh[1333], Fresh[1332]}), .outt ({new_AGEMA_signal_1596, n2025}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2179 ( .ina ({new_AGEMA_signal_1597, n2035}), .inb ({new_AGEMA_signal_1072, n2034}), .clk ( clk ), .rnd ({Fresh[1335], Fresh[1334]}), .outt ({new_AGEMA_signal_1674, n2036}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2196 ( .ina ({new_AGEMA_signal_1599, n2048}), .inb ({new_AGEMA_signal_1600, n2047}), .clk ( clk ), .rnd ({Fresh[1337], Fresh[1336]}), .outt ({new_AGEMA_signal_1675, n2049}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2207 ( .ina ({new_AGEMA_signal_970, n2719}), .inb ({new_AGEMA_signal_1601, n2059}), .clk ( clk ), .rnd ({Fresh[1339], Fresh[1338]}), .outt ({new_AGEMA_signal_1676, n2072}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2214 ( .ina ({new_AGEMA_signal_971, n2641}), .inb ({new_AGEMA_signal_1602, n2064}), .clk ( clk ), .rnd ({Fresh[1341], Fresh[1340]}), .outt ({new_AGEMA_signal_1677, n2067}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2230 ( .ina ({new_AGEMA_signal_974, n2699}), .inb ({new_AGEMA_signal_1603, n2077}), .clk ( clk ), .rnd ({Fresh[1343], Fresh[1342]}), .outt ({new_AGEMA_signal_1678, n2078}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2250 ( .ina ({new_AGEMA_signal_1500, n2091}), .inb ({new_AGEMA_signal_1604, n2158}), .clk ( clk ), .rnd ({Fresh[1345], Fresh[1344]}), .outt ({new_AGEMA_signal_1679, n2097}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2257 ( .ina ({new_AGEMA_signal_1605, n2095}), .inb ({new_AGEMA_signal_1355, n2094}), .clk ( clk ), .rnd ({Fresh[1347], Fresh[1346]}), .outt ({new_AGEMA_signal_1680, n2096}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2275 ( .ina ({SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1681, n2117}), .clk ( clk ), .rnd ({Fresh[1349], Fresh[1348]}), .outt ({new_AGEMA_signal_1735, n2128}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2285 ( .ina ({new_AGEMA_signal_1607, n2123}), .inb ({new_AGEMA_signal_1193, n2122}), .clk ( clk ), .rnd ({Fresh[1351], Fresh[1350]}), .outt ({new_AGEMA_signal_1682, n2124}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2301 ( .ina ({new_AGEMA_signal_1506, n2543}), .inb ({new_AGEMA_signal_1507, n2135}), .clk ( clk ), .rnd ({Fresh[1353], Fresh[1352]}), .outt ({new_AGEMA_signal_1608, n2148}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2310 ( .ina ({new_AGEMA_signal_1199, n2220}), .inb ({new_AGEMA_signal_1609, n2141}), .clk ( clk ), .rnd ({Fresh[1355], Fresh[1354]}), .outt ({new_AGEMA_signal_1683, n2142}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2325 ( .ina ({new_AGEMA_signal_1510, n2159}), .inb ({new_AGEMA_signal_1604, n2158}), .clk ( clk ), .rnd ({Fresh[1357], Fresh[1356]}), .outt ({new_AGEMA_signal_1684, n2168}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2332 ( .ina ({new_AGEMA_signal_1610, n2166}), .inb ({new_AGEMA_signal_1512, n2165}), .clk ( clk ), .rnd ({Fresh[1359], Fresh[1358]}), .outt ({new_AGEMA_signal_1685, n2167}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2347 ( .ina ({new_AGEMA_signal_1369, n2181}), .inb ({new_AGEMA_signal_1611, n2180}), .clk ( clk ), .rnd ({Fresh[1361], Fresh[1360]}), .outt ({new_AGEMA_signal_1686, n2184}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2361 ( .ina ({new_AGEMA_signal_1371, n2195}), .inb ({new_AGEMA_signal_1612, n2194}), .clk ( clk ), .rnd ({Fresh[1363], Fresh[1362]}), .outt ({new_AGEMA_signal_1687, n2197}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2373 ( .ina ({new_AGEMA_signal_1063, n2823}), .inb ({new_AGEMA_signal_1688, n2204}), .clk ( clk ), .rnd ({Fresh[1365], Fresh[1364]}), .outt ({new_AGEMA_signal_1741, n2205}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2390 ( .ina ({new_AGEMA_signal_1065, n2828}), .inb ({new_AGEMA_signal_1614, n2225}), .clk ( clk ), .rnd ({Fresh[1367], Fresh[1366]}), .outt ({new_AGEMA_signal_1689, n2232}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2395 ( .ina ({new_AGEMA_signal_1519, n2230}), .inb ({new_AGEMA_signal_1007, n2563}), .clk ( clk ), .rnd ({Fresh[1369], Fresh[1368]}), .outt ({new_AGEMA_signal_1615, n2231}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2401 ( .ina ({new_AGEMA_signal_1215, n2237}), .inb ({new_AGEMA_signal_1690, n2236}), .clk ( clk ), .rnd ({Fresh[1371], Fresh[1370]}), .outt ({new_AGEMA_signal_1743, n2239}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2413 ( .ina ({new_AGEMA_signal_1380, n2248}), .inb ({new_AGEMA_signal_1617, n2247}), .clk ( clk ), .rnd ({Fresh[1373], Fresh[1372]}), .outt ({new_AGEMA_signal_1691, n2250}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2428 ( .ina ({new_AGEMA_signal_970, n2719}), .inb ({new_AGEMA_signal_1619, n2264}), .clk ( clk ), .rnd ({Fresh[1375], Fresh[1374]}), .outt ({new_AGEMA_signal_1692, n2276}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2439 ( .ina ({new_AGEMA_signal_1620, n2271}), .inb ({new_AGEMA_signal_1386, n2270}), .clk ( clk ), .rnd ({Fresh[1377], Fresh[1376]}), .outt ({new_AGEMA_signal_1693, n2272}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2454 ( .ina ({new_AGEMA_signal_1527, n2286}), .inb ({new_AGEMA_signal_1528, n2285}), .clk ( clk ), .rnd ({Fresh[1379], Fresh[1378]}), .outt ({new_AGEMA_signal_1621, n2306}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2468 ( .ina ({new_AGEMA_signal_1623, n2295}), .inb ({new_AGEMA_signal_1230, n2294}), .clk ( clk ), .rnd ({Fresh[1381], Fresh[1380]}), .outt ({new_AGEMA_signal_1694, n2296}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2489 ( .ina ({new_AGEMA_signal_1395, n2323}), .inb ({new_AGEMA_signal_1624, n2322}), .clk ( clk ), .rnd ({Fresh[1383], Fresh[1382]}), .outt ({new_AGEMA_signal_1695, n2324}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2500 ( .ina ({new_AGEMA_signal_1397, n2334}), .inb ({new_AGEMA_signal_1625, n2333}), .clk ( clk ), .rnd ({Fresh[1385], Fresh[1384]}), .outt ({new_AGEMA_signal_1696, n2337}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2511 ( .ina ({new_AGEMA_signal_1627, n2345}), .inb ({new_AGEMA_signal_1239, n2344}), .clk ( clk ), .rnd ({Fresh[1387], Fresh[1386]}), .outt ({new_AGEMA_signal_1697, n2350}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2528 ( .ina ({new_AGEMA_signal_1628, n2361}), .inb ({new_AGEMA_signal_1403, n2360}), .clk ( clk ), .rnd ({Fresh[1389], Fresh[1388]}), .outt ({new_AGEMA_signal_1698, n2362}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2550 ( .ina ({new_AGEMA_signal_1246, n2467}), .inb ({new_AGEMA_signal_1541, n2388}), .clk ( clk ), .rnd ({Fresh[1391], Fresh[1390]}), .outt ({new_AGEMA_signal_1629, n2389}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2557 ( .ina ({new_AGEMA_signal_1249, n2394}), .inb ({new_AGEMA_signal_1630, n2393}), .clk ( clk ), .rnd ({Fresh[1393], Fresh[1392]}), .outt ({new_AGEMA_signal_1700, n2397}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2568 ( .ina ({new_AGEMA_signal_1409, n2406}), .inb ({new_AGEMA_signal_1543, n2405}), .clk ( clk ), .rnd ({Fresh[1395], Fresh[1394]}), .outt ({new_AGEMA_signal_1631, n2411}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2580 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1546, n2419}), .clk ( clk ), .rnd ({Fresh[1397], Fresh[1396]}), .outt ({new_AGEMA_signal_1634, n2420}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2593 ( .ina ({new_AGEMA_signal_1635, n2436}), .inb ({new_AGEMA_signal_1416, n2435}), .clk ( clk ), .rnd ({Fresh[1399], Fresh[1398]}), .outt ({new_AGEMA_signal_1703, n2440}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2614 ( .ina ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1638, n2461}), .clk ( clk ), .rnd ({Fresh[1401], Fresh[1400]}), .outt ({new_AGEMA_signal_1704, n2516}) ) ;
    mux2_HPC1 #(.security_order(1), .pipeline(0)) U2621 ( .ins ({SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_1552, n2469}), .ina ({new_AGEMA_signal_1110, n2468}), .clk ( clk ), .rnd ({Fresh[1403], Fresh[1402]}), .outt ({new_AGEMA_signal_1639, n2471}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2636 ( .ina ({new_AGEMA_signal_1144, n2761}), .inb ({new_AGEMA_signal_1640, n2484}), .clk ( clk ), .rnd ({Fresh[1405], Fresh[1404]}), .outt ({new_AGEMA_signal_1706, n2485}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2644 ( .ina ({new_AGEMA_signal_971, n2641}), .inb ({new_AGEMA_signal_1555, n2491}), .clk ( clk ), .rnd ({Fresh[1407], Fresh[1406]}), .outt ({new_AGEMA_signal_1641, n2502}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2651 ( .ina ({new_AGEMA_signal_1642, n2500}), .inb ({new_AGEMA_signal_1269, n2499}), .clk ( clk ), .rnd ({Fresh[1409], Fresh[1408]}), .outt ({new_AGEMA_signal_1707, n2501}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2657 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1708, n2508}), .clk ( clk ), .rnd ({Fresh[1411], Fresh[1410]}), .outt ({new_AGEMA_signal_1757, n2509}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2671 ( .ina ({new_AGEMA_signal_989, n2785}), .inb ({new_AGEMA_signal_1709, n2526}), .clk ( clk ), .rnd ({Fresh[1413], Fresh[1412]}), .outt ({new_AGEMA_signal_1758, n2527}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2680 ( .ina ({new_AGEMA_signal_1645, n2539}), .inb ({new_AGEMA_signal_985, n2538}), .clk ( clk ), .rnd ({Fresh[1415], Fresh[1414]}), .outt ({new_AGEMA_signal_1710, n2550}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2685 ( .ina ({new_AGEMA_signal_1646, n2548}), .inb ({new_AGEMA_signal_1434, n2547}), .clk ( clk ), .rnd ({Fresh[1417], Fresh[1416]}), .outt ({new_AGEMA_signal_1711, n2549}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2701 ( .ina ({new_AGEMA_signal_1647, n2568}), .inb ({new_AGEMA_signal_1648, n2567}), .clk ( clk ), .rnd ({Fresh[1419], Fresh[1418]}), .outt ({new_AGEMA_signal_1712, n2569}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2712 ( .ina ({new_AGEMA_signal_1649, n2583}), .inb ({new_AGEMA_signal_1443, n2582}), .clk ( clk ), .rnd ({Fresh[1421], Fresh[1420]}), .outt ({new_AGEMA_signal_1713, n2584}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2729 ( .ina ({new_AGEMA_signal_1445, n2605}), .inb ({new_AGEMA_signal_1566, n2604}), .clk ( clk ), .rnd ({Fresh[1423], Fresh[1422]}), .outt ({new_AGEMA_signal_1650, n2606}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2740 ( .ina ({new_AGEMA_signal_971, n2641}), .inb ({new_AGEMA_signal_1651, n2621}), .clk ( clk ), .rnd ({Fresh[1425], Fresh[1424]}), .outt ({new_AGEMA_signal_1715, n2622}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2747 ( .ina ({new_AGEMA_signal_1652, n2633}), .inb ({new_AGEMA_signal_1286, n2632}), .clk ( clk ), .rnd ({Fresh[1427], Fresh[1426]}), .outt ({new_AGEMA_signal_1716, n2634}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2761 ( .ina ({new_AGEMA_signal_1654, n2656}), .inb ({new_AGEMA_signal_1452, n2655}), .clk ( clk ), .rnd ({Fresh[1429], Fresh[1428]}), .outt ({new_AGEMA_signal_1717, n2657}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2783 ( .ina ({new_AGEMA_signal_1658, n2696}), .inb ({new_AGEMA_signal_1455, n2695}), .clk ( clk ), .rnd ({Fresh[1431], Fresh[1430]}), .outt ({new_AGEMA_signal_1718, n2697}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2795 ( .ina ({new_AGEMA_signal_970, n2719}), .inb ({new_AGEMA_signal_1659, n2718}), .clk ( clk ), .rnd ({Fresh[1433], Fresh[1432]}), .outt ({new_AGEMA_signal_1719, n2808}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2802 ( .ina ({new_AGEMA_signal_1660, n2730}), .inb ({new_AGEMA_signal_1067, n2809}), .clk ( clk ), .rnd ({Fresh[1435], Fresh[1434]}), .outt ({new_AGEMA_signal_1720, n2747}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2810 ( .ina ({new_AGEMA_signal_1661, n2745}), .inb ({new_AGEMA_signal_1662, n2744}), .clk ( clk ), .rnd ({Fresh[1437], Fresh[1436]}), .outt ({new_AGEMA_signal_1721, n2746}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2818 ( .ina ({new_AGEMA_signal_1663, n2759}), .inb ({new_AGEMA_signal_1579, n2758}), .clk ( clk ), .rnd ({Fresh[1439], Fresh[1438]}), .outt ({new_AGEMA_signal_1722, n2804}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2824 ( .ina ({new_AGEMA_signal_1664, n2771}), .inb ({new_AGEMA_signal_1463, n2770}), .clk ( clk ), .rnd ({Fresh[1441], Fresh[1440]}), .outt ({new_AGEMA_signal_1723, n2802}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2838 ( .ina ({new_AGEMA_signal_1582, n2798}), .inb ({new_AGEMA_signal_1583, n2797}), .clk ( clk ), .rnd ({Fresh[1443], Fresh[1442]}), .outt ({new_AGEMA_signal_1665, n2799}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2852 ( .ina ({new_AGEMA_signal_1666, n2826}), .inb ({new_AGEMA_signal_1308, n2825}), .clk ( clk ), .rnd ({Fresh[1445], Fresh[1444]}), .outt ({new_AGEMA_signal_1725, n2827}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2002 ( .ina ({new_AGEMA_signal_1585, n1934}), .inb ({new_AGEMA_signal_1667, n1933}), .clk ( clk ), .rnd ({Fresh[1447], Fresh[1446]}), .outt ({new_AGEMA_signal_1726, n1935}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2054 ( .ina ({new_AGEMA_signal_1668, n1958}), .inb ({new_AGEMA_signal_1049, n1957}), .clk ( clk ), .rnd ({Fresh[1449], Fresh[1448]}), .outt ({new_AGEMA_signal_1727, n1959}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2109 ( .ina ({new_AGEMA_signal_1670, n1982}), .inb ({new_AGEMA_signal_1593, n1981}), .clk ( clk ), .rnd ({Fresh[1451], Fresh[1450]}), .outt ({new_AGEMA_signal_1728, n1983}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2149 ( .ina ({new_AGEMA_signal_1487, n2012}), .inb ({new_AGEMA_signal_1672, n2011}), .clk ( clk ), .rnd ({Fresh[1453], Fresh[1452]}), .outt ({new_AGEMA_signal_1729, n2014}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2166 ( .ina ({new_AGEMA_signal_1069, n2026}), .inb ({new_AGEMA_signal_1596, n2025}), .clk ( clk ), .rnd ({Fresh[1455], Fresh[1454]}), .outt ({new_AGEMA_signal_1673, n2029}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2180 ( .ina ({new_AGEMA_signal_996, n2437}), .inb ({new_AGEMA_signal_1674, n2036}), .clk ( clk ), .rnd ({Fresh[1457], Fresh[1456]}), .outt ({new_AGEMA_signal_1731, n2037}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2197 ( .ina ({new_AGEMA_signal_1171, n2050}), .inb ({new_AGEMA_signal_1675, n2049}), .clk ( clk ), .rnd ({Fresh[1459], Fresh[1458]}), .outt ({new_AGEMA_signal_1732, n2052}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2219 ( .ina ({new_AGEMA_signal_1677, n2067}), .inb ({new_AGEMA_signal_1496, n2652}), .clk ( clk ), .rnd ({Fresh[1461], Fresh[1460]}), .outt ({new_AGEMA_signal_1733, n2070}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2258 ( .ina ({new_AGEMA_signal_1679, n2097}), .inb ({new_AGEMA_signal_1680, n2096}), .clk ( clk ), .rnd ({Fresh[1463], Fresh[1462]}), .outt ({new_AGEMA_signal_1734, n2098}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2287 ( .ina ({new_AGEMA_signal_1682, n2124}), .inb ({new_AGEMA_signal_1194, n2811}), .clk ( clk ), .rnd ({Fresh[1465], Fresh[1464]}), .outt ({new_AGEMA_signal_1736, n2125}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2311 ( .ina ({new_AGEMA_signal_1508, n2143}), .inb ({new_AGEMA_signal_1683, n2142}), .clk ( clk ), .rnd ({Fresh[1467], Fresh[1466]}), .outt ({new_AGEMA_signal_1737, n2145}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2333 ( .ina ({new_AGEMA_signal_1684, n2168}), .inb ({new_AGEMA_signal_1685, n2167}), .clk ( clk ), .rnd ({Fresh[1469], Fresh[1468]}), .outt ({new_AGEMA_signal_1738, n2169}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2350 ( .ina ({new_AGEMA_signal_1686, n2184}), .inb ({new_AGEMA_signal_1086, n2183}), .clk ( clk ), .rnd ({Fresh[1471], Fresh[1470]}), .outt ({new_AGEMA_signal_1739, n2185}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2365 ( .ina ({new_AGEMA_signal_1687, n2197}), .inb ({new_AGEMA_signal_1209, n2196}), .clk ( clk ), .rnd ({Fresh[1473], Fresh[1472]}), .outt ({new_AGEMA_signal_1740, n2198}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2396 ( .ina ({new_AGEMA_signal_1689, n2232}), .inb ({new_AGEMA_signal_1615, n2231}), .clk ( clk ), .rnd ({Fresh[1475], Fresh[1474]}), .outt ({new_AGEMA_signal_1742, n2312}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2404 ( .ina ({new_AGEMA_signal_1743, n2239}), .inb ({new_AGEMA_signal_1216, n2238}), .clk ( clk ), .rnd ({Fresh[1477], Fresh[1476]}), .outt ({new_AGEMA_signal_1781, n2258}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2415 ( .ina ({new_AGEMA_signal_1691, n2250}), .inb ({new_AGEMA_signal_1382, n2249}), .clk ( clk ), .rnd ({Fresh[1479], Fresh[1478]}), .outt ({new_AGEMA_signal_1744, n2251}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2440 ( .ina ({new_AGEMA_signal_1524, n2273}), .inb ({new_AGEMA_signal_1693, n2272}), .clk ( clk ), .rnd ({Fresh[1481], Fresh[1480]}), .outt ({new_AGEMA_signal_1745, n2274}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2469 ( .ina ({new_AGEMA_signal_1531, n2297}), .inb ({new_AGEMA_signal_1694, n2296}), .clk ( clk ), .rnd ({Fresh[1483], Fresh[1482]}), .outt ({new_AGEMA_signal_1746, n2302}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2490 ( .ina ({new_AGEMA_signal_1695, n2324}), .inb ({new_AGEMA_signal_1000, n2772}), .clk ( clk ), .rnd ({Fresh[1485], Fresh[1484]}), .outt ({new_AGEMA_signal_1747, n2339}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2503 ( .ina ({new_AGEMA_signal_1696, n2337}), .inb ({new_AGEMA_signal_1626, n2336}), .clk ( clk ), .rnd ({Fresh[1487], Fresh[1486]}), .outt ({new_AGEMA_signal_1748, n2338}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2515 ( .ina ({new_AGEMA_signal_1697, n2350}), .inb ({new_AGEMA_signal_1240, n2349}), .clk ( clk ), .rnd ({Fresh[1489], Fresh[1488]}), .outt ({new_AGEMA_signal_1749, n2351}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2529 ( .ina ({new_AGEMA_signal_1102, n2363}), .inb ({new_AGEMA_signal_1698, n2362}), .clk ( clk ), .rnd ({Fresh[1491], Fresh[1490]}), .outt ({new_AGEMA_signal_1750, n2365}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2551 ( .ina ({new_AGEMA_signal_1629, n2389}), .inb ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[1493], Fresh[1492]}), .outt ({new_AGEMA_signal_1699, n2399}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2560 ( .ina ({new_AGEMA_signal_1700, n2397}), .inb ({new_AGEMA_signal_1251, n2396}), .clk ( clk ), .rnd ({Fresh[1495], Fresh[1494]}), .outt ({new_AGEMA_signal_1751, n2398}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2572 ( .ina ({new_AGEMA_signal_1631, n2411}), .inb ({new_AGEMA_signal_1632, n2410}), .clk ( clk ), .rnd ({Fresh[1497], Fresh[1496]}), .outt ({new_AGEMA_signal_1701, n2423}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2581 ( .ina ({new_AGEMA_signal_1633, n2421}), .inb ({new_AGEMA_signal_1634, n2420}), .clk ( clk ), .rnd ({Fresh[1499], Fresh[1498]}), .outt ({new_AGEMA_signal_1702, n2422}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2596 ( .ina ({new_AGEMA_signal_1703, n2440}), .inb ({new_AGEMA_signal_1417, n2439}), .clk ( clk ), .rnd ({Fresh[1501], Fresh[1500]}), .outt ({new_AGEMA_signal_1753, n2441}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2623 ( .ina ({new_AGEMA_signal_1639, n2471}), .inb ({new_AGEMA_signal_1261, n2470}), .clk ( clk ), .rnd ({Fresh[1503], Fresh[1502]}), .outt ({new_AGEMA_signal_1705, n2479}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2637 ( .ina ({new_AGEMA_signal_1706, n2485}), .inb ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .rnd ({Fresh[1505], Fresh[1504]}), .outt ({new_AGEMA_signal_1755, n2512}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2652 ( .ina ({new_AGEMA_signal_1641, n2502}), .inb ({new_AGEMA_signal_1707, n2501}), .clk ( clk ), .rnd ({Fresh[1507], Fresh[1506]}), .outt ({new_AGEMA_signal_1756, n2510}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2686 ( .ina ({new_AGEMA_signal_1710, n2550}), .inb ({new_AGEMA_signal_1711, n2549}), .clk ( clk ), .rnd ({Fresh[1509], Fresh[1508]}), .outt ({new_AGEMA_signal_1759, n2552}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2702 ( .ina ({new_AGEMA_signal_1044, n2570}), .inb ({new_AGEMA_signal_1712, n2569}), .clk ( clk ), .rnd ({Fresh[1511], Fresh[1510]}), .outt ({new_AGEMA_signal_1760, n2593}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2713 ( .ina ({new_AGEMA_signal_1441, n2585}), .inb ({new_AGEMA_signal_1713, n2584}), .clk ( clk ), .rnd ({Fresh[1513], Fresh[1512]}), .outt ({new_AGEMA_signal_1761, n2589}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2730 ( .ina ({new_AGEMA_signal_1279, n2607}), .inb ({new_AGEMA_signal_1650, n2606}), .clk ( clk ), .rnd ({Fresh[1515], Fresh[1514]}), .outt ({new_AGEMA_signal_1714, n2608}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2748 ( .ina ({new_AGEMA_signal_958, n2635}), .inb ({new_AGEMA_signal_1716, n2634}), .clk ( clk ), .rnd ({Fresh[1517], Fresh[1516]}), .outt ({new_AGEMA_signal_1763, n2636}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2762 ( .ina ({new_AGEMA_signal_1478, n2658}), .inb ({new_AGEMA_signal_1717, n2657}), .clk ( clk ), .rnd ({Fresh[1519], Fresh[1518]}), .outt ({new_AGEMA_signal_1764, n2659}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2784 ( .ina ({new_AGEMA_signal_1573, n2698}), .inb ({new_AGEMA_signal_1718, n2697}), .clk ( clk ), .rnd ({Fresh[1521], Fresh[1520]}), .outt ({new_AGEMA_signal_1765, n2702}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2811 ( .ina ({new_AGEMA_signal_1720, n2747}), .inb ({new_AGEMA_signal_1721, n2746}), .clk ( clk ), .rnd ({Fresh[1523], Fresh[1522]}), .outt ({new_AGEMA_signal_1766, n2806}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2839 ( .ina ({new_AGEMA_signal_1581, n2800}), .inb ({new_AGEMA_signal_1665, n2799}), .clk ( clk ), .rnd ({Fresh[1525], Fresh[1524]}), .outt ({new_AGEMA_signal_1724, n2801}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2853 ( .ina ({new_AGEMA_signal_1065, n2828}), .inb ({new_AGEMA_signal_1725, n2827}), .clk ( clk ), .rnd ({Fresh[1527], Fresh[1526]}), .outt ({new_AGEMA_signal_1768, n2829}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2003 ( .ina ({new_AGEMA_signal_1470, n1936}), .inb ({new_AGEMA_signal_1726, n1935}), .clk ( clk ), .rnd ({Fresh[1529], Fresh[1528]}), .outt ({new_AGEMA_signal_1769, n1941}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2059 ( .ina ({new_AGEMA_signal_1727, n1959}), .inb ({new_AGEMA_signal_1478, n2658}), .clk ( clk ), .rnd ({Fresh[1531], Fresh[1530]}), .outt ({new_AGEMA_signal_1770, n1960}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2110 ( .ina ({new_AGEMA_signal_1669, n1984}), .inb ({new_AGEMA_signal_1728, n1983}), .clk ( clk ), .rnd ({Fresh[1533], Fresh[1532]}), .outt ({new_AGEMA_signal_1771, n1988}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2153 ( .ina ({new_AGEMA_signal_1729, n2014}), .inb ({new_AGEMA_signal_1335, n2013}), .clk ( clk ), .rnd ({Fresh[1535], Fresh[1534]}), .outt ({new_AGEMA_signal_1772, n2015}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2169 ( .ina ({new_AGEMA_signal_1673, n2029}), .inb ({new_AGEMA_signal_1071, n2028}), .clk ( clk ), .rnd ({Fresh[1537], Fresh[1536]}), .outt ({new_AGEMA_signal_1730, n2030}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2200 ( .ina ({new_AGEMA_signal_1732, n2052}), .inb ({new_AGEMA_signal_1341, n2051}), .clk ( clk ), .rnd ({Fresh[1539], Fresh[1538]}), .outt ({new_AGEMA_signal_1774, n2053}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2222 ( .ina ({new_AGEMA_signal_1733, n2070}), .inb ({new_AGEMA_signal_1346, n2069}), .clk ( clk ), .rnd ({Fresh[1541], Fresh[1540]}), .outt ({new_AGEMA_signal_1775, n2071}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2259 ( .ina ({new_AGEMA_signal_1499, n2099}), .inb ({new_AGEMA_signal_1734, n2098}), .clk ( clk ), .rnd ({Fresh[1543], Fresh[1542]}), .outt ({new_AGEMA_signal_1776, n2103}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2288 ( .ina ({new_AGEMA_signal_1079, n2544}), .inb ({new_AGEMA_signal_1736, n2125}), .clk ( clk ), .rnd ({Fresh[1545], Fresh[1544]}), .outt ({new_AGEMA_signal_1777, n2126}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2314 ( .ina ({new_AGEMA_signal_1737, n2145}), .inb ({new_AGEMA_signal_1363, n2144}), .clk ( clk ), .rnd ({Fresh[1547], Fresh[1546]}), .outt ({new_AGEMA_signal_1778, n2146}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2334 ( .ina ({new_AGEMA_signal_1365, n2170}), .inb ({new_AGEMA_signal_1738, n2169}), .clk ( clk ), .rnd ({Fresh[1549], Fresh[1548]}), .outt ({new_AGEMA_signal_1779, n2173}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2351 ( .ina ({new_AGEMA_signal_1084, n2186}), .inb ({new_AGEMA_signal_1739, n2185}), .clk ( clk ), .rnd ({Fresh[1551], Fresh[1550]}), .outt ({new_AGEMA_signal_1780, n2187}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2416 ( .ina ({new_AGEMA_signal_996, n2437}), .inb ({new_AGEMA_signal_1744, n2251}), .clk ( clk ), .rnd ({Fresh[1553], Fresh[1552]}), .outt ({new_AGEMA_signal_1782, n2256}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2441 ( .ina ({new_AGEMA_signal_1745, n2274}), .inb ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[1555], Fresh[1554]}), .outt ({new_AGEMA_signal_1783, n2275}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2474 ( .ina ({new_AGEMA_signal_1746, n2302}), .inb ({new_AGEMA_signal_1533, n2301}), .clk ( clk ), .rnd ({Fresh[1557], Fresh[1556]}), .outt ({new_AGEMA_signal_1784, n2303}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2504 ( .ina ({new_AGEMA_signal_1747, n2339}), .inb ({new_AGEMA_signal_1748, n2338}), .clk ( clk ), .rnd ({Fresh[1559], Fresh[1558]}), .outt ({new_AGEMA_signal_1785, n2382}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2516 ( .ina ({new_AGEMA_signal_1749, n2351}), .inb ({new_AGEMA_signal_971, n2641}), .clk ( clk ), .rnd ({Fresh[1561], Fresh[1560]}), .outt ({new_AGEMA_signal_1786, n2380}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2531 ( .ina ({new_AGEMA_signal_1750, n2365}), .inb ({new_AGEMA_signal_1245, n2364}), .clk ( clk ), .rnd ({Fresh[1563], Fresh[1562]}), .outt ({new_AGEMA_signal_1787, n2366}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2561 ( .ina ({new_AGEMA_signal_1699, n2399}), .inb ({new_AGEMA_signal_1751, n2398}), .clk ( clk ), .rnd ({Fresh[1565], Fresh[1564]}), .outt ({new_AGEMA_signal_1788, n2425}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2582 ( .ina ({new_AGEMA_signal_1701, n2423}), .inb ({new_AGEMA_signal_1702, n2422}), .clk ( clk ), .rnd ({Fresh[1567], Fresh[1566]}), .outt ({new_AGEMA_signal_1752, n2424}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2597 ( .ina ({new_AGEMA_signal_1031, n2688}), .inb ({new_AGEMA_signal_1753, n2441}), .clk ( clk ), .rnd ({Fresh[1569], Fresh[1568]}), .outt ({new_AGEMA_signal_1789, n2451}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2631 ( .ina ({new_AGEMA_signal_1705, n2479}), .inb ({new_AGEMA_signal_1553, n2478}), .clk ( clk ), .rnd ({Fresh[1571], Fresh[1570]}), .outt ({new_AGEMA_signal_1754, n2514}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2658 ( .ina ({new_AGEMA_signal_1756, n2510}), .inb ({new_AGEMA_signal_1757, n2509}), .clk ( clk ), .rnd ({Fresh[1573], Fresh[1572]}), .outt ({new_AGEMA_signal_1790, n2511}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2688 ( .ina ({new_AGEMA_signal_1759, n2552}), .inb ({new_AGEMA_signal_1435, n2551}), .clk ( clk ), .rnd ({Fresh[1575], Fresh[1574]}), .outt ({new_AGEMA_signal_1791, n2671}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2716 ( .ina ({new_AGEMA_signal_1761, n2589}), .inb ({new_AGEMA_signal_1444, n2588}), .clk ( clk ), .rnd ({Fresh[1577], Fresh[1576]}), .outt ({new_AGEMA_signal_1792, n2590}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2731 ( .ina ({new_AGEMA_signal_1714, n2608}), .inb ({new_AGEMA_signal_1050, n2766}), .clk ( clk ), .rnd ({Fresh[1579], Fresh[1578]}), .outt ({new_AGEMA_signal_1762, n2623}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2763 ( .ina ({new_AGEMA_signal_1653, n2660}), .inb ({new_AGEMA_signal_1764, n2659}), .clk ( clk ), .rnd ({Fresh[1581], Fresh[1580]}), .outt ({new_AGEMA_signal_1794, n2667}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2786 ( .ina ({new_AGEMA_signal_1765, n2702}), .inb ({new_AGEMA_signal_1293, n2701}), .clk ( clk ), .rnd ({Fresh[1583], Fresh[1582]}), .outt ({new_AGEMA_signal_1795, n2703}) ) ;
    mux2_HPC1 #(.security_order(1), .pipeline(0)) U2840 ( .ins ({SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1723, n2802}), .ina ({new_AGEMA_signal_1724, n2801}), .clk ( clk ), .rnd ({Fresh[1585], Fresh[1584]}), .outt ({new_AGEMA_signal_1767, n2803}) ) ;

    /* cells in depth 17 */

    /* cells in depth 18 */
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2016 ( .ina ({new_AGEMA_signal_1769, n1941}), .inb ({new_AGEMA_signal_1587, n1940}), .clk ( clk ), .rnd ({Fresh[1587], Fresh[1586]}), .outt ({new_AGEMA_signal_1797, n2019}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2060 ( .ina ({new_AGEMA_signal_1588, n1961}), .inb ({new_AGEMA_signal_1770, n1960}), .clk ( clk ), .rnd ({Fresh[1589], Fresh[1588]}), .outt ({new_AGEMA_signal_1798, n2002}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2116 ( .ina ({new_AGEMA_signal_1771, n1988}), .inb ({new_AGEMA_signal_1485, n1987}), .clk ( clk ), .rnd ({Fresh[1591], Fresh[1590]}), .outt ({new_AGEMA_signal_1799, n1989}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2154 ( .ina ({new_AGEMA_signal_1065, n2828}), .inb ({new_AGEMA_signal_1772, n2015}), .clk ( clk ), .rnd ({Fresh[1593], Fresh[1592]}), .outt ({new_AGEMA_signal_1800, n2016}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2170 ( .ina ({new_AGEMA_signal_986, n2742}), .inb ({new_AGEMA_signal_1730, n2030}), .clk ( clk ), .rnd ({Fresh[1595], Fresh[1594]}), .outt ({new_AGEMA_signal_1773, n2038}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2201 ( .ina ({new_AGEMA_signal_1598, n2054}), .inb ({new_AGEMA_signal_1774, n2053}), .clk ( clk ), .rnd ({Fresh[1597], Fresh[1596]}), .outt ({new_AGEMA_signal_1802, n2111}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2223 ( .ina ({new_AGEMA_signal_1676, n2072}), .inb ({new_AGEMA_signal_1775, n2071}), .clk ( clk ), .rnd ({Fresh[1599], Fresh[1598]}), .outt ({new_AGEMA_signal_1803, n2079}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2263 ( .ina ({new_AGEMA_signal_1776, n2103}), .inb ({new_AGEMA_signal_1503, n2102}), .clk ( clk ), .rnd ({Fresh[1601], Fresh[1600]}), .outt ({new_AGEMA_signal_1804, n2104}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2289 ( .ina ({new_AGEMA_signal_1023, n2672}), .inb ({new_AGEMA_signal_1777, n2126}), .clk ( clk ), .rnd ({Fresh[1603], Fresh[1602]}), .outt ({new_AGEMA_signal_1805, n2127}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2315 ( .ina ({new_AGEMA_signal_1065, n2828}), .inb ({new_AGEMA_signal_1778, n2146}), .clk ( clk ), .rnd ({Fresh[1605], Fresh[1604]}), .outt ({new_AGEMA_signal_1806, n2147}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2336 ( .ina ({new_AGEMA_signal_1779, n2173}), .inb ({new_AGEMA_signal_1368, n2172}), .clk ( clk ), .rnd ({Fresh[1607], Fresh[1606]}), .outt ({new_AGEMA_signal_1807, n2208}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2352 ( .ina ({new_AGEMA_signal_1780, n2187}), .inb ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .rnd ({Fresh[1609], Fresh[1608]}), .outt ({new_AGEMA_signal_1808, n2199}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2420 ( .ina ({new_AGEMA_signal_1782, n2256}), .inb ({new_AGEMA_signal_1618, n2255}), .clk ( clk ), .rnd ({Fresh[1611], Fresh[1610]}), .outt ({new_AGEMA_signal_1809, n2257}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2442 ( .ina ({new_AGEMA_signal_1692, n2276}), .inb ({new_AGEMA_signal_1783, n2275}), .clk ( clk ), .rnd ({Fresh[1613], Fresh[1612]}), .outt ({new_AGEMA_signal_1810, n2281}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2475 ( .ina ({new_AGEMA_signal_1622, n2304}), .inb ({new_AGEMA_signal_1784, n2303}), .clk ( clk ), .rnd ({Fresh[1615], Fresh[1614]}), .outt ({new_AGEMA_signal_1811, n2305}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2532 ( .ina ({new_AGEMA_signal_1400, n2367}), .inb ({new_AGEMA_signal_1787, n2366}), .clk ( clk ), .rnd ({Fresh[1617], Fresh[1616]}), .outt ({new_AGEMA_signal_1812, n2368}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2583 ( .ina ({new_AGEMA_signal_1788, n2425}), .inb ({new_AGEMA_signal_1752, n2424}), .clk ( clk ), .rnd ({Fresh[1619], Fresh[1618]}), .outt ({new_AGEMA_signal_1813, n2426}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2605 ( .ina ({new_AGEMA_signal_1789, n2451}), .inb ({new_AGEMA_signal_1636, n2450}), .clk ( clk ), .rnd ({Fresh[1621], Fresh[1620]}), .outt ({new_AGEMA_signal_1814, n2457}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2659 ( .ina ({new_AGEMA_signal_1755, n2512}), .inb ({new_AGEMA_signal_1790, n2511}), .clk ( clk ), .rnd ({Fresh[1623], Fresh[1622]}), .outt ({new_AGEMA_signal_1815, n2513}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2717 ( .ina ({new_AGEMA_signal_1564, n2591}), .inb ({new_AGEMA_signal_1792, n2590}), .clk ( clk ), .rnd ({Fresh[1625], Fresh[1624]}), .outt ({new_AGEMA_signal_1816, n2592}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2741 ( .ina ({new_AGEMA_signal_1762, n2623}), .inb ({new_AGEMA_signal_1715, n2622}), .clk ( clk ), .rnd ({Fresh[1627], Fresh[1626]}), .outt ({new_AGEMA_signal_1793, n2637}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2767 ( .ina ({new_AGEMA_signal_1794, n2667}), .inb ({new_AGEMA_signal_1655, n2666}), .clk ( clk ), .rnd ({Fresh[1629], Fresh[1628]}), .outt ({new_AGEMA_signal_1818, n2668}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2787 ( .ina ({new_AGEMA_signal_1657, n2704}), .inb ({new_AGEMA_signal_1795, n2703}), .clk ( clk ), .rnd ({Fresh[1631], Fresh[1630]}), .outt ({new_AGEMA_signal_1819, n2705}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2841 ( .ina ({new_AGEMA_signal_1722, n2804}), .inb ({new_AGEMA_signal_1767, n2803}), .clk ( clk ), .rnd ({Fresh[1633], Fresh[1632]}), .outt ({new_AGEMA_signal_1796, n2805}) ) ;

    /* cells in depth 19 */

    /* cells in depth 20 */
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2117 ( .ina ({new_AGEMA_signal_1590, n1990}), .inb ({new_AGEMA_signal_1799, n1989}), .clk ( clk ), .rnd ({Fresh[1635], Fresh[1634]}), .outt ({new_AGEMA_signal_1821, n2000}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2181 ( .ina ({new_AGEMA_signal_1773, n2038}), .inb ({new_AGEMA_signal_1731, n2037}), .clk ( clk ), .rnd ({Fresh[1637], Fresh[1636]}), .outt ({new_AGEMA_signal_1801, n2113}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2231 ( .ina ({new_AGEMA_signal_1803, n2079}), .inb ({new_AGEMA_signal_1678, n2078}), .clk ( clk ), .rnd ({Fresh[1639], Fresh[1638]}), .outt ({new_AGEMA_signal_1822, n2109}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2264 ( .ina ({new_AGEMA_signal_1498, n2105}), .inb ({new_AGEMA_signal_1804, n2104}), .clk ( clk ), .rnd ({Fresh[1641], Fresh[1640]}), .outt ({new_AGEMA_signal_1823, n2107}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2290 ( .ina ({new_AGEMA_signal_1735, n2128}), .inb ({new_AGEMA_signal_1805, n2127}), .clk ( clk ), .rnd ({Fresh[1643], Fresh[1642]}), .outt ({new_AGEMA_signal_1824, n2212}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2316 ( .ina ({new_AGEMA_signal_1608, n2148}), .inb ({new_AGEMA_signal_1806, n2147}), .clk ( clk ), .rnd ({Fresh[1645], Fresh[1644]}), .outt ({new_AGEMA_signal_1825, n2149}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2366 ( .ina ({new_AGEMA_signal_1808, n2199}), .inb ({new_AGEMA_signal_1740, n2198}), .clk ( clk ), .rnd ({Fresh[1647], Fresh[1646]}), .outt ({new_AGEMA_signal_1826, n2206}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2421 ( .ina ({new_AGEMA_signal_1781, n2258}), .inb ({new_AGEMA_signal_1809, n2257}), .clk ( clk ), .rnd ({Fresh[1649], Fresh[1648]}), .outt ({new_AGEMA_signal_1827, n2310}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2447 ( .ina ({new_AGEMA_signal_1810, n2281}), .inb ({new_AGEMA_signal_1526, n2280}), .clk ( clk ), .rnd ({Fresh[1651], Fresh[1650]}), .outt ({new_AGEMA_signal_1828, n2308}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2476 ( .ina ({new_AGEMA_signal_1621, n2306}), .inb ({new_AGEMA_signal_1811, n2305}), .clk ( clk ), .rnd ({Fresh[1653], Fresh[1652]}), .outt ({new_AGEMA_signal_1829, n2307}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2533 ( .ina ({new_AGEMA_signal_970, n2719}), .inb ({new_AGEMA_signal_1812, n2368}), .clk ( clk ), .rnd ({Fresh[1655], Fresh[1654]}), .outt ({new_AGEMA_signal_1830, n2370}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2611 ( .ina ({new_AGEMA_signal_1814, n2457}), .inb ({new_AGEMA_signal_1637, n2456}), .clk ( clk ), .rnd ({Fresh[1657], Fresh[1656]}), .outt ({new_AGEMA_signal_1831, n2530}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2660 ( .ina ({new_AGEMA_signal_1754, n2514}), .inb ({new_AGEMA_signal_1815, n2513}), .clk ( clk ), .rnd ({Fresh[1659], Fresh[1658]}), .outt ({new_AGEMA_signal_1832, n2515}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2718 ( .ina ({new_AGEMA_signal_1760, n2593}), .inb ({new_AGEMA_signal_1816, n2592}), .clk ( clk ), .rnd ({Fresh[1661], Fresh[1660]}), .outt ({new_AGEMA_signal_1833, n2639}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2749 ( .ina ({new_AGEMA_signal_1793, n2637}), .inb ({new_AGEMA_signal_1763, n2636}), .clk ( clk ), .rnd ({Fresh[1663], Fresh[1662]}), .outt ({new_AGEMA_signal_1817, n2638}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2788 ( .ina ({new_AGEMA_signal_1656, n2706}), .inb ({new_AGEMA_signal_1819, n2705}), .clk ( clk ), .rnd ({Fresh[1665], Fresh[1664]}), .outt ({new_AGEMA_signal_1834, n2832}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2842 ( .ina ({new_AGEMA_signal_1766, n2806}), .inb ({new_AGEMA_signal_1796, n2805}), .clk ( clk ), .rnd ({Fresh[1667], Fresh[1666]}), .outt ({new_AGEMA_signal_1820, n2807}) ) ;

    /* cells in depth 21 */

    /* cells in depth 22 */
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2129 ( .ina ({new_AGEMA_signal_1821, n2000}), .inb ({new_AGEMA_signal_1671, n1999}), .clk ( clk ), .rnd ({Fresh[1669], Fresh[1668]}), .outt ({new_AGEMA_signal_1836, n2001}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2267 ( .ina ({new_AGEMA_signal_1823, n2107}), .inb ({new_AGEMA_signal_1357, n2106}), .clk ( clk ), .rnd ({Fresh[1671], Fresh[1670]}), .outt ({new_AGEMA_signal_1837, n2108}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2317 ( .ina ({new_AGEMA_signal_1197, n2150}), .inb ({new_AGEMA_signal_1825, n2149}), .clk ( clk ), .rnd ({Fresh[1673], Fresh[1672]}), .outt ({new_AGEMA_signal_1838, n2153}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2374 ( .ina ({new_AGEMA_signal_1826, n2206}), .inb ({new_AGEMA_signal_1741, n2205}), .clk ( clk ), .rnd ({Fresh[1675], Fresh[1674]}), .outt ({new_AGEMA_signal_1839, n2207}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2477 ( .ina ({new_AGEMA_signal_1828, n2308}), .inb ({new_AGEMA_signal_1829, n2307}), .clk ( clk ), .rnd ({Fresh[1677], Fresh[1676]}), .outt ({new_AGEMA_signal_1840, n2309}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2535 ( .ina ({new_AGEMA_signal_1830, n2370}), .inb ({new_AGEMA_signal_1540, n2369}), .clk ( clk ), .rnd ({Fresh[1679], Fresh[1678]}), .outt ({new_AGEMA_signal_1841, n2373}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2661 ( .ina ({new_AGEMA_signal_1704, n2516}), .inb ({new_AGEMA_signal_1832, n2515}), .clk ( clk ), .rnd ({Fresh[1681], Fresh[1680]}), .outt ({new_AGEMA_signal_1842, n2528}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2750 ( .ina ({new_AGEMA_signal_1833, n2639}), .inb ({new_AGEMA_signal_1817, n2638}), .clk ( clk ), .rnd ({Fresh[1683], Fresh[1682]}), .outt ({new_AGEMA_signal_1843, n2669}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2843 ( .ina ({new_AGEMA_signal_1719, n2808}), .inb ({new_AGEMA_signal_1820, n2807}), .clk ( clk ), .rnd ({Fresh[1685], Fresh[1684]}), .outt ({new_AGEMA_signal_1835, n2830}) ) ;

    /* cells in depth 23 */

    /* cells in depth 24 */
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2130 ( .ina ({new_AGEMA_signal_1798, n2002}), .inb ({new_AGEMA_signal_1836, n2001}), .clk ( clk ), .rnd ({Fresh[1687], Fresh[1686]}), .outt ({new_AGEMA_signal_1845, n2017}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2268 ( .ina ({new_AGEMA_signal_1822, n2109}), .inb ({new_AGEMA_signal_1837, n2108}), .clk ( clk ), .rnd ({Fresh[1689], Fresh[1688]}), .outt ({new_AGEMA_signal_1846, n2110}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2319 ( .ina ({new_AGEMA_signal_1838, n2153}), .inb ({new_AGEMA_signal_1364, n2152}), .clk ( clk ), .rnd ({Fresh[1691], Fresh[1690]}), .outt ({new_AGEMA_signal_1847, n2154}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2375 ( .ina ({new_AGEMA_signal_1807, n2208}), .inb ({new_AGEMA_signal_1839, n2207}), .clk ( clk ), .rnd ({Fresh[1693], Fresh[1692]}), .outt ({new_AGEMA_signal_1848, n2209}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2478 ( .ina ({new_AGEMA_signal_1827, n2310}), .inb ({new_AGEMA_signal_1840, n2309}), .clk ( clk ), .rnd ({Fresh[1695], Fresh[1694]}), .outt ({new_AGEMA_signal_1849, n2311}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2537 ( .ina ({new_AGEMA_signal_1841, n2373}), .inb ({new_AGEMA_signal_1404, n2372}), .clk ( clk ), .rnd ({Fresh[1697], Fresh[1696]}), .outt ({new_AGEMA_signal_1850, n2374}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2672 ( .ina ({new_AGEMA_signal_1842, n2528}), .inb ({new_AGEMA_signal_1758, n2527}), .clk ( clk ), .rnd ({Fresh[1699], Fresh[1698]}), .outt ({new_AGEMA_signal_1851, n2529}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2768 ( .ina ({new_AGEMA_signal_1843, n2669}), .inb ({new_AGEMA_signal_1818, n2668}), .clk ( clk ), .rnd ({Fresh[1701], Fresh[1700]}), .outt ({new_AGEMA_signal_1852, n2670}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2854 ( .ina ({new_AGEMA_signal_1835, n2830}), .inb ({new_AGEMA_signal_1768, n2829}), .clk ( clk ), .rnd ({Fresh[1703], Fresh[1702]}), .outt ({new_AGEMA_signal_1844, n2831}) ) ;

    /* cells in depth 25 */

    /* cells in depth 26 */
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2155 ( .ina ({new_AGEMA_signal_1845, n2017}), .inb ({new_AGEMA_signal_1800, n2016}), .clk ( clk ), .rnd ({Fresh[1705], Fresh[1704]}), .outt ({new_AGEMA_signal_1854, n2018}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2269 ( .ina ({new_AGEMA_signal_1802, n2111}), .inb ({new_AGEMA_signal_1846, n2110}), .clk ( clk ), .rnd ({Fresh[1707], Fresh[1706]}), .outt ({new_AGEMA_signal_1855, n2112}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2320 ( .ina ({new_AGEMA_signal_1359, n2155}), .inb ({new_AGEMA_signal_1847, n2154}), .clk ( clk ), .rnd ({Fresh[1709], Fresh[1708]}), .outt ({new_AGEMA_signal_1856, n2210}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2479 ( .ina ({new_AGEMA_signal_1742, n2312}), .inb ({new_AGEMA_signal_1849, n2311}), .clk ( clk ), .rnd ({Fresh[1711], Fresh[1710]}), .outt ({new_AGEMA_signal_1857, N470}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2538 ( .ina ({new_AGEMA_signal_1241, n2375}), .inb ({new_AGEMA_signal_1850, n2374}), .clk ( clk ), .rnd ({Fresh[1713], Fresh[1712]}), .outt ({new_AGEMA_signal_1858, n2378}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2673 ( .ina ({new_AGEMA_signal_1831, n2530}), .inb ({new_AGEMA_signal_1851, n2529}), .clk ( clk ), .rnd ({Fresh[1715], Fresh[1714]}), .outt ({new_AGEMA_signal_1859, N639}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2769 ( .ina ({new_AGEMA_signal_1791, n2671}), .inb ({new_AGEMA_signal_1852, n2670}), .clk ( clk ), .rnd ({Fresh[1717], Fresh[1716]}), .outt ({new_AGEMA_signal_1860, N723}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2855 ( .ina ({new_AGEMA_signal_1834, n2832}), .inb ({new_AGEMA_signal_1844, n2831}), .clk ( clk ), .rnd ({Fresh[1719], Fresh[1718]}), .outt ({new_AGEMA_signal_1853, N789}) ) ;

    /* cells in depth 27 */

    /* cells in depth 28 */
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2156 ( .ina ({new_AGEMA_signal_1797, n2019}), .inb ({new_AGEMA_signal_1854, n2018}), .clk ( clk ), .rnd ({Fresh[1721], Fresh[1720]}), .outt ({new_AGEMA_signal_1861, N169}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2270 ( .ina ({new_AGEMA_signal_1801, n2113}), .inb ({new_AGEMA_signal_1855, n2112}), .clk ( clk ), .rnd ({Fresh[1723], Fresh[1722]}), .outt ({new_AGEMA_signal_1862, N277}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2376 ( .ina ({new_AGEMA_signal_1856, n2210}), .inb ({new_AGEMA_signal_1848, n2209}), .clk ( clk ), .rnd ({Fresh[1725], Fresh[1724]}), .outt ({new_AGEMA_signal_1863, n2211}) ) ;
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2540 ( .ina ({new_AGEMA_signal_1858, n2378}), .inb ({new_AGEMA_signal_1405, n2377}), .clk ( clk ), .rnd ({Fresh[1727], Fresh[1726]}), .outt ({new_AGEMA_signal_1864, n2379}) ) ;

    /* cells in depth 29 */

    /* cells in depth 30 */
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2377 ( .ina ({new_AGEMA_signal_1824, n2212}), .inb ({new_AGEMA_signal_1863, n2211}), .clk ( clk ), .rnd ({Fresh[1729], Fresh[1728]}), .outt ({new_AGEMA_signal_1865, N379}) ) ;
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2541 ( .ina ({new_AGEMA_signal_1786, n2380}), .inb ({new_AGEMA_signal_1864, n2379}), .clk ( clk ), .rnd ({Fresh[1731], Fresh[1730]}), .outt ({new_AGEMA_signal_1866, n2381}) ) ;

    /* cells in depth 31 */

    /* cells in depth 32 */
    nor_HPC1 #(.security_order(1), .pipeline(0)) U2542 ( .ina ({new_AGEMA_signal_1785, n2382}), .inb ({new_AGEMA_signal_1866, n2381}), .clk ( clk ), .rnd ({Fresh[1733], Fresh[1732]}), .outt ({new_AGEMA_signal_1867, n2427}) ) ;

    /* cells in depth 33 */

    /* cells in depth 34 */
    nand_HPC1 #(.security_order(1), .pipeline(0)) U2584 ( .ina ({new_AGEMA_signal_1867, n2427}), .inb ({new_AGEMA_signal_1813, n2426}), .clk ( clk ), .rnd ({Fresh[1735], Fresh[1734]}), .outt ({new_AGEMA_signal_1868, N563}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) SO_reg_7_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1861, N169}), .Q ({SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) SO_reg_6_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1862, N277}), .Q ({SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) SO_reg_5_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1865, N379}), .Q ({SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) SO_reg_4_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1857, N470}), .Q ({SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) SO_reg_3_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1868, N563}), .Q ({SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) SO_reg_2_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1859, N639}), .Q ({SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) SO_reg_1_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1860, N723}), .Q ({SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) SO_reg_0_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1853, N789}), .Q ({SO_s1[0], SO_s0[0]}) ) ;
endmodule
