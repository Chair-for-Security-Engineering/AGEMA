
module SkinnyTop_HPC2_ClockGating_d2 ( Plaintext_s0, Key_s0, clk, rst, Key_s1, 
        Key_s2, Plaintext_s1, Plaintext_s2, Fresh, Ciphertext_s0, done, 
        Ciphertext_s1, Ciphertext_s2, Synch );
  input [63:0] Plaintext_s0;
  input [63:0] Key_s0;
  input [63:0] Key_s1;
  input [63:0] Key_s2;
  input [63:0] Plaintext_s1;
  input [63:0] Plaintext_s2;
  input [191:0] Fresh;
  output [63:0] Ciphertext_s0;
  output [63:0] Ciphertext_s1;
  output [63:0] Ciphertext_s2;
  input clk, rst;
  output done, Synch;
  wire   SubCellInst_SboxInst_0_n3, new_AGEMA_signal_1171,
         new_AGEMA_signal_1170, SubCellInst_SboxInst_0_XX_1_,
         new_AGEMA_signal_1175, new_AGEMA_signal_1174,
         SubCellInst_SboxInst_0_XX_2_, new_AGEMA_signal_1743,
         new_AGEMA_signal_1742, SubCellInst_SboxInst_0_Q0,
         new_AGEMA_signal_1745, new_AGEMA_signal_1744,
         SubCellInst_SboxInst_0_Q1, new_AGEMA_signal_1747,
         new_AGEMA_signal_1746, SubCellInst_SboxInst_0_Q4,
         new_AGEMA_signal_1749, new_AGEMA_signal_1748,
         SubCellInst_SboxInst_0_Q6, new_AGEMA_signal_1937,
         new_AGEMA_signal_1936, SubCellInst_SboxInst_0_L1,
         new_AGEMA_signal_1751, new_AGEMA_signal_1750,
         SubCellInst_SboxInst_0_L2, SubCellInst_SboxInst_1_n3,
         new_AGEMA_signal_1183, new_AGEMA_signal_1182,
         SubCellInst_SboxInst_1_XX_1_, new_AGEMA_signal_1187,
         new_AGEMA_signal_1186, SubCellInst_SboxInst_1_XX_2_,
         new_AGEMA_signal_1755, new_AGEMA_signal_1754,
         SubCellInst_SboxInst_1_Q0, new_AGEMA_signal_1757,
         new_AGEMA_signal_1756, SubCellInst_SboxInst_1_Q1,
         new_AGEMA_signal_1759, new_AGEMA_signal_1758,
         SubCellInst_SboxInst_1_Q4, new_AGEMA_signal_1761,
         new_AGEMA_signal_1760, SubCellInst_SboxInst_1_Q6,
         new_AGEMA_signal_1943, new_AGEMA_signal_1942,
         SubCellInst_SboxInst_1_L1, new_AGEMA_signal_1763,
         new_AGEMA_signal_1762, SubCellInst_SboxInst_1_L2,
         SubCellInst_SboxInst_2_n3, new_AGEMA_signal_1195,
         new_AGEMA_signal_1194, SubCellInst_SboxInst_2_XX_1_,
         new_AGEMA_signal_1199, new_AGEMA_signal_1198,
         SubCellInst_SboxInst_2_XX_2_, new_AGEMA_signal_1767,
         new_AGEMA_signal_1766, SubCellInst_SboxInst_2_Q0,
         new_AGEMA_signal_1769, new_AGEMA_signal_1768,
         SubCellInst_SboxInst_2_Q1, new_AGEMA_signal_1771,
         new_AGEMA_signal_1770, SubCellInst_SboxInst_2_Q4,
         new_AGEMA_signal_1773, new_AGEMA_signal_1772,
         SubCellInst_SboxInst_2_Q6, new_AGEMA_signal_1949,
         new_AGEMA_signal_1948, SubCellInst_SboxInst_2_L1,
         new_AGEMA_signal_1775, new_AGEMA_signal_1774,
         SubCellInst_SboxInst_2_L2, SubCellInst_SboxInst_3_n3,
         new_AGEMA_signal_1207, new_AGEMA_signal_1206,
         SubCellInst_SboxInst_3_XX_1_, new_AGEMA_signal_1211,
         new_AGEMA_signal_1210, SubCellInst_SboxInst_3_XX_2_,
         new_AGEMA_signal_1779, new_AGEMA_signal_1778,
         SubCellInst_SboxInst_3_Q0, new_AGEMA_signal_1781,
         new_AGEMA_signal_1780, SubCellInst_SboxInst_3_Q1,
         new_AGEMA_signal_1783, new_AGEMA_signal_1782,
         SubCellInst_SboxInst_3_Q4, new_AGEMA_signal_1785,
         new_AGEMA_signal_1784, SubCellInst_SboxInst_3_Q6,
         new_AGEMA_signal_1955, new_AGEMA_signal_1954,
         SubCellInst_SboxInst_3_L1, new_AGEMA_signal_1787,
         new_AGEMA_signal_1786, SubCellInst_SboxInst_3_L2,
         SubCellInst_SboxInst_4_n3, new_AGEMA_signal_1219,
         new_AGEMA_signal_1218, SubCellInst_SboxInst_4_XX_1_,
         new_AGEMA_signal_1223, new_AGEMA_signal_1222,
         SubCellInst_SboxInst_4_XX_2_, new_AGEMA_signal_1791,
         new_AGEMA_signal_1790, SubCellInst_SboxInst_4_Q0,
         new_AGEMA_signal_1793, new_AGEMA_signal_1792,
         SubCellInst_SboxInst_4_Q1, new_AGEMA_signal_1795,
         new_AGEMA_signal_1794, SubCellInst_SboxInst_4_Q4,
         new_AGEMA_signal_1797, new_AGEMA_signal_1796,
         SubCellInst_SboxInst_4_Q6, new_AGEMA_signal_1961,
         new_AGEMA_signal_1960, SubCellInst_SboxInst_4_L1,
         new_AGEMA_signal_1799, new_AGEMA_signal_1798,
         SubCellInst_SboxInst_4_L2, SubCellInst_SboxInst_5_n3,
         new_AGEMA_signal_1231, new_AGEMA_signal_1230,
         SubCellInst_SboxInst_5_XX_1_, new_AGEMA_signal_1235,
         new_AGEMA_signal_1234, SubCellInst_SboxInst_5_XX_2_,
         new_AGEMA_signal_1803, new_AGEMA_signal_1802,
         SubCellInst_SboxInst_5_Q0, new_AGEMA_signal_1805,
         new_AGEMA_signal_1804, SubCellInst_SboxInst_5_Q1,
         new_AGEMA_signal_1807, new_AGEMA_signal_1806,
         SubCellInst_SboxInst_5_Q4, new_AGEMA_signal_1809,
         new_AGEMA_signal_1808, SubCellInst_SboxInst_5_Q6,
         new_AGEMA_signal_1967, new_AGEMA_signal_1966,
         SubCellInst_SboxInst_5_L1, new_AGEMA_signal_1811,
         new_AGEMA_signal_1810, SubCellInst_SboxInst_5_L2,
         SubCellInst_SboxInst_6_n3, new_AGEMA_signal_1243,
         new_AGEMA_signal_1242, SubCellInst_SboxInst_6_XX_1_,
         new_AGEMA_signal_1247, new_AGEMA_signal_1246,
         SubCellInst_SboxInst_6_XX_2_, new_AGEMA_signal_1815,
         new_AGEMA_signal_1814, SubCellInst_SboxInst_6_Q0,
         new_AGEMA_signal_1817, new_AGEMA_signal_1816,
         SubCellInst_SboxInst_6_Q1, new_AGEMA_signal_1819,
         new_AGEMA_signal_1818, SubCellInst_SboxInst_6_Q4,
         new_AGEMA_signal_1821, new_AGEMA_signal_1820,
         SubCellInst_SboxInst_6_Q6, new_AGEMA_signal_1973,
         new_AGEMA_signal_1972, SubCellInst_SboxInst_6_L1,
         new_AGEMA_signal_1823, new_AGEMA_signal_1822,
         SubCellInst_SboxInst_6_L2, SubCellInst_SboxInst_7_n3,
         new_AGEMA_signal_1255, new_AGEMA_signal_1254,
         SubCellInst_SboxInst_7_XX_1_, new_AGEMA_signal_1259,
         new_AGEMA_signal_1258, SubCellInst_SboxInst_7_XX_2_,
         new_AGEMA_signal_1827, new_AGEMA_signal_1826,
         SubCellInst_SboxInst_7_Q0, new_AGEMA_signal_1829,
         new_AGEMA_signal_1828, SubCellInst_SboxInst_7_Q1,
         new_AGEMA_signal_1831, new_AGEMA_signal_1830,
         SubCellInst_SboxInst_7_Q4, new_AGEMA_signal_1833,
         new_AGEMA_signal_1832, SubCellInst_SboxInst_7_Q6,
         new_AGEMA_signal_1979, new_AGEMA_signal_1978,
         SubCellInst_SboxInst_7_L1, new_AGEMA_signal_1835,
         new_AGEMA_signal_1834, SubCellInst_SboxInst_7_L2,
         SubCellInst_SboxInst_8_n3, new_AGEMA_signal_1267,
         new_AGEMA_signal_1266, SubCellInst_SboxInst_8_XX_1_,
         new_AGEMA_signal_1271, new_AGEMA_signal_1270,
         SubCellInst_SboxInst_8_XX_2_, new_AGEMA_signal_1839,
         new_AGEMA_signal_1838, SubCellInst_SboxInst_8_Q0,
         new_AGEMA_signal_1841, new_AGEMA_signal_1840,
         SubCellInst_SboxInst_8_Q1, new_AGEMA_signal_1843,
         new_AGEMA_signal_1842, SubCellInst_SboxInst_8_Q4,
         new_AGEMA_signal_1845, new_AGEMA_signal_1844,
         SubCellInst_SboxInst_8_Q6, new_AGEMA_signal_1985,
         new_AGEMA_signal_1984, SubCellInst_SboxInst_8_L1,
         new_AGEMA_signal_1847, new_AGEMA_signal_1846,
         SubCellInst_SboxInst_8_L2, SubCellInst_SboxInst_9_n3,
         new_AGEMA_signal_1279, new_AGEMA_signal_1278,
         SubCellInst_SboxInst_9_XX_1_, new_AGEMA_signal_1283,
         new_AGEMA_signal_1282, SubCellInst_SboxInst_9_XX_2_,
         new_AGEMA_signal_1851, new_AGEMA_signal_1850,
         SubCellInst_SboxInst_9_Q0, new_AGEMA_signal_1853,
         new_AGEMA_signal_1852, SubCellInst_SboxInst_9_Q1,
         new_AGEMA_signal_1855, new_AGEMA_signal_1854,
         SubCellInst_SboxInst_9_Q4, new_AGEMA_signal_1857,
         new_AGEMA_signal_1856, SubCellInst_SboxInst_9_Q6,
         new_AGEMA_signal_1991, new_AGEMA_signal_1990,
         SubCellInst_SboxInst_9_L1, new_AGEMA_signal_1859,
         new_AGEMA_signal_1858, SubCellInst_SboxInst_9_L2,
         SubCellInst_SboxInst_10_n3, new_AGEMA_signal_1291,
         new_AGEMA_signal_1290, SubCellInst_SboxInst_10_XX_1_,
         new_AGEMA_signal_1295, new_AGEMA_signal_1294,
         SubCellInst_SboxInst_10_XX_2_, new_AGEMA_signal_1863,
         new_AGEMA_signal_1862, SubCellInst_SboxInst_10_Q0,
         new_AGEMA_signal_1865, new_AGEMA_signal_1864,
         SubCellInst_SboxInst_10_Q1, new_AGEMA_signal_1867,
         new_AGEMA_signal_1866, SubCellInst_SboxInst_10_Q4,
         new_AGEMA_signal_1869, new_AGEMA_signal_1868,
         SubCellInst_SboxInst_10_Q6, new_AGEMA_signal_1997,
         new_AGEMA_signal_1996, SubCellInst_SboxInst_10_L1,
         new_AGEMA_signal_1871, new_AGEMA_signal_1870,
         SubCellInst_SboxInst_10_L2, SubCellInst_SboxInst_11_n3,
         new_AGEMA_signal_1303, new_AGEMA_signal_1302,
         SubCellInst_SboxInst_11_XX_1_, new_AGEMA_signal_1307,
         new_AGEMA_signal_1306, SubCellInst_SboxInst_11_XX_2_,
         new_AGEMA_signal_1875, new_AGEMA_signal_1874,
         SubCellInst_SboxInst_11_Q0, new_AGEMA_signal_1877,
         new_AGEMA_signal_1876, SubCellInst_SboxInst_11_Q1,
         new_AGEMA_signal_1879, new_AGEMA_signal_1878,
         SubCellInst_SboxInst_11_Q4, new_AGEMA_signal_1881,
         new_AGEMA_signal_1880, SubCellInst_SboxInst_11_Q6,
         new_AGEMA_signal_2003, new_AGEMA_signal_2002,
         SubCellInst_SboxInst_11_L1, new_AGEMA_signal_1883,
         new_AGEMA_signal_1882, SubCellInst_SboxInst_11_L2,
         SubCellInst_SboxInst_12_n3, new_AGEMA_signal_1315,
         new_AGEMA_signal_1314, SubCellInst_SboxInst_12_XX_1_,
         new_AGEMA_signal_1319, new_AGEMA_signal_1318,
         SubCellInst_SboxInst_12_XX_2_, new_AGEMA_signal_1887,
         new_AGEMA_signal_1886, SubCellInst_SboxInst_12_Q0,
         new_AGEMA_signal_1889, new_AGEMA_signal_1888,
         SubCellInst_SboxInst_12_Q1, new_AGEMA_signal_1891,
         new_AGEMA_signal_1890, SubCellInst_SboxInst_12_Q4,
         new_AGEMA_signal_1893, new_AGEMA_signal_1892,
         SubCellInst_SboxInst_12_Q6, new_AGEMA_signal_2009,
         new_AGEMA_signal_2008, SubCellInst_SboxInst_12_L1,
         new_AGEMA_signal_1895, new_AGEMA_signal_1894,
         SubCellInst_SboxInst_12_L2, SubCellInst_SboxInst_13_n3,
         new_AGEMA_signal_1327, new_AGEMA_signal_1326,
         SubCellInst_SboxInst_13_XX_1_, new_AGEMA_signal_1331,
         new_AGEMA_signal_1330, SubCellInst_SboxInst_13_XX_2_,
         new_AGEMA_signal_1899, new_AGEMA_signal_1898,
         SubCellInst_SboxInst_13_Q0, new_AGEMA_signal_1901,
         new_AGEMA_signal_1900, SubCellInst_SboxInst_13_Q1,
         new_AGEMA_signal_1903, new_AGEMA_signal_1902,
         SubCellInst_SboxInst_13_Q4, new_AGEMA_signal_1905,
         new_AGEMA_signal_1904, SubCellInst_SboxInst_13_Q6,
         new_AGEMA_signal_2015, new_AGEMA_signal_2014,
         SubCellInst_SboxInst_13_L1, new_AGEMA_signal_1907,
         new_AGEMA_signal_1906, SubCellInst_SboxInst_13_L2,
         SubCellInst_SboxInst_14_n3, new_AGEMA_signal_1339,
         new_AGEMA_signal_1338, SubCellInst_SboxInst_14_XX_1_,
         new_AGEMA_signal_1343, new_AGEMA_signal_1342,
         SubCellInst_SboxInst_14_XX_2_, new_AGEMA_signal_1911,
         new_AGEMA_signal_1910, SubCellInst_SboxInst_14_Q0,
         new_AGEMA_signal_1913, new_AGEMA_signal_1912,
         SubCellInst_SboxInst_14_Q1, new_AGEMA_signal_1915,
         new_AGEMA_signal_1914, SubCellInst_SboxInst_14_Q4,
         new_AGEMA_signal_1917, new_AGEMA_signal_1916,
         SubCellInst_SboxInst_14_Q6, new_AGEMA_signal_2021,
         new_AGEMA_signal_2020, SubCellInst_SboxInst_14_L1,
         new_AGEMA_signal_1919, new_AGEMA_signal_1918,
         SubCellInst_SboxInst_14_L2, SubCellInst_SboxInst_15_n3,
         new_AGEMA_signal_1351, new_AGEMA_signal_1350,
         SubCellInst_SboxInst_15_XX_1_, new_AGEMA_signal_1355,
         new_AGEMA_signal_1354, SubCellInst_SboxInst_15_XX_2_,
         new_AGEMA_signal_1923, new_AGEMA_signal_1922,
         SubCellInst_SboxInst_15_Q0, new_AGEMA_signal_1925,
         new_AGEMA_signal_1924, SubCellInst_SboxInst_15_Q1,
         new_AGEMA_signal_1927, new_AGEMA_signal_1926,
         SubCellInst_SboxInst_15_Q4, new_AGEMA_signal_1929,
         new_AGEMA_signal_1928, SubCellInst_SboxInst_15_Q6,
         new_AGEMA_signal_2027, new_AGEMA_signal_2026,
         SubCellInst_SboxInst_15_L1, new_AGEMA_signal_1931,
         new_AGEMA_signal_1930, SubCellInst_SboxInst_15_L2,
         new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1357,
         new_AGEMA_signal_1356, new_AGEMA_signal_1367, new_AGEMA_signal_1366,
         new_AGEMA_signal_1363, new_AGEMA_signal_1362, new_AGEMA_signal_1373,
         new_AGEMA_signal_1372, new_AGEMA_signal_1369, new_AGEMA_signal_1368,
         new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1375,
         new_AGEMA_signal_1374, new_AGEMA_signal_1385, new_AGEMA_signal_1384,
         new_AGEMA_signal_1381, new_AGEMA_signal_1380, new_AGEMA_signal_1391,
         new_AGEMA_signal_1390, new_AGEMA_signal_1387, new_AGEMA_signal_1386,
         new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1393,
         new_AGEMA_signal_1392, new_AGEMA_signal_1403, new_AGEMA_signal_1402,
         new_AGEMA_signal_1399, new_AGEMA_signal_1398, new_AGEMA_signal_1409,
         new_AGEMA_signal_1408, new_AGEMA_signal_1405, new_AGEMA_signal_1404,
         new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1411,
         new_AGEMA_signal_1410, new_AGEMA_signal_1421, new_AGEMA_signal_1420,
         new_AGEMA_signal_1417, new_AGEMA_signal_1416, new_AGEMA_signal_1427,
         new_AGEMA_signal_1426, new_AGEMA_signal_1423, new_AGEMA_signal_1422,
         new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1429,
         new_AGEMA_signal_1428, new_AGEMA_signal_1439, new_AGEMA_signal_1438,
         new_AGEMA_signal_1435, new_AGEMA_signal_1434, new_AGEMA_signal_1445,
         new_AGEMA_signal_1444, new_AGEMA_signal_1441, new_AGEMA_signal_1440,
         new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1447,
         new_AGEMA_signal_1446, new_AGEMA_signal_1457, new_AGEMA_signal_1456,
         new_AGEMA_signal_1453, new_AGEMA_signal_1452, new_AGEMA_signal_1463,
         new_AGEMA_signal_1462, new_AGEMA_signal_1459, new_AGEMA_signal_1458,
         new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1465,
         new_AGEMA_signal_1464, new_AGEMA_signal_1475, new_AGEMA_signal_1474,
         new_AGEMA_signal_1471, new_AGEMA_signal_1470, new_AGEMA_signal_1481,
         new_AGEMA_signal_1480, new_AGEMA_signal_1477, new_AGEMA_signal_1476,
         new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1483,
         new_AGEMA_signal_1482, new_AGEMA_signal_1493, new_AGEMA_signal_1492,
         new_AGEMA_signal_1489, new_AGEMA_signal_1488, new_AGEMA_signal_1499,
         new_AGEMA_signal_1498, new_AGEMA_signal_1495, new_AGEMA_signal_1494,
         new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1501,
         new_AGEMA_signal_1500, new_AGEMA_signal_1511, new_AGEMA_signal_1510,
         new_AGEMA_signal_1507, new_AGEMA_signal_1506, new_AGEMA_signal_1517,
         new_AGEMA_signal_1516, new_AGEMA_signal_1513, new_AGEMA_signal_1512,
         new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1519,
         new_AGEMA_signal_1518, new_AGEMA_signal_1529, new_AGEMA_signal_1528,
         new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1535,
         new_AGEMA_signal_1534, new_AGEMA_signal_1531, new_AGEMA_signal_1530,
         new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1537,
         new_AGEMA_signal_1536, new_AGEMA_signal_1547, new_AGEMA_signal_1546,
         new_AGEMA_signal_1543, new_AGEMA_signal_1542, new_AGEMA_signal_1553,
         new_AGEMA_signal_1552, new_AGEMA_signal_1549, new_AGEMA_signal_1548,
         new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1555,
         new_AGEMA_signal_1554, new_AGEMA_signal_1565, new_AGEMA_signal_1564,
         new_AGEMA_signal_1561, new_AGEMA_signal_1560, new_AGEMA_signal_1571,
         new_AGEMA_signal_1570, new_AGEMA_signal_1567, new_AGEMA_signal_1566,
         new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1573,
         new_AGEMA_signal_1572, new_AGEMA_signal_1583, new_AGEMA_signal_1582,
         new_AGEMA_signal_1579, new_AGEMA_signal_1578, new_AGEMA_signal_1589,
         new_AGEMA_signal_1588, new_AGEMA_signal_1585, new_AGEMA_signal_1584,
         new_AGEMA_signal_1595, new_AGEMA_signal_1594, new_AGEMA_signal_1591,
         new_AGEMA_signal_1590, new_AGEMA_signal_1601, new_AGEMA_signal_1600,
         new_AGEMA_signal_1597, new_AGEMA_signal_1596, new_AGEMA_signal_1607,
         new_AGEMA_signal_1606, new_AGEMA_signal_1603, new_AGEMA_signal_1602,
         new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1609,
         new_AGEMA_signal_1608, new_AGEMA_signal_1619, new_AGEMA_signal_1618,
         new_AGEMA_signal_1615, new_AGEMA_signal_1614, new_AGEMA_signal_1625,
         new_AGEMA_signal_1624, new_AGEMA_signal_1621, new_AGEMA_signal_1620,
         new_AGEMA_signal_1631, new_AGEMA_signal_1630, new_AGEMA_signal_1627,
         new_AGEMA_signal_1626, new_AGEMA_signal_1637, new_AGEMA_signal_1636,
         new_AGEMA_signal_1633, new_AGEMA_signal_1632, new_AGEMA_signal_1643,
         new_AGEMA_signal_1642, new_AGEMA_signal_1639, new_AGEMA_signal_1638,
         new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1645,
         new_AGEMA_signal_1644, new_AGEMA_signal_1655, new_AGEMA_signal_1654,
         new_AGEMA_signal_1651, new_AGEMA_signal_1650, new_AGEMA_signal_1661,
         new_AGEMA_signal_1660, new_AGEMA_signal_1657, new_AGEMA_signal_1656,
         new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1663,
         new_AGEMA_signal_1662, new_AGEMA_signal_1673, new_AGEMA_signal_1672,
         new_AGEMA_signal_1669, new_AGEMA_signal_1668, new_AGEMA_signal_1679,
         new_AGEMA_signal_1678, new_AGEMA_signal_1675, new_AGEMA_signal_1674,
         new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1681,
         new_AGEMA_signal_1680, new_AGEMA_signal_1691, new_AGEMA_signal_1690,
         new_AGEMA_signal_1687, new_AGEMA_signal_1686, new_AGEMA_signal_1697,
         new_AGEMA_signal_1696, new_AGEMA_signal_1693, new_AGEMA_signal_1692,
         new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1699,
         new_AGEMA_signal_1698, new_AGEMA_signal_1709, new_AGEMA_signal_1708,
         new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1715,
         new_AGEMA_signal_1714, new_AGEMA_signal_1711, new_AGEMA_signal_1710,
         new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1717,
         new_AGEMA_signal_1716, new_AGEMA_signal_1727, new_AGEMA_signal_1726,
         new_AGEMA_signal_1723, new_AGEMA_signal_1722, new_AGEMA_signal_1733,
         new_AGEMA_signal_1732, new_AGEMA_signal_1729, new_AGEMA_signal_1728,
         new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1735,
         new_AGEMA_signal_1734, FSM_1, clk_gated, new_AGEMA_signal_2681,
         new_AGEMA_signal_2680, new_AGEMA_signal_2667, new_AGEMA_signal_2666,
         new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2787,
         new_AGEMA_signal_2786, new_AGEMA_signal_2685, new_AGEMA_signal_2684,
         new_AGEMA_signal_2671, new_AGEMA_signal_2670, new_AGEMA_signal_2805,
         new_AGEMA_signal_2804, new_AGEMA_signal_2791, new_AGEMA_signal_2790,
         new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2675,
         new_AGEMA_signal_2674, new_AGEMA_signal_2809, new_AGEMA_signal_2808,
         new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2921,
         new_AGEMA_signal_2920, new_AGEMA_signal_2903, new_AGEMA_signal_2902,
         new_AGEMA_signal_3007, new_AGEMA_signal_3006, new_AGEMA_signal_2991,
         new_AGEMA_signal_2990, new_AGEMA_signal_2693, new_AGEMA_signal_2692,
         new_AGEMA_signal_2655, new_AGEMA_signal_2654, new_AGEMA_signal_2813,
         new_AGEMA_signal_2812, new_AGEMA_signal_2773, new_AGEMA_signal_2772,
         new_AGEMA_signal_2697, new_AGEMA_signal_2696, new_AGEMA_signal_2659,
         new_AGEMA_signal_2658, new_AGEMA_signal_2817, new_AGEMA_signal_2816,
         new_AGEMA_signal_2777, new_AGEMA_signal_2776, new_AGEMA_signal_2933,
         new_AGEMA_signal_2932, new_AGEMA_signal_2883, new_AGEMA_signal_2882,
         new_AGEMA_signal_3019, new_AGEMA_signal_3018, new_AGEMA_signal_2979,
         new_AGEMA_signal_2978, new_AGEMA_signal_2701, new_AGEMA_signal_2700,
         new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2821,
         new_AGEMA_signal_2820, new_AGEMA_signal_2783, new_AGEMA_signal_2782,
         new_AGEMA_signal_2479, new_AGEMA_signal_2478, new_AGEMA_signal_2457,
         new_AGEMA_signal_2456, new_AGEMA_signal_2585, new_AGEMA_signal_2584,
         new_AGEMA_signal_2545, new_AGEMA_signal_2544, new_AGEMA_signal_2483,
         new_AGEMA_signal_2482, new_AGEMA_signal_2461, new_AGEMA_signal_2460,
         new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2549,
         new_AGEMA_signal_2548, new_AGEMA_signal_2487, new_AGEMA_signal_2486,
         new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2593,
         new_AGEMA_signal_2592, new_AGEMA_signal_2553, new_AGEMA_signal_2552,
         new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2633,
         new_AGEMA_signal_2632, new_AGEMA_signal_2837, new_AGEMA_signal_2836,
         new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2721,
         new_AGEMA_signal_2720, new_AGEMA_signal_2639, new_AGEMA_signal_2638,
         new_AGEMA_signal_2841, new_AGEMA_signal_2840, new_AGEMA_signal_2757,
         new_AGEMA_signal_2756, new_AGEMA_signal_2725, new_AGEMA_signal_2724,
         new_AGEMA_signal_2643, new_AGEMA_signal_2642, new_AGEMA_signal_2845,
         new_AGEMA_signal_2844, new_AGEMA_signal_2763, new_AGEMA_signal_2762,
         new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2649,
         new_AGEMA_signal_2648, new_AGEMA_signal_2849, new_AGEMA_signal_2848,
         new_AGEMA_signal_2767, new_AGEMA_signal_2766, new_AGEMA_signal_2957,
         new_AGEMA_signal_2956, new_AGEMA_signal_2871, new_AGEMA_signal_2870,
         new_AGEMA_signal_3043, new_AGEMA_signal_3042, new_AGEMA_signal_2971,
         new_AGEMA_signal_2970, new_AGEMA_signal_2285, new_AGEMA_signal_2284,
         SubCellInst_SboxInst_0_YY_1_, new_AGEMA_signal_2157,
         new_AGEMA_signal_2156, SubCellInst_SboxInst_0_YY_0_,
         new_AGEMA_signal_1933, new_AGEMA_signal_1932,
         SubCellInst_SboxInst_0_T0, new_AGEMA_signal_2029,
         new_AGEMA_signal_2028, SubCellInst_SboxInst_0_Q2,
         new_AGEMA_signal_1935, new_AGEMA_signal_1934,
         SubCellInst_SboxInst_0_T2, new_AGEMA_signal_2031,
         new_AGEMA_signal_2030, SubCellInst_SboxInst_0_Q7,
         new_AGEMA_signal_2033, new_AGEMA_signal_2032,
         SubCellInst_SboxInst_0_L3, new_AGEMA_signal_2289,
         new_AGEMA_signal_2288, SubCellInst_SboxInst_1_YY_1_,
         new_AGEMA_signal_2165, new_AGEMA_signal_2164,
         SubCellInst_SboxInst_1_YY_0_, new_AGEMA_signal_1939,
         new_AGEMA_signal_1938, SubCellInst_SboxInst_1_T0,
         new_AGEMA_signal_2037, new_AGEMA_signal_2036,
         SubCellInst_SboxInst_1_Q2, new_AGEMA_signal_1941,
         new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2,
         new_AGEMA_signal_2039, new_AGEMA_signal_2038,
         SubCellInst_SboxInst_1_Q7, new_AGEMA_signal_2041,
         new_AGEMA_signal_2040, SubCellInst_SboxInst_1_L3,
         new_AGEMA_signal_2293, new_AGEMA_signal_2292,
         SubCellInst_SboxInst_2_YY_1_, new_AGEMA_signal_2173,
         new_AGEMA_signal_2172, SubCellInst_SboxInst_2_YY_0_,
         new_AGEMA_signal_1945, new_AGEMA_signal_1944,
         SubCellInst_SboxInst_2_T0, new_AGEMA_signal_2045,
         new_AGEMA_signal_2044, SubCellInst_SboxInst_2_Q2,
         new_AGEMA_signal_1947, new_AGEMA_signal_1946,
         SubCellInst_SboxInst_2_T2, new_AGEMA_signal_2047,
         new_AGEMA_signal_2046, SubCellInst_SboxInst_2_Q7,
         new_AGEMA_signal_2049, new_AGEMA_signal_2048,
         SubCellInst_SboxInst_2_L3, new_AGEMA_signal_2297,
         new_AGEMA_signal_2296, SubCellInst_SboxInst_3_YY_1_,
         new_AGEMA_signal_2181, new_AGEMA_signal_2180,
         SubCellInst_SboxInst_3_YY_0_, new_AGEMA_signal_1951,
         new_AGEMA_signal_1950, SubCellInst_SboxInst_3_T0,
         new_AGEMA_signal_2053, new_AGEMA_signal_2052,
         SubCellInst_SboxInst_3_Q2, new_AGEMA_signal_1953,
         new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2,
         new_AGEMA_signal_2055, new_AGEMA_signal_2054,
         SubCellInst_SboxInst_3_Q7, new_AGEMA_signal_2057,
         new_AGEMA_signal_2056, SubCellInst_SboxInst_3_L3,
         new_AGEMA_signal_2301, new_AGEMA_signal_2300,
         SubCellInst_SboxInst_4_YY_1_, new_AGEMA_signal_2189,
         new_AGEMA_signal_2188, SubCellInst_SboxInst_4_YY_0_,
         new_AGEMA_signal_1957, new_AGEMA_signal_1956,
         SubCellInst_SboxInst_4_T0, new_AGEMA_signal_2061,
         new_AGEMA_signal_2060, SubCellInst_SboxInst_4_Q2,
         new_AGEMA_signal_1959, new_AGEMA_signal_1958,
         SubCellInst_SboxInst_4_T2, new_AGEMA_signal_2063,
         new_AGEMA_signal_2062, SubCellInst_SboxInst_4_Q7,
         new_AGEMA_signal_2065, new_AGEMA_signal_2064,
         SubCellInst_SboxInst_4_L3, new_AGEMA_signal_2305,
         new_AGEMA_signal_2304, SubCellInst_SboxInst_5_YY_1_,
         new_AGEMA_signal_2197, new_AGEMA_signal_2196,
         SubCellInst_SboxInst_5_YY_0_, new_AGEMA_signal_1963,
         new_AGEMA_signal_1962, SubCellInst_SboxInst_5_T0,
         new_AGEMA_signal_2069, new_AGEMA_signal_2068,
         SubCellInst_SboxInst_5_Q2, new_AGEMA_signal_1965,
         new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2,
         new_AGEMA_signal_2071, new_AGEMA_signal_2070,
         SubCellInst_SboxInst_5_Q7, new_AGEMA_signal_2073,
         new_AGEMA_signal_2072, SubCellInst_SboxInst_5_L3,
         new_AGEMA_signal_2309, new_AGEMA_signal_2308,
         SubCellInst_SboxInst_6_YY_1_, new_AGEMA_signal_2205,
         new_AGEMA_signal_2204, SubCellInst_SboxInst_6_YY_0_,
         new_AGEMA_signal_1969, new_AGEMA_signal_1968,
         SubCellInst_SboxInst_6_T0, new_AGEMA_signal_2077,
         new_AGEMA_signal_2076, SubCellInst_SboxInst_6_Q2,
         new_AGEMA_signal_1971, new_AGEMA_signal_1970,
         SubCellInst_SboxInst_6_T2, new_AGEMA_signal_2079,
         new_AGEMA_signal_2078, SubCellInst_SboxInst_6_Q7,
         new_AGEMA_signal_2081, new_AGEMA_signal_2080,
         SubCellInst_SboxInst_6_L3, new_AGEMA_signal_2313,
         new_AGEMA_signal_2312, SubCellInst_SboxInst_7_YY_1_,
         new_AGEMA_signal_2213, new_AGEMA_signal_2212,
         SubCellInst_SboxInst_7_YY_0_, new_AGEMA_signal_1975,
         new_AGEMA_signal_1974, SubCellInst_SboxInst_7_T0,
         new_AGEMA_signal_2085, new_AGEMA_signal_2084,
         SubCellInst_SboxInst_7_Q2, new_AGEMA_signal_1977,
         new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2,
         new_AGEMA_signal_2087, new_AGEMA_signal_2086,
         SubCellInst_SboxInst_7_Q7, new_AGEMA_signal_2089,
         new_AGEMA_signal_2088, SubCellInst_SboxInst_7_L3,
         new_AGEMA_signal_2317, new_AGEMA_signal_2316,
         SubCellInst_SboxInst_8_YY_1_, new_AGEMA_signal_2221,
         new_AGEMA_signal_2220, SubCellInst_SboxInst_8_YY_0_,
         new_AGEMA_signal_1981, new_AGEMA_signal_1980,
         SubCellInst_SboxInst_8_T0, new_AGEMA_signal_2093,
         new_AGEMA_signal_2092, SubCellInst_SboxInst_8_Q2,
         new_AGEMA_signal_1983, new_AGEMA_signal_1982,
         SubCellInst_SboxInst_8_T2, new_AGEMA_signal_2095,
         new_AGEMA_signal_2094, SubCellInst_SboxInst_8_Q7,
         new_AGEMA_signal_2097, new_AGEMA_signal_2096,
         SubCellInst_SboxInst_8_L3, new_AGEMA_signal_2321,
         new_AGEMA_signal_2320, SubCellInst_SboxInst_9_YY_1_,
         new_AGEMA_signal_2229, new_AGEMA_signal_2228,
         SubCellInst_SboxInst_9_YY_0_, new_AGEMA_signal_1987,
         new_AGEMA_signal_1986, SubCellInst_SboxInst_9_T0,
         new_AGEMA_signal_2101, new_AGEMA_signal_2100,
         SubCellInst_SboxInst_9_Q2, new_AGEMA_signal_1989,
         new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2,
         new_AGEMA_signal_2103, new_AGEMA_signal_2102,
         SubCellInst_SboxInst_9_Q7, new_AGEMA_signal_2105,
         new_AGEMA_signal_2104, SubCellInst_SboxInst_9_L3,
         new_AGEMA_signal_2325, new_AGEMA_signal_2324,
         SubCellInst_SboxInst_10_YY_1_, new_AGEMA_signal_2237,
         new_AGEMA_signal_2236, SubCellInst_SboxInst_10_YY_0_,
         new_AGEMA_signal_1993, new_AGEMA_signal_1992,
         SubCellInst_SboxInst_10_T0, new_AGEMA_signal_2109,
         new_AGEMA_signal_2108, SubCellInst_SboxInst_10_Q2,
         new_AGEMA_signal_1995, new_AGEMA_signal_1994,
         SubCellInst_SboxInst_10_T2, new_AGEMA_signal_2111,
         new_AGEMA_signal_2110, SubCellInst_SboxInst_10_Q7,
         new_AGEMA_signal_2113, new_AGEMA_signal_2112,
         SubCellInst_SboxInst_10_L3, SubCellOutput_47, SubCellOutput_46,
         SubCellOutput_45, SubCellOutput_44, SubCellOutput_29,
         new_AGEMA_signal_2329, new_AGEMA_signal_2328,
         SubCellInst_SboxInst_11_YY_1_, new_AGEMA_signal_2245,
         new_AGEMA_signal_2244, SubCellInst_SboxInst_11_YY_0_,
         new_AGEMA_signal_1999, new_AGEMA_signal_1998,
         SubCellInst_SboxInst_11_T0, new_AGEMA_signal_2117,
         new_AGEMA_signal_2116, SubCellInst_SboxInst_11_Q2,
         new_AGEMA_signal_2001, new_AGEMA_signal_2000,
         SubCellInst_SboxInst_11_T2, new_AGEMA_signal_2119,
         new_AGEMA_signal_2118, SubCellInst_SboxInst_11_Q7,
         new_AGEMA_signal_2121, new_AGEMA_signal_2120,
         SubCellInst_SboxInst_11_L3, new_AGEMA_signal_2333,
         new_AGEMA_signal_2332, SubCellInst_SboxInst_12_YY_1_,
         new_AGEMA_signal_2253, new_AGEMA_signal_2252,
         SubCellInst_SboxInst_12_YY_0_, new_AGEMA_signal_2005,
         new_AGEMA_signal_2004, SubCellInst_SboxInst_12_T0,
         new_AGEMA_signal_2125, new_AGEMA_signal_2124,
         SubCellInst_SboxInst_12_Q2, new_AGEMA_signal_2007,
         new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2,
         new_AGEMA_signal_2127, new_AGEMA_signal_2126,
         SubCellInst_SboxInst_12_Q7, new_AGEMA_signal_2129,
         new_AGEMA_signal_2128, SubCellInst_SboxInst_12_L3,
         new_AGEMA_signal_2337, new_AGEMA_signal_2336,
         SubCellInst_SboxInst_13_YY_1_, new_AGEMA_signal_2261,
         new_AGEMA_signal_2260, SubCellInst_SboxInst_13_YY_0_,
         new_AGEMA_signal_2011, new_AGEMA_signal_2010,
         SubCellInst_SboxInst_13_T0, new_AGEMA_signal_2133,
         new_AGEMA_signal_2132, SubCellInst_SboxInst_13_Q2,
         new_AGEMA_signal_2013, new_AGEMA_signal_2012,
         SubCellInst_SboxInst_13_T2, new_AGEMA_signal_2135,
         new_AGEMA_signal_2134, SubCellInst_SboxInst_13_Q7,
         new_AGEMA_signal_2137, new_AGEMA_signal_2136,
         SubCellInst_SboxInst_13_L3, new_AGEMA_signal_2341,
         new_AGEMA_signal_2340, SubCellInst_SboxInst_14_YY_1_,
         new_AGEMA_signal_2269, new_AGEMA_signal_2268,
         SubCellInst_SboxInst_14_YY_0_, new_AGEMA_signal_2017,
         new_AGEMA_signal_2016, SubCellInst_SboxInst_14_T0,
         new_AGEMA_signal_2141, new_AGEMA_signal_2140,
         SubCellInst_SboxInst_14_Q2, new_AGEMA_signal_2019,
         new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2,
         new_AGEMA_signal_2143, new_AGEMA_signal_2142,
         SubCellInst_SboxInst_14_Q7, new_AGEMA_signal_2145,
         new_AGEMA_signal_2144, SubCellInst_SboxInst_14_L3,
         new_AGEMA_signal_2345, new_AGEMA_signal_2344,
         SubCellInst_SboxInst_15_YY_1_, new_AGEMA_signal_2277,
         new_AGEMA_signal_2276, SubCellInst_SboxInst_15_YY_0_,
         new_AGEMA_signal_2023, new_AGEMA_signal_2022,
         SubCellInst_SboxInst_15_T0, new_AGEMA_signal_2149,
         new_AGEMA_signal_2148, SubCellInst_SboxInst_15_Q2,
         new_AGEMA_signal_2025, new_AGEMA_signal_2024,
         SubCellInst_SboxInst_15_T2, new_AGEMA_signal_2151,
         new_AGEMA_signal_2150, SubCellInst_SboxInst_15_Q7,
         new_AGEMA_signal_2153, new_AGEMA_signal_2152,
         SubCellInst_SboxInst_15_L3, new_AGEMA_signal_2437,
         new_AGEMA_signal_2436, new_AGEMA_signal_2349, new_AGEMA_signal_2348,
         AddConstXOR_AddConstXOR_XORInst_0_2_n1, new_AGEMA_signal_2523,
         new_AGEMA_signal_2522, new_AGEMA_signal_2439, new_AGEMA_signal_2438,
         AddConstXOR_AddConstXOR_XORInst_0_3_n1, new_AGEMA_signal_2441,
         new_AGEMA_signal_2440, new_AGEMA_signal_2351, new_AGEMA_signal_2350,
         AddConstXOR_AddConstXOR_XORInst_1_2_n1, new_AGEMA_signal_2527,
         new_AGEMA_signal_2526, new_AGEMA_signal_2443, new_AGEMA_signal_2442,
         AddConstXOR_AddConstXOR_XORInst_1_3_n1, new_AGEMA_signal_2445,
         new_AGEMA_signal_2444, new_AGEMA_signal_2353, new_AGEMA_signal_2352,
         AddRoundTweakeyXOR_XORInst_0_2_n1, new_AGEMA_signal_2531,
         new_AGEMA_signal_2530, new_AGEMA_signal_2447, new_AGEMA_signal_2446,
         AddRoundTweakeyXOR_XORInst_0_3_n1, new_AGEMA_signal_2449,
         new_AGEMA_signal_2448, new_AGEMA_signal_2355, new_AGEMA_signal_2354,
         AddRoundTweakeyXOR_XORInst_1_2_n1, new_AGEMA_signal_2535,
         new_AGEMA_signal_2534, new_AGEMA_signal_2451, new_AGEMA_signal_2450,
         AddRoundTweakeyXOR_XORInst_1_3_n1, new_AGEMA_signal_2453,
         new_AGEMA_signal_2452, new_AGEMA_signal_2357, new_AGEMA_signal_2356,
         AddRoundTweakeyXOR_XORInst_2_2_n1, new_AGEMA_signal_2539,
         new_AGEMA_signal_2538, new_AGEMA_signal_2455, new_AGEMA_signal_2454,
         AddRoundTweakeyXOR_XORInst_2_3_n1, new_AGEMA_signal_2617,
         new_AGEMA_signal_2616, new_AGEMA_signal_2541, new_AGEMA_signal_2540,
         AddRoundTweakeyXOR_XORInst_3_2_n1, new_AGEMA_signal_2743,
         new_AGEMA_signal_2742, new_AGEMA_signal_2619, new_AGEMA_signal_2618,
         AddRoundTweakeyXOR_XORInst_3_3_n1, new_AGEMA_signal_2359,
         new_AGEMA_signal_2358, AddRoundTweakeyXOR_XORInst_4_2_n1,
         new_AGEMA_signal_2459, new_AGEMA_signal_2458,
         AddRoundTweakeyXOR_XORInst_4_3_n1, new_AGEMA_signal_2361,
         new_AGEMA_signal_2360, AddRoundTweakeyXOR_XORInst_5_2_n1,
         new_AGEMA_signal_2463, new_AGEMA_signal_2462,
         AddRoundTweakeyXOR_XORInst_5_3_n1, new_AGEMA_signal_2363,
         new_AGEMA_signal_2362, AddRoundTweakeyXOR_XORInst_6_2_n1,
         new_AGEMA_signal_2467, new_AGEMA_signal_2466,
         AddRoundTweakeyXOR_XORInst_6_3_n1, new_AGEMA_signal_2555,
         new_AGEMA_signal_2554, AddRoundTweakeyXOR_XORInst_7_2_n1,
         new_AGEMA_signal_2635, new_AGEMA_signal_2634,
         AddRoundTweakeyXOR_XORInst_7_3_n1, new_AGEMA_signal_2365,
         new_AGEMA_signal_2364, MCInst_MCR0_XORInst_0_2_n1,
         new_AGEMA_signal_2559, new_AGEMA_signal_2558,
         MCInst_MCR0_XORInst_0_2_n2, new_AGEMA_signal_2469,
         new_AGEMA_signal_2468, MCInst_MCR0_XORInst_0_3_n1,
         new_AGEMA_signal_2641, new_AGEMA_signal_2640,
         MCInst_MCR0_XORInst_0_3_n2, new_AGEMA_signal_2367,
         new_AGEMA_signal_2366, MCInst_MCR0_XORInst_1_2_n1,
         new_AGEMA_signal_2563, new_AGEMA_signal_2562,
         MCInst_MCR0_XORInst_1_2_n2, new_AGEMA_signal_2471,
         new_AGEMA_signal_2470, MCInst_MCR0_XORInst_1_3_n1,
         new_AGEMA_signal_2645, new_AGEMA_signal_2644,
         MCInst_MCR0_XORInst_1_3_n2, new_AGEMA_signal_2369,
         new_AGEMA_signal_2368, MCInst_MCR0_XORInst_2_2_n1,
         new_AGEMA_signal_2567, new_AGEMA_signal_2566,
         MCInst_MCR0_XORInst_2_2_n2, new_AGEMA_signal_2473,
         new_AGEMA_signal_2472, MCInst_MCR0_XORInst_2_3_n1,
         new_AGEMA_signal_2651, new_AGEMA_signal_2650,
         MCInst_MCR0_XORInst_2_3_n2, new_AGEMA_signal_2371,
         new_AGEMA_signal_2370, MCInst_MCR0_XORInst_3_2_n1,
         new_AGEMA_signal_2769, new_AGEMA_signal_2768,
         MCInst_MCR0_XORInst_3_2_n2, new_AGEMA_signal_2475,
         new_AGEMA_signal_2474, MCInst_MCR0_XORInst_3_3_n1,
         new_AGEMA_signal_2873, new_AGEMA_signal_2872,
         MCInst_MCR0_XORInst_3_3_n2, new_AGEMA_signal_2571,
         new_AGEMA_signal_2570, MCInst_MCR2_XORInst_0_2_n1,
         new_AGEMA_signal_2657, new_AGEMA_signal_2656,
         MCInst_MCR2_XORInst_0_3_n1, new_AGEMA_signal_2573,
         new_AGEMA_signal_2572, MCInst_MCR2_XORInst_1_2_n1,
         new_AGEMA_signal_2661, new_AGEMA_signal_2660,
         MCInst_MCR2_XORInst_1_3_n1, new_AGEMA_signal_2779,
         new_AGEMA_signal_2778, MCInst_MCR2_XORInst_2_2_n1,
         new_AGEMA_signal_2885, new_AGEMA_signal_2884,
         MCInst_MCR2_XORInst_2_3_n1, new_AGEMA_signal_2575,
         new_AGEMA_signal_2574, MCInst_MCR2_XORInst_3_2_n1,
         new_AGEMA_signal_2665, new_AGEMA_signal_2664,
         MCInst_MCR2_XORInst_3_3_n1, new_AGEMA_signal_2577,
         new_AGEMA_signal_2576, MCInst_MCR3_XORInst_0_2_n1,
         new_AGEMA_signal_2669, new_AGEMA_signal_2668,
         MCInst_MCR3_XORInst_0_3_n1, new_AGEMA_signal_2579,
         new_AGEMA_signal_2578, MCInst_MCR3_XORInst_1_2_n1,
         new_AGEMA_signal_2673, new_AGEMA_signal_2672,
         MCInst_MCR3_XORInst_1_3_n1, new_AGEMA_signal_2581,
         new_AGEMA_signal_2580, MCInst_MCR3_XORInst_2_2_n1,
         new_AGEMA_signal_2677, new_AGEMA_signal_2676,
         MCInst_MCR3_XORInst_2_3_n1, new_AGEMA_signal_2797,
         new_AGEMA_signal_2796, MCInst_MCR3_XORInst_3_2_n1,
         new_AGEMA_signal_2905, new_AGEMA_signal_2904,
         MCInst_MCR3_XORInst_3_3_n1, new_AGEMA_signal_2909,
         new_AGEMA_signal_2908, new_AGEMA_signal_2891, new_AGEMA_signal_2890,
         new_AGEMA_signal_2995, new_AGEMA_signal_2994, new_AGEMA_signal_2983,
         new_AGEMA_signal_2982, new_AGEMA_signal_2913, new_AGEMA_signal_2912,
         new_AGEMA_signal_2895, new_AGEMA_signal_2894, new_AGEMA_signal_2999,
         new_AGEMA_signal_2998, new_AGEMA_signal_2985, new_AGEMA_signal_2984,
         new_AGEMA_signal_2917, new_AGEMA_signal_2916, new_AGEMA_signal_2899,
         new_AGEMA_signal_2898, new_AGEMA_signal_3003, new_AGEMA_signal_3002,
         new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_3059,
         new_AGEMA_signal_3058, new_AGEMA_signal_3053, new_AGEMA_signal_3052,
         new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3073,
         new_AGEMA_signal_3072, new_AGEMA_signal_2925, new_AGEMA_signal_2924,
         new_AGEMA_signal_2875, new_AGEMA_signal_2874, new_AGEMA_signal_3011,
         new_AGEMA_signal_3010, new_AGEMA_signal_2973, new_AGEMA_signal_2972,
         new_AGEMA_signal_2929, new_AGEMA_signal_2928, new_AGEMA_signal_2879,
         new_AGEMA_signal_2878, new_AGEMA_signal_3015, new_AGEMA_signal_3014,
         new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_3063,
         new_AGEMA_signal_3062, new_AGEMA_signal_3049, new_AGEMA_signal_3048,
         new_AGEMA_signal_3081, new_AGEMA_signal_3080, new_AGEMA_signal_3071,
         new_AGEMA_signal_3070, new_AGEMA_signal_2937, new_AGEMA_signal_2936,
         new_AGEMA_signal_2887, new_AGEMA_signal_2886, new_AGEMA_signal_3023,
         new_AGEMA_signal_3022, new_AGEMA_signal_2981, new_AGEMA_signal_2980,
         new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2621,
         new_AGEMA_signal_2620, new_AGEMA_signal_2825, new_AGEMA_signal_2824,
         new_AGEMA_signal_2745, new_AGEMA_signal_2744, new_AGEMA_signal_2709,
         new_AGEMA_signal_2708, new_AGEMA_signal_2625, new_AGEMA_signal_2624,
         new_AGEMA_signal_2829, new_AGEMA_signal_2828, new_AGEMA_signal_2747,
         new_AGEMA_signal_2746, new_AGEMA_signal_2713, new_AGEMA_signal_2712,
         new_AGEMA_signal_2629, new_AGEMA_signal_2628, new_AGEMA_signal_2833,
         new_AGEMA_signal_2832, new_AGEMA_signal_2749, new_AGEMA_signal_2748,
         new_AGEMA_signal_2941, new_AGEMA_signal_2940, new_AGEMA_signal_2855,
         new_AGEMA_signal_2854, new_AGEMA_signal_3027, new_AGEMA_signal_3026,
         new_AGEMA_signal_2961, new_AGEMA_signal_2960, new_AGEMA_signal_2945,
         new_AGEMA_signal_2944, new_AGEMA_signal_2859, new_AGEMA_signal_2858,
         new_AGEMA_signal_3031, new_AGEMA_signal_3030, new_AGEMA_signal_2963,
         new_AGEMA_signal_2962, new_AGEMA_signal_2949, new_AGEMA_signal_2948,
         new_AGEMA_signal_2863, new_AGEMA_signal_2862, new_AGEMA_signal_3035,
         new_AGEMA_signal_3034, new_AGEMA_signal_2965, new_AGEMA_signal_2964,
         new_AGEMA_signal_2953, new_AGEMA_signal_2952, new_AGEMA_signal_2867,
         new_AGEMA_signal_2866, new_AGEMA_signal_3039, new_AGEMA_signal_3038,
         new_AGEMA_signal_2967, new_AGEMA_signal_2966, new_AGEMA_signal_3067,
         new_AGEMA_signal_3066, new_AGEMA_signal_3045, new_AGEMA_signal_3044,
         new_AGEMA_signal_3085, new_AGEMA_signal_3084, new_AGEMA_signal_3069,
         new_AGEMA_signal_3068, new_AGEMA_signal_2159, new_AGEMA_signal_2158,
         SubCellInst_SboxInst_0_T1, new_AGEMA_signal_2287,
         new_AGEMA_signal_2286, SubCellInst_SboxInst_0_L0,
         new_AGEMA_signal_2161, new_AGEMA_signal_2160,
         SubCellInst_SboxInst_0_T3, new_AGEMA_signal_2373,
         new_AGEMA_signal_2372, SubCellInst_SboxInst_0_YY_3,
         new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2489,
         new_AGEMA_signal_2488, new_AGEMA_signal_2167, new_AGEMA_signal_2166,
         SubCellInst_SboxInst_1_T1, new_AGEMA_signal_2291,
         new_AGEMA_signal_2290, SubCellInst_SboxInst_1_L0,
         new_AGEMA_signal_2169, new_AGEMA_signal_2168,
         SubCellInst_SboxInst_1_T3, new_AGEMA_signal_2377,
         new_AGEMA_signal_2376, SubCellInst_SboxInst_1_YY_3,
         new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2491,
         new_AGEMA_signal_2490, new_AGEMA_signal_2175, new_AGEMA_signal_2174,
         SubCellInst_SboxInst_2_T1, new_AGEMA_signal_2295,
         new_AGEMA_signal_2294, SubCellInst_SboxInst_2_L0,
         new_AGEMA_signal_2177, new_AGEMA_signal_2176,
         SubCellInst_SboxInst_2_T3, new_AGEMA_signal_2381,
         new_AGEMA_signal_2380, SubCellInst_SboxInst_2_YY_3,
         new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2493,
         new_AGEMA_signal_2492, new_AGEMA_signal_2183, new_AGEMA_signal_2182,
         SubCellInst_SboxInst_3_T1, new_AGEMA_signal_2299,
         new_AGEMA_signal_2298, SubCellInst_SboxInst_3_L0,
         new_AGEMA_signal_2185, new_AGEMA_signal_2184,
         SubCellInst_SboxInst_3_T3, new_AGEMA_signal_2385,
         new_AGEMA_signal_2384, SubCellInst_SboxInst_3_YY_3,
         new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2495,
         new_AGEMA_signal_2494, new_AGEMA_signal_2191, new_AGEMA_signal_2190,
         SubCellInst_SboxInst_4_T1, new_AGEMA_signal_2303,
         new_AGEMA_signal_2302, SubCellInst_SboxInst_4_L0,
         new_AGEMA_signal_2193, new_AGEMA_signal_2192,
         SubCellInst_SboxInst_4_T3, new_AGEMA_signal_2389,
         new_AGEMA_signal_2388, SubCellInst_SboxInst_4_YY_3,
         new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2497,
         new_AGEMA_signal_2496, new_AGEMA_signal_2199, new_AGEMA_signal_2198,
         SubCellInst_SboxInst_5_T1, new_AGEMA_signal_2307,
         new_AGEMA_signal_2306, SubCellInst_SboxInst_5_L0,
         new_AGEMA_signal_2201, new_AGEMA_signal_2200,
         SubCellInst_SboxInst_5_T3, new_AGEMA_signal_2393,
         new_AGEMA_signal_2392, SubCellInst_SboxInst_5_YY_3,
         new_AGEMA_signal_2395, new_AGEMA_signal_2394, new_AGEMA_signal_2499,
         new_AGEMA_signal_2498, new_AGEMA_signal_2207, new_AGEMA_signal_2206,
         SubCellInst_SboxInst_6_T1, new_AGEMA_signal_2311,
         new_AGEMA_signal_2310, SubCellInst_SboxInst_6_L0,
         new_AGEMA_signal_2209, new_AGEMA_signal_2208,
         SubCellInst_SboxInst_6_T3, new_AGEMA_signal_2397,
         new_AGEMA_signal_2396, SubCellInst_SboxInst_6_YY_3,
         new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2501,
         new_AGEMA_signal_2500, new_AGEMA_signal_2215, new_AGEMA_signal_2214,
         SubCellInst_SboxInst_7_T1, new_AGEMA_signal_2315,
         new_AGEMA_signal_2314, SubCellInst_SboxInst_7_L0,
         new_AGEMA_signal_2217, new_AGEMA_signal_2216,
         SubCellInst_SboxInst_7_T3, new_AGEMA_signal_2401,
         new_AGEMA_signal_2400, SubCellInst_SboxInst_7_YY_3,
         new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2223,
         new_AGEMA_signal_2222, SubCellInst_SboxInst_8_T1,
         new_AGEMA_signal_2319, new_AGEMA_signal_2318,
         SubCellInst_SboxInst_8_L0, new_AGEMA_signal_2225,
         new_AGEMA_signal_2224, SubCellInst_SboxInst_8_T3,
         new_AGEMA_signal_2405, new_AGEMA_signal_2404,
         SubCellInst_SboxInst_8_YY_3, new_AGEMA_signal_2407,
         new_AGEMA_signal_2406, new_AGEMA_signal_2505, new_AGEMA_signal_2504,
         new_AGEMA_signal_2231, new_AGEMA_signal_2230,
         SubCellInst_SboxInst_9_T1, new_AGEMA_signal_2323,
         new_AGEMA_signal_2322, SubCellInst_SboxInst_9_L0,
         new_AGEMA_signal_2233, new_AGEMA_signal_2232,
         SubCellInst_SboxInst_9_T3, new_AGEMA_signal_2409,
         new_AGEMA_signal_2408, SubCellInst_SboxInst_9_YY_3,
         new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2507,
         new_AGEMA_signal_2506, new_AGEMA_signal_2239, new_AGEMA_signal_2238,
         SubCellInst_SboxInst_10_T1, new_AGEMA_signal_2327,
         new_AGEMA_signal_2326, SubCellInst_SboxInst_10_L0,
         new_AGEMA_signal_2241, new_AGEMA_signal_2240,
         SubCellInst_SboxInst_10_T3, new_AGEMA_signal_2413,
         new_AGEMA_signal_2412, SubCellInst_SboxInst_10_YY_3,
         new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2509,
         new_AGEMA_signal_2508, new_AGEMA_signal_2247, new_AGEMA_signal_2246,
         SubCellInst_SboxInst_11_T1, new_AGEMA_signal_2331,
         new_AGEMA_signal_2330, SubCellInst_SboxInst_11_L0,
         new_AGEMA_signal_2249, new_AGEMA_signal_2248,
         SubCellInst_SboxInst_11_T3, new_AGEMA_signal_2417,
         new_AGEMA_signal_2416, SubCellInst_SboxInst_11_YY_3,
         new_AGEMA_signal_2419, new_AGEMA_signal_2418, new_AGEMA_signal_2511,
         new_AGEMA_signal_2510, new_AGEMA_signal_2255, new_AGEMA_signal_2254,
         SubCellInst_SboxInst_12_T1, new_AGEMA_signal_2335,
         new_AGEMA_signal_2334, SubCellInst_SboxInst_12_L0,
         new_AGEMA_signal_2257, new_AGEMA_signal_2256,
         SubCellInst_SboxInst_12_T3, new_AGEMA_signal_2421,
         new_AGEMA_signal_2420, SubCellInst_SboxInst_12_YY_3,
         new_AGEMA_signal_2423, new_AGEMA_signal_2422, new_AGEMA_signal_2513,
         new_AGEMA_signal_2512, new_AGEMA_signal_2263, new_AGEMA_signal_2262,
         SubCellInst_SboxInst_13_T1, new_AGEMA_signal_2339,
         new_AGEMA_signal_2338, SubCellInst_SboxInst_13_L0,
         new_AGEMA_signal_2265, new_AGEMA_signal_2264,
         SubCellInst_SboxInst_13_T3, new_AGEMA_signal_2425,
         new_AGEMA_signal_2424, SubCellInst_SboxInst_13_YY_3,
         new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2515,
         new_AGEMA_signal_2514, new_AGEMA_signal_2271, new_AGEMA_signal_2270,
         SubCellInst_SboxInst_14_T1, new_AGEMA_signal_2343,
         new_AGEMA_signal_2342, SubCellInst_SboxInst_14_L0,
         new_AGEMA_signal_2273, new_AGEMA_signal_2272,
         SubCellInst_SboxInst_14_T3, new_AGEMA_signal_2429,
         new_AGEMA_signal_2428, SubCellInst_SboxInst_14_YY_3,
         new_AGEMA_signal_2431, new_AGEMA_signal_2430, new_AGEMA_signal_2517,
         new_AGEMA_signal_2516, new_AGEMA_signal_2279, new_AGEMA_signal_2278,
         SubCellInst_SboxInst_15_T1, new_AGEMA_signal_2347,
         new_AGEMA_signal_2346, SubCellInst_SboxInst_15_L0,
         new_AGEMA_signal_2281, new_AGEMA_signal_2280,
         SubCellInst_SboxInst_15_T3, new_AGEMA_signal_2433,
         new_AGEMA_signal_2432, SubCellInst_SboxInst_15_YY_3,
         new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2519,
         new_AGEMA_signal_2518, new_AGEMA_signal_2595, new_AGEMA_signal_2594,
         new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2521,
         new_AGEMA_signal_2520, AddConstXOR_AddConstXOR_XORInst_0_0_n1,
         new_AGEMA_signal_2731, new_AGEMA_signal_2730, new_AGEMA_signal_2599,
         new_AGEMA_signal_2598, AddConstXOR_AddConstXOR_XORInst_0_1_n1,
         new_AGEMA_signal_2601, new_AGEMA_signal_2600, new_AGEMA_signal_2525,
         new_AGEMA_signal_2524, AddConstXOR_AddConstXOR_XORInst_1_0_n1,
         new_AGEMA_signal_2733, new_AGEMA_signal_2732, new_AGEMA_signal_2603,
         new_AGEMA_signal_2602, AddConstXOR_AddConstXOR_XORInst_1_1_n1,
         new_AGEMA_signal_2605, new_AGEMA_signal_2604, new_AGEMA_signal_2529,
         new_AGEMA_signal_2528, AddRoundTweakeyXOR_XORInst_0_0_n1,
         new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2607,
         new_AGEMA_signal_2606, AddRoundTweakeyXOR_XORInst_0_1_n1,
         new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2533,
         new_AGEMA_signal_2532, AddRoundTweakeyXOR_XORInst_1_0_n1,
         new_AGEMA_signal_2737, new_AGEMA_signal_2736, new_AGEMA_signal_2611,
         new_AGEMA_signal_2610, AddRoundTweakeyXOR_XORInst_1_1_n1,
         new_AGEMA_signal_2613, new_AGEMA_signal_2612, new_AGEMA_signal_2537,
         new_AGEMA_signal_2536, AddRoundTweakeyXOR_XORInst_2_0_n1,
         new_AGEMA_signal_2739, new_AGEMA_signal_2738, new_AGEMA_signal_2615,
         new_AGEMA_signal_2614, AddRoundTweakeyXOR_XORInst_2_1_n1,
         new_AGEMA_signal_2851, new_AGEMA_signal_2850, new_AGEMA_signal_2741,
         new_AGEMA_signal_2740, AddRoundTweakeyXOR_XORInst_3_0_n1,
         new_AGEMA_signal_2959, new_AGEMA_signal_2958, new_AGEMA_signal_2853,
         new_AGEMA_signal_2852, AddRoundTweakeyXOR_XORInst_3_1_n1,
         new_AGEMA_signal_2543, new_AGEMA_signal_2542,
         AddRoundTweakeyXOR_XORInst_4_0_n1, new_AGEMA_signal_2623,
         new_AGEMA_signal_2622, AddRoundTweakeyXOR_XORInst_4_1_n1,
         new_AGEMA_signal_2547, new_AGEMA_signal_2546,
         AddRoundTweakeyXOR_XORInst_5_0_n1, new_AGEMA_signal_2627,
         new_AGEMA_signal_2626, AddRoundTweakeyXOR_XORInst_5_1_n1,
         new_AGEMA_signal_2551, new_AGEMA_signal_2550,
         AddRoundTweakeyXOR_XORInst_6_0_n1, new_AGEMA_signal_2631,
         new_AGEMA_signal_2630, AddRoundTweakeyXOR_XORInst_6_1_n1,
         new_AGEMA_signal_2751, new_AGEMA_signal_2750,
         AddRoundTweakeyXOR_XORInst_7_0_n1, new_AGEMA_signal_2857,
         new_AGEMA_signal_2856, AddRoundTweakeyXOR_XORInst_7_1_n1,
         new_AGEMA_signal_2557, new_AGEMA_signal_2556,
         MCInst_MCR0_XORInst_0_0_n1, new_AGEMA_signal_2755,
         new_AGEMA_signal_2754, MCInst_MCR0_XORInst_0_0_n2,
         new_AGEMA_signal_2637, new_AGEMA_signal_2636,
         MCInst_MCR0_XORInst_0_1_n1, new_AGEMA_signal_2861,
         new_AGEMA_signal_2860, MCInst_MCR0_XORInst_0_1_n2,
         new_AGEMA_signal_2561, new_AGEMA_signal_2560,
         MCInst_MCR0_XORInst_1_0_n1, new_AGEMA_signal_2759,
         new_AGEMA_signal_2758, MCInst_MCR0_XORInst_1_0_n2,
         new_AGEMA_signal_2761, new_AGEMA_signal_2760,
         MCInst_MCR0_XORInst_1_1_n1, new_AGEMA_signal_2865,
         new_AGEMA_signal_2864, MCInst_MCR0_XORInst_1_1_n2,
         new_AGEMA_signal_2565, new_AGEMA_signal_2564,
         MCInst_MCR0_XORInst_2_0_n1, new_AGEMA_signal_2765,
         new_AGEMA_signal_2764, MCInst_MCR0_XORInst_2_0_n2,
         new_AGEMA_signal_2647, new_AGEMA_signal_2646,
         MCInst_MCR0_XORInst_2_1_n1, new_AGEMA_signal_2869,
         new_AGEMA_signal_2868, MCInst_MCR0_XORInst_2_1_n2,
         new_AGEMA_signal_2569, new_AGEMA_signal_2568,
         MCInst_MCR0_XORInst_3_0_n1, new_AGEMA_signal_2969,
         new_AGEMA_signal_2968, MCInst_MCR0_XORInst_3_0_n2,
         new_AGEMA_signal_2653, new_AGEMA_signal_2652,
         MCInst_MCR0_XORInst_3_1_n1, new_AGEMA_signal_3047,
         new_AGEMA_signal_3046, MCInst_MCR0_XORInst_3_1_n2,
         new_AGEMA_signal_2771, new_AGEMA_signal_2770,
         MCInst_MCR2_XORInst_0_0_n1, new_AGEMA_signal_2877,
         new_AGEMA_signal_2876, MCInst_MCR2_XORInst_0_1_n1,
         new_AGEMA_signal_2775, new_AGEMA_signal_2774,
         MCInst_MCR2_XORInst_1_0_n1, new_AGEMA_signal_2881,
         new_AGEMA_signal_2880, MCInst_MCR2_XORInst_1_1_n1,
         new_AGEMA_signal_2977, new_AGEMA_signal_2976,
         MCInst_MCR2_XORInst_2_0_n1, new_AGEMA_signal_3051,
         new_AGEMA_signal_3050, MCInst_MCR2_XORInst_2_1_n1,
         new_AGEMA_signal_2781, new_AGEMA_signal_2780,
         MCInst_MCR2_XORInst_3_0_n1, new_AGEMA_signal_2889,
         new_AGEMA_signal_2888, MCInst_MCR2_XORInst_3_1_n1,
         new_AGEMA_signal_2785, new_AGEMA_signal_2784,
         MCInst_MCR3_XORInst_0_0_n1, new_AGEMA_signal_2893,
         new_AGEMA_signal_2892, MCInst_MCR3_XORInst_0_1_n1,
         new_AGEMA_signal_2789, new_AGEMA_signal_2788,
         MCInst_MCR3_XORInst_1_0_n1, new_AGEMA_signal_2897,
         new_AGEMA_signal_2896, MCInst_MCR3_XORInst_1_1_n1,
         new_AGEMA_signal_2793, new_AGEMA_signal_2792,
         MCInst_MCR3_XORInst_2_0_n1, new_AGEMA_signal_2901,
         new_AGEMA_signal_2900, MCInst_MCR3_XORInst_2_1_n1,
         new_AGEMA_signal_2989, new_AGEMA_signal_2988,
         MCInst_MCR3_XORInst_3_0_n1, new_AGEMA_signal_3055,
         new_AGEMA_signal_3054, MCInst_MCR3_XORInst_3_1_n1, n13, n14, n15, n16,
         n17, n18, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         ClockGatingInst_n11, ClockGatingInst_n10, ClockGatingInst_n9,
         ClockGatingInst_n8, ClockGatingInst_n7, ClockGatingInst_n6,
         ClockGatingInst_n4, ClockGatingInst_n3, ClockGatingInst_n2,
         ClockGatingInst_n1, ClockGatingInst_LatchedEnable, ClockGatingInst_N7,
         ClockGatingInst_ShiftRegister_5_, SubCellInst_SboxInst_0_AND1_U1_n36,
         SubCellInst_SboxInst_0_AND1_U1_n35,
         SubCellInst_SboxInst_0_AND1_U1_n34,
         SubCellInst_SboxInst_0_AND1_U1_n33,
         SubCellInst_SboxInst_0_AND1_U1_n32,
         SubCellInst_SboxInst_0_AND1_U1_n31,
         SubCellInst_SboxInst_0_AND1_U1_n30,
         SubCellInst_SboxInst_0_AND1_U1_n29,
         SubCellInst_SboxInst_0_AND1_U1_n28,
         SubCellInst_SboxInst_0_AND1_U1_n27,
         SubCellInst_SboxInst_0_AND1_U1_n26,
         SubCellInst_SboxInst_0_AND1_U1_n25,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_0_AND3_U1_n36,
         SubCellInst_SboxInst_0_AND3_U1_n35,
         SubCellInst_SboxInst_0_AND3_U1_n34,
         SubCellInst_SboxInst_0_AND3_U1_n33,
         SubCellInst_SboxInst_0_AND3_U1_n32,
         SubCellInst_SboxInst_0_AND3_U1_n31,
         SubCellInst_SboxInst_0_AND3_U1_n30,
         SubCellInst_SboxInst_0_AND3_U1_n29,
         SubCellInst_SboxInst_0_AND3_U1_n28,
         SubCellInst_SboxInst_0_AND3_U1_n27,
         SubCellInst_SboxInst_0_AND3_U1_n26,
         SubCellInst_SboxInst_0_AND3_U1_n25,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND1_U1_n36,
         SubCellInst_SboxInst_1_AND1_U1_n35,
         SubCellInst_SboxInst_1_AND1_U1_n34,
         SubCellInst_SboxInst_1_AND1_U1_n33,
         SubCellInst_SboxInst_1_AND1_U1_n32,
         SubCellInst_SboxInst_1_AND1_U1_n31,
         SubCellInst_SboxInst_1_AND1_U1_n30,
         SubCellInst_SboxInst_1_AND1_U1_n29,
         SubCellInst_SboxInst_1_AND1_U1_n28,
         SubCellInst_SboxInst_1_AND1_U1_n27,
         SubCellInst_SboxInst_1_AND1_U1_n26,
         SubCellInst_SboxInst_1_AND1_U1_n25,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND3_U1_n36,
         SubCellInst_SboxInst_1_AND3_U1_n35,
         SubCellInst_SboxInst_1_AND3_U1_n34,
         SubCellInst_SboxInst_1_AND3_U1_n33,
         SubCellInst_SboxInst_1_AND3_U1_n32,
         SubCellInst_SboxInst_1_AND3_U1_n31,
         SubCellInst_SboxInst_1_AND3_U1_n30,
         SubCellInst_SboxInst_1_AND3_U1_n29,
         SubCellInst_SboxInst_1_AND3_U1_n28,
         SubCellInst_SboxInst_1_AND3_U1_n27,
         SubCellInst_SboxInst_1_AND3_U1_n26,
         SubCellInst_SboxInst_1_AND3_U1_n25,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND1_U1_n36,
         SubCellInst_SboxInst_2_AND1_U1_n35,
         SubCellInst_SboxInst_2_AND1_U1_n34,
         SubCellInst_SboxInst_2_AND1_U1_n33,
         SubCellInst_SboxInst_2_AND1_U1_n32,
         SubCellInst_SboxInst_2_AND1_U1_n31,
         SubCellInst_SboxInst_2_AND1_U1_n30,
         SubCellInst_SboxInst_2_AND1_U1_n29,
         SubCellInst_SboxInst_2_AND1_U1_n28,
         SubCellInst_SboxInst_2_AND1_U1_n27,
         SubCellInst_SboxInst_2_AND1_U1_n26,
         SubCellInst_SboxInst_2_AND1_U1_n25,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND3_U1_n36,
         SubCellInst_SboxInst_2_AND3_U1_n35,
         SubCellInst_SboxInst_2_AND3_U1_n34,
         SubCellInst_SboxInst_2_AND3_U1_n33,
         SubCellInst_SboxInst_2_AND3_U1_n32,
         SubCellInst_SboxInst_2_AND3_U1_n31,
         SubCellInst_SboxInst_2_AND3_U1_n30,
         SubCellInst_SboxInst_2_AND3_U1_n29,
         SubCellInst_SboxInst_2_AND3_U1_n28,
         SubCellInst_SboxInst_2_AND3_U1_n27,
         SubCellInst_SboxInst_2_AND3_U1_n26,
         SubCellInst_SboxInst_2_AND3_U1_n25,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND1_U1_n36,
         SubCellInst_SboxInst_3_AND1_U1_n35,
         SubCellInst_SboxInst_3_AND1_U1_n34,
         SubCellInst_SboxInst_3_AND1_U1_n33,
         SubCellInst_SboxInst_3_AND1_U1_n32,
         SubCellInst_SboxInst_3_AND1_U1_n31,
         SubCellInst_SboxInst_3_AND1_U1_n30,
         SubCellInst_SboxInst_3_AND1_U1_n29,
         SubCellInst_SboxInst_3_AND1_U1_n28,
         SubCellInst_SboxInst_3_AND1_U1_n27,
         SubCellInst_SboxInst_3_AND1_U1_n26,
         SubCellInst_SboxInst_3_AND1_U1_n25,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND3_U1_n36,
         SubCellInst_SboxInst_3_AND3_U1_n35,
         SubCellInst_SboxInst_3_AND3_U1_n34,
         SubCellInst_SboxInst_3_AND3_U1_n33,
         SubCellInst_SboxInst_3_AND3_U1_n32,
         SubCellInst_SboxInst_3_AND3_U1_n31,
         SubCellInst_SboxInst_3_AND3_U1_n30,
         SubCellInst_SboxInst_3_AND3_U1_n29,
         SubCellInst_SboxInst_3_AND3_U1_n28,
         SubCellInst_SboxInst_3_AND3_U1_n27,
         SubCellInst_SboxInst_3_AND3_U1_n26,
         SubCellInst_SboxInst_3_AND3_U1_n25,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND1_U1_n36,
         SubCellInst_SboxInst_4_AND1_U1_n35,
         SubCellInst_SboxInst_4_AND1_U1_n34,
         SubCellInst_SboxInst_4_AND1_U1_n33,
         SubCellInst_SboxInst_4_AND1_U1_n32,
         SubCellInst_SboxInst_4_AND1_U1_n31,
         SubCellInst_SboxInst_4_AND1_U1_n30,
         SubCellInst_SboxInst_4_AND1_U1_n29,
         SubCellInst_SboxInst_4_AND1_U1_n28,
         SubCellInst_SboxInst_4_AND1_U1_n27,
         SubCellInst_SboxInst_4_AND1_U1_n26,
         SubCellInst_SboxInst_4_AND1_U1_n25,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND3_U1_n36,
         SubCellInst_SboxInst_4_AND3_U1_n35,
         SubCellInst_SboxInst_4_AND3_U1_n34,
         SubCellInst_SboxInst_4_AND3_U1_n33,
         SubCellInst_SboxInst_4_AND3_U1_n32,
         SubCellInst_SboxInst_4_AND3_U1_n31,
         SubCellInst_SboxInst_4_AND3_U1_n30,
         SubCellInst_SboxInst_4_AND3_U1_n29,
         SubCellInst_SboxInst_4_AND3_U1_n28,
         SubCellInst_SboxInst_4_AND3_U1_n27,
         SubCellInst_SboxInst_4_AND3_U1_n26,
         SubCellInst_SboxInst_4_AND3_U1_n25,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND1_U1_n36,
         SubCellInst_SboxInst_5_AND1_U1_n35,
         SubCellInst_SboxInst_5_AND1_U1_n34,
         SubCellInst_SboxInst_5_AND1_U1_n33,
         SubCellInst_SboxInst_5_AND1_U1_n32,
         SubCellInst_SboxInst_5_AND1_U1_n31,
         SubCellInst_SboxInst_5_AND1_U1_n30,
         SubCellInst_SboxInst_5_AND1_U1_n29,
         SubCellInst_SboxInst_5_AND1_U1_n28,
         SubCellInst_SboxInst_5_AND1_U1_n27,
         SubCellInst_SboxInst_5_AND1_U1_n26,
         SubCellInst_SboxInst_5_AND1_U1_n25,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND3_U1_n36,
         SubCellInst_SboxInst_5_AND3_U1_n35,
         SubCellInst_SboxInst_5_AND3_U1_n34,
         SubCellInst_SboxInst_5_AND3_U1_n33,
         SubCellInst_SboxInst_5_AND3_U1_n32,
         SubCellInst_SboxInst_5_AND3_U1_n31,
         SubCellInst_SboxInst_5_AND3_U1_n30,
         SubCellInst_SboxInst_5_AND3_U1_n29,
         SubCellInst_SboxInst_5_AND3_U1_n28,
         SubCellInst_SboxInst_5_AND3_U1_n27,
         SubCellInst_SboxInst_5_AND3_U1_n26,
         SubCellInst_SboxInst_5_AND3_U1_n25,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND1_U1_n36,
         SubCellInst_SboxInst_6_AND1_U1_n35,
         SubCellInst_SboxInst_6_AND1_U1_n34,
         SubCellInst_SboxInst_6_AND1_U1_n33,
         SubCellInst_SboxInst_6_AND1_U1_n32,
         SubCellInst_SboxInst_6_AND1_U1_n31,
         SubCellInst_SboxInst_6_AND1_U1_n30,
         SubCellInst_SboxInst_6_AND1_U1_n29,
         SubCellInst_SboxInst_6_AND1_U1_n28,
         SubCellInst_SboxInst_6_AND1_U1_n27,
         SubCellInst_SboxInst_6_AND1_U1_n26,
         SubCellInst_SboxInst_6_AND1_U1_n25,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND3_U1_n36,
         SubCellInst_SboxInst_6_AND3_U1_n35,
         SubCellInst_SboxInst_6_AND3_U1_n34,
         SubCellInst_SboxInst_6_AND3_U1_n33,
         SubCellInst_SboxInst_6_AND3_U1_n32,
         SubCellInst_SboxInst_6_AND3_U1_n31,
         SubCellInst_SboxInst_6_AND3_U1_n30,
         SubCellInst_SboxInst_6_AND3_U1_n29,
         SubCellInst_SboxInst_6_AND3_U1_n28,
         SubCellInst_SboxInst_6_AND3_U1_n27,
         SubCellInst_SboxInst_6_AND3_U1_n26,
         SubCellInst_SboxInst_6_AND3_U1_n25,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND1_U1_n36,
         SubCellInst_SboxInst_7_AND1_U1_n35,
         SubCellInst_SboxInst_7_AND1_U1_n34,
         SubCellInst_SboxInst_7_AND1_U1_n33,
         SubCellInst_SboxInst_7_AND1_U1_n32,
         SubCellInst_SboxInst_7_AND1_U1_n31,
         SubCellInst_SboxInst_7_AND1_U1_n30,
         SubCellInst_SboxInst_7_AND1_U1_n29,
         SubCellInst_SboxInst_7_AND1_U1_n28,
         SubCellInst_SboxInst_7_AND1_U1_n27,
         SubCellInst_SboxInst_7_AND1_U1_n26,
         SubCellInst_SboxInst_7_AND1_U1_n25,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND3_U1_n36,
         SubCellInst_SboxInst_7_AND3_U1_n35,
         SubCellInst_SboxInst_7_AND3_U1_n34,
         SubCellInst_SboxInst_7_AND3_U1_n33,
         SubCellInst_SboxInst_7_AND3_U1_n32,
         SubCellInst_SboxInst_7_AND3_U1_n31,
         SubCellInst_SboxInst_7_AND3_U1_n30,
         SubCellInst_SboxInst_7_AND3_U1_n29,
         SubCellInst_SboxInst_7_AND3_U1_n28,
         SubCellInst_SboxInst_7_AND3_U1_n27,
         SubCellInst_SboxInst_7_AND3_U1_n26,
         SubCellInst_SboxInst_7_AND3_U1_n25,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND1_U1_n36,
         SubCellInst_SboxInst_8_AND1_U1_n35,
         SubCellInst_SboxInst_8_AND1_U1_n34,
         SubCellInst_SboxInst_8_AND1_U1_n33,
         SubCellInst_SboxInst_8_AND1_U1_n32,
         SubCellInst_SboxInst_8_AND1_U1_n31,
         SubCellInst_SboxInst_8_AND1_U1_n30,
         SubCellInst_SboxInst_8_AND1_U1_n29,
         SubCellInst_SboxInst_8_AND1_U1_n28,
         SubCellInst_SboxInst_8_AND1_U1_n27,
         SubCellInst_SboxInst_8_AND1_U1_n26,
         SubCellInst_SboxInst_8_AND1_U1_n25,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND3_U1_n36,
         SubCellInst_SboxInst_8_AND3_U1_n35,
         SubCellInst_SboxInst_8_AND3_U1_n34,
         SubCellInst_SboxInst_8_AND3_U1_n33,
         SubCellInst_SboxInst_8_AND3_U1_n32,
         SubCellInst_SboxInst_8_AND3_U1_n31,
         SubCellInst_SboxInst_8_AND3_U1_n30,
         SubCellInst_SboxInst_8_AND3_U1_n29,
         SubCellInst_SboxInst_8_AND3_U1_n28,
         SubCellInst_SboxInst_8_AND3_U1_n27,
         SubCellInst_SboxInst_8_AND3_U1_n26,
         SubCellInst_SboxInst_8_AND3_U1_n25,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND1_U1_n36,
         SubCellInst_SboxInst_9_AND1_U1_n35,
         SubCellInst_SboxInst_9_AND1_U1_n34,
         SubCellInst_SboxInst_9_AND1_U1_n33,
         SubCellInst_SboxInst_9_AND1_U1_n32,
         SubCellInst_SboxInst_9_AND1_U1_n31,
         SubCellInst_SboxInst_9_AND1_U1_n30,
         SubCellInst_SboxInst_9_AND1_U1_n29,
         SubCellInst_SboxInst_9_AND1_U1_n28,
         SubCellInst_SboxInst_9_AND1_U1_n27,
         SubCellInst_SboxInst_9_AND1_U1_n26,
         SubCellInst_SboxInst_9_AND1_U1_n25,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND3_U1_n36,
         SubCellInst_SboxInst_9_AND3_U1_n35,
         SubCellInst_SboxInst_9_AND3_U1_n34,
         SubCellInst_SboxInst_9_AND3_U1_n33,
         SubCellInst_SboxInst_9_AND3_U1_n32,
         SubCellInst_SboxInst_9_AND3_U1_n31,
         SubCellInst_SboxInst_9_AND3_U1_n30,
         SubCellInst_SboxInst_9_AND3_U1_n29,
         SubCellInst_SboxInst_9_AND3_U1_n28,
         SubCellInst_SboxInst_9_AND3_U1_n27,
         SubCellInst_SboxInst_9_AND3_U1_n26,
         SubCellInst_SboxInst_9_AND3_U1_n25,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND1_U1_n36,
         SubCellInst_SboxInst_10_AND1_U1_n35,
         SubCellInst_SboxInst_10_AND1_U1_n34,
         SubCellInst_SboxInst_10_AND1_U1_n33,
         SubCellInst_SboxInst_10_AND1_U1_n32,
         SubCellInst_SboxInst_10_AND1_U1_n31,
         SubCellInst_SboxInst_10_AND1_U1_n30,
         SubCellInst_SboxInst_10_AND1_U1_n29,
         SubCellInst_SboxInst_10_AND1_U1_n28,
         SubCellInst_SboxInst_10_AND1_U1_n27,
         SubCellInst_SboxInst_10_AND1_U1_n26,
         SubCellInst_SboxInst_10_AND1_U1_n25,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND3_U1_n36,
         SubCellInst_SboxInst_10_AND3_U1_n35,
         SubCellInst_SboxInst_10_AND3_U1_n34,
         SubCellInst_SboxInst_10_AND3_U1_n33,
         SubCellInst_SboxInst_10_AND3_U1_n32,
         SubCellInst_SboxInst_10_AND3_U1_n31,
         SubCellInst_SboxInst_10_AND3_U1_n30,
         SubCellInst_SboxInst_10_AND3_U1_n29,
         SubCellInst_SboxInst_10_AND3_U1_n28,
         SubCellInst_SboxInst_10_AND3_U1_n27,
         SubCellInst_SboxInst_10_AND3_U1_n26,
         SubCellInst_SboxInst_10_AND3_U1_n25,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND1_U1_n36,
         SubCellInst_SboxInst_11_AND1_U1_n35,
         SubCellInst_SboxInst_11_AND1_U1_n34,
         SubCellInst_SboxInst_11_AND1_U1_n33,
         SubCellInst_SboxInst_11_AND1_U1_n32,
         SubCellInst_SboxInst_11_AND1_U1_n31,
         SubCellInst_SboxInst_11_AND1_U1_n30,
         SubCellInst_SboxInst_11_AND1_U1_n29,
         SubCellInst_SboxInst_11_AND1_U1_n28,
         SubCellInst_SboxInst_11_AND1_U1_n27,
         SubCellInst_SboxInst_11_AND1_U1_n26,
         SubCellInst_SboxInst_11_AND1_U1_n25,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND3_U1_n36,
         SubCellInst_SboxInst_11_AND3_U1_n35,
         SubCellInst_SboxInst_11_AND3_U1_n34,
         SubCellInst_SboxInst_11_AND3_U1_n33,
         SubCellInst_SboxInst_11_AND3_U1_n32,
         SubCellInst_SboxInst_11_AND3_U1_n31,
         SubCellInst_SboxInst_11_AND3_U1_n30,
         SubCellInst_SboxInst_11_AND3_U1_n29,
         SubCellInst_SboxInst_11_AND3_U1_n28,
         SubCellInst_SboxInst_11_AND3_U1_n27,
         SubCellInst_SboxInst_11_AND3_U1_n26,
         SubCellInst_SboxInst_11_AND3_U1_n25,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND1_U1_n36,
         SubCellInst_SboxInst_12_AND1_U1_n35,
         SubCellInst_SboxInst_12_AND1_U1_n34,
         SubCellInst_SboxInst_12_AND1_U1_n33,
         SubCellInst_SboxInst_12_AND1_U1_n32,
         SubCellInst_SboxInst_12_AND1_U1_n31,
         SubCellInst_SboxInst_12_AND1_U1_n30,
         SubCellInst_SboxInst_12_AND1_U1_n29,
         SubCellInst_SboxInst_12_AND1_U1_n28,
         SubCellInst_SboxInst_12_AND1_U1_n27,
         SubCellInst_SboxInst_12_AND1_U1_n26,
         SubCellInst_SboxInst_12_AND1_U1_n25,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND3_U1_n36,
         SubCellInst_SboxInst_12_AND3_U1_n35,
         SubCellInst_SboxInst_12_AND3_U1_n34,
         SubCellInst_SboxInst_12_AND3_U1_n33,
         SubCellInst_SboxInst_12_AND3_U1_n32,
         SubCellInst_SboxInst_12_AND3_U1_n31,
         SubCellInst_SboxInst_12_AND3_U1_n30,
         SubCellInst_SboxInst_12_AND3_U1_n29,
         SubCellInst_SboxInst_12_AND3_U1_n28,
         SubCellInst_SboxInst_12_AND3_U1_n27,
         SubCellInst_SboxInst_12_AND3_U1_n26,
         SubCellInst_SboxInst_12_AND3_U1_n25,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND1_U1_n36,
         SubCellInst_SboxInst_13_AND1_U1_n35,
         SubCellInst_SboxInst_13_AND1_U1_n34,
         SubCellInst_SboxInst_13_AND1_U1_n33,
         SubCellInst_SboxInst_13_AND1_U1_n32,
         SubCellInst_SboxInst_13_AND1_U1_n31,
         SubCellInst_SboxInst_13_AND1_U1_n30,
         SubCellInst_SboxInst_13_AND1_U1_n29,
         SubCellInst_SboxInst_13_AND1_U1_n28,
         SubCellInst_SboxInst_13_AND1_U1_n27,
         SubCellInst_SboxInst_13_AND1_U1_n26,
         SubCellInst_SboxInst_13_AND1_U1_n25,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND3_U1_n36,
         SubCellInst_SboxInst_13_AND3_U1_n35,
         SubCellInst_SboxInst_13_AND3_U1_n34,
         SubCellInst_SboxInst_13_AND3_U1_n33,
         SubCellInst_SboxInst_13_AND3_U1_n32,
         SubCellInst_SboxInst_13_AND3_U1_n31,
         SubCellInst_SboxInst_13_AND3_U1_n30,
         SubCellInst_SboxInst_13_AND3_U1_n29,
         SubCellInst_SboxInst_13_AND3_U1_n28,
         SubCellInst_SboxInst_13_AND3_U1_n27,
         SubCellInst_SboxInst_13_AND3_U1_n26,
         SubCellInst_SboxInst_13_AND3_U1_n25,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND1_U1_n36,
         SubCellInst_SboxInst_14_AND1_U1_n35,
         SubCellInst_SboxInst_14_AND1_U1_n34,
         SubCellInst_SboxInst_14_AND1_U1_n33,
         SubCellInst_SboxInst_14_AND1_U1_n32,
         SubCellInst_SboxInst_14_AND1_U1_n31,
         SubCellInst_SboxInst_14_AND1_U1_n30,
         SubCellInst_SboxInst_14_AND1_U1_n29,
         SubCellInst_SboxInst_14_AND1_U1_n28,
         SubCellInst_SboxInst_14_AND1_U1_n27,
         SubCellInst_SboxInst_14_AND1_U1_n26,
         SubCellInst_SboxInst_14_AND1_U1_n25,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND3_U1_n36,
         SubCellInst_SboxInst_14_AND3_U1_n35,
         SubCellInst_SboxInst_14_AND3_U1_n34,
         SubCellInst_SboxInst_14_AND3_U1_n33,
         SubCellInst_SboxInst_14_AND3_U1_n32,
         SubCellInst_SboxInst_14_AND3_U1_n31,
         SubCellInst_SboxInst_14_AND3_U1_n30,
         SubCellInst_SboxInst_14_AND3_U1_n29,
         SubCellInst_SboxInst_14_AND3_U1_n28,
         SubCellInst_SboxInst_14_AND3_U1_n27,
         SubCellInst_SboxInst_14_AND3_U1_n26,
         SubCellInst_SboxInst_14_AND3_U1_n25,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND1_U1_n36,
         SubCellInst_SboxInst_15_AND1_U1_n35,
         SubCellInst_SboxInst_15_AND1_U1_n34,
         SubCellInst_SboxInst_15_AND1_U1_n33,
         SubCellInst_SboxInst_15_AND1_U1_n32,
         SubCellInst_SboxInst_15_AND1_U1_n31,
         SubCellInst_SboxInst_15_AND1_U1_n30,
         SubCellInst_SboxInst_15_AND1_U1_n29,
         SubCellInst_SboxInst_15_AND1_U1_n28,
         SubCellInst_SboxInst_15_AND1_U1_n27,
         SubCellInst_SboxInst_15_AND1_U1_n26,
         SubCellInst_SboxInst_15_AND1_U1_n25,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND3_U1_n36,
         SubCellInst_SboxInst_15_AND3_U1_n35,
         SubCellInst_SboxInst_15_AND3_U1_n34,
         SubCellInst_SboxInst_15_AND3_U1_n33,
         SubCellInst_SboxInst_15_AND3_U1_n32,
         SubCellInst_SboxInst_15_AND3_U1_n31,
         SubCellInst_SboxInst_15_AND3_U1_n30,
         SubCellInst_SboxInst_15_AND3_U1_n29,
         SubCellInst_SboxInst_15_AND3_U1_n28,
         SubCellInst_SboxInst_15_AND3_U1_n27,
         SubCellInst_SboxInst_15_AND3_U1_n26,
         SubCellInst_SboxInst_15_AND3_U1_n25,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_0_AND2_U1_n36,
         SubCellInst_SboxInst_0_AND2_U1_n35,
         SubCellInst_SboxInst_0_AND2_U1_n34,
         SubCellInst_SboxInst_0_AND2_U1_n33,
         SubCellInst_SboxInst_0_AND2_U1_n32,
         SubCellInst_SboxInst_0_AND2_U1_n31,
         SubCellInst_SboxInst_0_AND2_U1_n30,
         SubCellInst_SboxInst_0_AND2_U1_n29,
         SubCellInst_SboxInst_0_AND2_U1_n28,
         SubCellInst_SboxInst_0_AND2_U1_n27,
         SubCellInst_SboxInst_0_AND2_U1_n26,
         SubCellInst_SboxInst_0_AND2_U1_n25,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_0_AND4_U1_n36,
         SubCellInst_SboxInst_0_AND4_U1_n35,
         SubCellInst_SboxInst_0_AND4_U1_n34,
         SubCellInst_SboxInst_0_AND4_U1_n33,
         SubCellInst_SboxInst_0_AND4_U1_n32,
         SubCellInst_SboxInst_0_AND4_U1_n31,
         SubCellInst_SboxInst_0_AND4_U1_n30,
         SubCellInst_SboxInst_0_AND4_U1_n29,
         SubCellInst_SboxInst_0_AND4_U1_n28,
         SubCellInst_SboxInst_0_AND4_U1_n27,
         SubCellInst_SboxInst_0_AND4_U1_n26,
         SubCellInst_SboxInst_0_AND4_U1_n25,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND2_U1_n36,
         SubCellInst_SboxInst_1_AND2_U1_n35,
         SubCellInst_SboxInst_1_AND2_U1_n34,
         SubCellInst_SboxInst_1_AND2_U1_n33,
         SubCellInst_SboxInst_1_AND2_U1_n32,
         SubCellInst_SboxInst_1_AND2_U1_n31,
         SubCellInst_SboxInst_1_AND2_U1_n30,
         SubCellInst_SboxInst_1_AND2_U1_n29,
         SubCellInst_SboxInst_1_AND2_U1_n28,
         SubCellInst_SboxInst_1_AND2_U1_n27,
         SubCellInst_SboxInst_1_AND2_U1_n26,
         SubCellInst_SboxInst_1_AND2_U1_n25,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND4_U1_n36,
         SubCellInst_SboxInst_1_AND4_U1_n35,
         SubCellInst_SboxInst_1_AND4_U1_n34,
         SubCellInst_SboxInst_1_AND4_U1_n33,
         SubCellInst_SboxInst_1_AND4_U1_n32,
         SubCellInst_SboxInst_1_AND4_U1_n31,
         SubCellInst_SboxInst_1_AND4_U1_n30,
         SubCellInst_SboxInst_1_AND4_U1_n29,
         SubCellInst_SboxInst_1_AND4_U1_n28,
         SubCellInst_SboxInst_1_AND4_U1_n27,
         SubCellInst_SboxInst_1_AND4_U1_n26,
         SubCellInst_SboxInst_1_AND4_U1_n25,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND2_U1_n36,
         SubCellInst_SboxInst_2_AND2_U1_n35,
         SubCellInst_SboxInst_2_AND2_U1_n34,
         SubCellInst_SboxInst_2_AND2_U1_n33,
         SubCellInst_SboxInst_2_AND2_U1_n32,
         SubCellInst_SboxInst_2_AND2_U1_n31,
         SubCellInst_SboxInst_2_AND2_U1_n30,
         SubCellInst_SboxInst_2_AND2_U1_n29,
         SubCellInst_SboxInst_2_AND2_U1_n28,
         SubCellInst_SboxInst_2_AND2_U1_n27,
         SubCellInst_SboxInst_2_AND2_U1_n26,
         SubCellInst_SboxInst_2_AND2_U1_n25,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND4_U1_n36,
         SubCellInst_SboxInst_2_AND4_U1_n35,
         SubCellInst_SboxInst_2_AND4_U1_n34,
         SubCellInst_SboxInst_2_AND4_U1_n33,
         SubCellInst_SboxInst_2_AND4_U1_n32,
         SubCellInst_SboxInst_2_AND4_U1_n31,
         SubCellInst_SboxInst_2_AND4_U1_n30,
         SubCellInst_SboxInst_2_AND4_U1_n29,
         SubCellInst_SboxInst_2_AND4_U1_n28,
         SubCellInst_SboxInst_2_AND4_U1_n27,
         SubCellInst_SboxInst_2_AND4_U1_n26,
         SubCellInst_SboxInst_2_AND4_U1_n25,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND2_U1_n36,
         SubCellInst_SboxInst_3_AND2_U1_n35,
         SubCellInst_SboxInst_3_AND2_U1_n34,
         SubCellInst_SboxInst_3_AND2_U1_n33,
         SubCellInst_SboxInst_3_AND2_U1_n32,
         SubCellInst_SboxInst_3_AND2_U1_n31,
         SubCellInst_SboxInst_3_AND2_U1_n30,
         SubCellInst_SboxInst_3_AND2_U1_n29,
         SubCellInst_SboxInst_3_AND2_U1_n28,
         SubCellInst_SboxInst_3_AND2_U1_n27,
         SubCellInst_SboxInst_3_AND2_U1_n26,
         SubCellInst_SboxInst_3_AND2_U1_n25,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND4_U1_n36,
         SubCellInst_SboxInst_3_AND4_U1_n35,
         SubCellInst_SboxInst_3_AND4_U1_n34,
         SubCellInst_SboxInst_3_AND4_U1_n33,
         SubCellInst_SboxInst_3_AND4_U1_n32,
         SubCellInst_SboxInst_3_AND4_U1_n31,
         SubCellInst_SboxInst_3_AND4_U1_n30,
         SubCellInst_SboxInst_3_AND4_U1_n29,
         SubCellInst_SboxInst_3_AND4_U1_n28,
         SubCellInst_SboxInst_3_AND4_U1_n27,
         SubCellInst_SboxInst_3_AND4_U1_n26,
         SubCellInst_SboxInst_3_AND4_U1_n25,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND2_U1_n36,
         SubCellInst_SboxInst_4_AND2_U1_n35,
         SubCellInst_SboxInst_4_AND2_U1_n34,
         SubCellInst_SboxInst_4_AND2_U1_n33,
         SubCellInst_SboxInst_4_AND2_U1_n32,
         SubCellInst_SboxInst_4_AND2_U1_n31,
         SubCellInst_SboxInst_4_AND2_U1_n30,
         SubCellInst_SboxInst_4_AND2_U1_n29,
         SubCellInst_SboxInst_4_AND2_U1_n28,
         SubCellInst_SboxInst_4_AND2_U1_n27,
         SubCellInst_SboxInst_4_AND2_U1_n26,
         SubCellInst_SboxInst_4_AND2_U1_n25,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND4_U1_n36,
         SubCellInst_SboxInst_4_AND4_U1_n35,
         SubCellInst_SboxInst_4_AND4_U1_n34,
         SubCellInst_SboxInst_4_AND4_U1_n33,
         SubCellInst_SboxInst_4_AND4_U1_n32,
         SubCellInst_SboxInst_4_AND4_U1_n31,
         SubCellInst_SboxInst_4_AND4_U1_n30,
         SubCellInst_SboxInst_4_AND4_U1_n29,
         SubCellInst_SboxInst_4_AND4_U1_n28,
         SubCellInst_SboxInst_4_AND4_U1_n27,
         SubCellInst_SboxInst_4_AND4_U1_n26,
         SubCellInst_SboxInst_4_AND4_U1_n25,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND2_U1_n36,
         SubCellInst_SboxInst_5_AND2_U1_n35,
         SubCellInst_SboxInst_5_AND2_U1_n34,
         SubCellInst_SboxInst_5_AND2_U1_n33,
         SubCellInst_SboxInst_5_AND2_U1_n32,
         SubCellInst_SboxInst_5_AND2_U1_n31,
         SubCellInst_SboxInst_5_AND2_U1_n30,
         SubCellInst_SboxInst_5_AND2_U1_n29,
         SubCellInst_SboxInst_5_AND2_U1_n28,
         SubCellInst_SboxInst_5_AND2_U1_n27,
         SubCellInst_SboxInst_5_AND2_U1_n26,
         SubCellInst_SboxInst_5_AND2_U1_n25,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND4_U1_n36,
         SubCellInst_SboxInst_5_AND4_U1_n35,
         SubCellInst_SboxInst_5_AND4_U1_n34,
         SubCellInst_SboxInst_5_AND4_U1_n33,
         SubCellInst_SboxInst_5_AND4_U1_n32,
         SubCellInst_SboxInst_5_AND4_U1_n31,
         SubCellInst_SboxInst_5_AND4_U1_n30,
         SubCellInst_SboxInst_5_AND4_U1_n29,
         SubCellInst_SboxInst_5_AND4_U1_n28,
         SubCellInst_SboxInst_5_AND4_U1_n27,
         SubCellInst_SboxInst_5_AND4_U1_n26,
         SubCellInst_SboxInst_5_AND4_U1_n25,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND2_U1_n36,
         SubCellInst_SboxInst_6_AND2_U1_n35,
         SubCellInst_SboxInst_6_AND2_U1_n34,
         SubCellInst_SboxInst_6_AND2_U1_n33,
         SubCellInst_SboxInst_6_AND2_U1_n32,
         SubCellInst_SboxInst_6_AND2_U1_n31,
         SubCellInst_SboxInst_6_AND2_U1_n30,
         SubCellInst_SboxInst_6_AND2_U1_n29,
         SubCellInst_SboxInst_6_AND2_U1_n28,
         SubCellInst_SboxInst_6_AND2_U1_n27,
         SubCellInst_SboxInst_6_AND2_U1_n26,
         SubCellInst_SboxInst_6_AND2_U1_n25,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND4_U1_n36,
         SubCellInst_SboxInst_6_AND4_U1_n35,
         SubCellInst_SboxInst_6_AND4_U1_n34,
         SubCellInst_SboxInst_6_AND4_U1_n33,
         SubCellInst_SboxInst_6_AND4_U1_n32,
         SubCellInst_SboxInst_6_AND4_U1_n31,
         SubCellInst_SboxInst_6_AND4_U1_n30,
         SubCellInst_SboxInst_6_AND4_U1_n29,
         SubCellInst_SboxInst_6_AND4_U1_n28,
         SubCellInst_SboxInst_6_AND4_U1_n27,
         SubCellInst_SboxInst_6_AND4_U1_n26,
         SubCellInst_SboxInst_6_AND4_U1_n25,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND2_U1_n36,
         SubCellInst_SboxInst_7_AND2_U1_n35,
         SubCellInst_SboxInst_7_AND2_U1_n34,
         SubCellInst_SboxInst_7_AND2_U1_n33,
         SubCellInst_SboxInst_7_AND2_U1_n32,
         SubCellInst_SboxInst_7_AND2_U1_n31,
         SubCellInst_SboxInst_7_AND2_U1_n30,
         SubCellInst_SboxInst_7_AND2_U1_n29,
         SubCellInst_SboxInst_7_AND2_U1_n28,
         SubCellInst_SboxInst_7_AND2_U1_n27,
         SubCellInst_SboxInst_7_AND2_U1_n26,
         SubCellInst_SboxInst_7_AND2_U1_n25,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND4_U1_n36,
         SubCellInst_SboxInst_7_AND4_U1_n35,
         SubCellInst_SboxInst_7_AND4_U1_n34,
         SubCellInst_SboxInst_7_AND4_U1_n33,
         SubCellInst_SboxInst_7_AND4_U1_n32,
         SubCellInst_SboxInst_7_AND4_U1_n31,
         SubCellInst_SboxInst_7_AND4_U1_n30,
         SubCellInst_SboxInst_7_AND4_U1_n29,
         SubCellInst_SboxInst_7_AND4_U1_n28,
         SubCellInst_SboxInst_7_AND4_U1_n27,
         SubCellInst_SboxInst_7_AND4_U1_n26,
         SubCellInst_SboxInst_7_AND4_U1_n25,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND2_U1_n36,
         SubCellInst_SboxInst_8_AND2_U1_n35,
         SubCellInst_SboxInst_8_AND2_U1_n34,
         SubCellInst_SboxInst_8_AND2_U1_n33,
         SubCellInst_SboxInst_8_AND2_U1_n32,
         SubCellInst_SboxInst_8_AND2_U1_n31,
         SubCellInst_SboxInst_8_AND2_U1_n30,
         SubCellInst_SboxInst_8_AND2_U1_n29,
         SubCellInst_SboxInst_8_AND2_U1_n28,
         SubCellInst_SboxInst_8_AND2_U1_n27,
         SubCellInst_SboxInst_8_AND2_U1_n26,
         SubCellInst_SboxInst_8_AND2_U1_n25,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND4_U1_n36,
         SubCellInst_SboxInst_8_AND4_U1_n35,
         SubCellInst_SboxInst_8_AND4_U1_n34,
         SubCellInst_SboxInst_8_AND4_U1_n33,
         SubCellInst_SboxInst_8_AND4_U1_n32,
         SubCellInst_SboxInst_8_AND4_U1_n31,
         SubCellInst_SboxInst_8_AND4_U1_n30,
         SubCellInst_SboxInst_8_AND4_U1_n29,
         SubCellInst_SboxInst_8_AND4_U1_n28,
         SubCellInst_SboxInst_8_AND4_U1_n27,
         SubCellInst_SboxInst_8_AND4_U1_n26,
         SubCellInst_SboxInst_8_AND4_U1_n25,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND2_U1_n36,
         SubCellInst_SboxInst_9_AND2_U1_n35,
         SubCellInst_SboxInst_9_AND2_U1_n34,
         SubCellInst_SboxInst_9_AND2_U1_n33,
         SubCellInst_SboxInst_9_AND2_U1_n32,
         SubCellInst_SboxInst_9_AND2_U1_n31,
         SubCellInst_SboxInst_9_AND2_U1_n30,
         SubCellInst_SboxInst_9_AND2_U1_n29,
         SubCellInst_SboxInst_9_AND2_U1_n28,
         SubCellInst_SboxInst_9_AND2_U1_n27,
         SubCellInst_SboxInst_9_AND2_U1_n26,
         SubCellInst_SboxInst_9_AND2_U1_n25,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND4_U1_n36,
         SubCellInst_SboxInst_9_AND4_U1_n35,
         SubCellInst_SboxInst_9_AND4_U1_n34,
         SubCellInst_SboxInst_9_AND4_U1_n33,
         SubCellInst_SboxInst_9_AND4_U1_n32,
         SubCellInst_SboxInst_9_AND4_U1_n31,
         SubCellInst_SboxInst_9_AND4_U1_n30,
         SubCellInst_SboxInst_9_AND4_U1_n29,
         SubCellInst_SboxInst_9_AND4_U1_n28,
         SubCellInst_SboxInst_9_AND4_U1_n27,
         SubCellInst_SboxInst_9_AND4_U1_n26,
         SubCellInst_SboxInst_9_AND4_U1_n25,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND2_U1_n36,
         SubCellInst_SboxInst_10_AND2_U1_n35,
         SubCellInst_SboxInst_10_AND2_U1_n34,
         SubCellInst_SboxInst_10_AND2_U1_n33,
         SubCellInst_SboxInst_10_AND2_U1_n32,
         SubCellInst_SboxInst_10_AND2_U1_n31,
         SubCellInst_SboxInst_10_AND2_U1_n30,
         SubCellInst_SboxInst_10_AND2_U1_n29,
         SubCellInst_SboxInst_10_AND2_U1_n28,
         SubCellInst_SboxInst_10_AND2_U1_n27,
         SubCellInst_SboxInst_10_AND2_U1_n26,
         SubCellInst_SboxInst_10_AND2_U1_n25,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND4_U1_n36,
         SubCellInst_SboxInst_10_AND4_U1_n35,
         SubCellInst_SboxInst_10_AND4_U1_n34,
         SubCellInst_SboxInst_10_AND4_U1_n33,
         SubCellInst_SboxInst_10_AND4_U1_n32,
         SubCellInst_SboxInst_10_AND4_U1_n31,
         SubCellInst_SboxInst_10_AND4_U1_n30,
         SubCellInst_SboxInst_10_AND4_U1_n29,
         SubCellInst_SboxInst_10_AND4_U1_n28,
         SubCellInst_SboxInst_10_AND4_U1_n27,
         SubCellInst_SboxInst_10_AND4_U1_n26,
         SubCellInst_SboxInst_10_AND4_U1_n25,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND2_U1_n36,
         SubCellInst_SboxInst_11_AND2_U1_n35,
         SubCellInst_SboxInst_11_AND2_U1_n34,
         SubCellInst_SboxInst_11_AND2_U1_n33,
         SubCellInst_SboxInst_11_AND2_U1_n32,
         SubCellInst_SboxInst_11_AND2_U1_n31,
         SubCellInst_SboxInst_11_AND2_U1_n30,
         SubCellInst_SboxInst_11_AND2_U1_n29,
         SubCellInst_SboxInst_11_AND2_U1_n28,
         SubCellInst_SboxInst_11_AND2_U1_n27,
         SubCellInst_SboxInst_11_AND2_U1_n26,
         SubCellInst_SboxInst_11_AND2_U1_n25,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND4_U1_n36,
         SubCellInst_SboxInst_11_AND4_U1_n35,
         SubCellInst_SboxInst_11_AND4_U1_n34,
         SubCellInst_SboxInst_11_AND4_U1_n33,
         SubCellInst_SboxInst_11_AND4_U1_n32,
         SubCellInst_SboxInst_11_AND4_U1_n31,
         SubCellInst_SboxInst_11_AND4_U1_n30,
         SubCellInst_SboxInst_11_AND4_U1_n29,
         SubCellInst_SboxInst_11_AND4_U1_n28,
         SubCellInst_SboxInst_11_AND4_U1_n27,
         SubCellInst_SboxInst_11_AND4_U1_n26,
         SubCellInst_SboxInst_11_AND4_U1_n25,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND2_U1_n36,
         SubCellInst_SboxInst_12_AND2_U1_n35,
         SubCellInst_SboxInst_12_AND2_U1_n34,
         SubCellInst_SboxInst_12_AND2_U1_n33,
         SubCellInst_SboxInst_12_AND2_U1_n32,
         SubCellInst_SboxInst_12_AND2_U1_n31,
         SubCellInst_SboxInst_12_AND2_U1_n30,
         SubCellInst_SboxInst_12_AND2_U1_n29,
         SubCellInst_SboxInst_12_AND2_U1_n28,
         SubCellInst_SboxInst_12_AND2_U1_n27,
         SubCellInst_SboxInst_12_AND2_U1_n26,
         SubCellInst_SboxInst_12_AND2_U1_n25,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND4_U1_n36,
         SubCellInst_SboxInst_12_AND4_U1_n35,
         SubCellInst_SboxInst_12_AND4_U1_n34,
         SubCellInst_SboxInst_12_AND4_U1_n33,
         SubCellInst_SboxInst_12_AND4_U1_n32,
         SubCellInst_SboxInst_12_AND4_U1_n31,
         SubCellInst_SboxInst_12_AND4_U1_n30,
         SubCellInst_SboxInst_12_AND4_U1_n29,
         SubCellInst_SboxInst_12_AND4_U1_n28,
         SubCellInst_SboxInst_12_AND4_U1_n27,
         SubCellInst_SboxInst_12_AND4_U1_n26,
         SubCellInst_SboxInst_12_AND4_U1_n25,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND2_U1_n36,
         SubCellInst_SboxInst_13_AND2_U1_n35,
         SubCellInst_SboxInst_13_AND2_U1_n34,
         SubCellInst_SboxInst_13_AND2_U1_n33,
         SubCellInst_SboxInst_13_AND2_U1_n32,
         SubCellInst_SboxInst_13_AND2_U1_n31,
         SubCellInst_SboxInst_13_AND2_U1_n30,
         SubCellInst_SboxInst_13_AND2_U1_n29,
         SubCellInst_SboxInst_13_AND2_U1_n28,
         SubCellInst_SboxInst_13_AND2_U1_n27,
         SubCellInst_SboxInst_13_AND2_U1_n26,
         SubCellInst_SboxInst_13_AND2_U1_n25,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND4_U1_n36,
         SubCellInst_SboxInst_13_AND4_U1_n35,
         SubCellInst_SboxInst_13_AND4_U1_n34,
         SubCellInst_SboxInst_13_AND4_U1_n33,
         SubCellInst_SboxInst_13_AND4_U1_n32,
         SubCellInst_SboxInst_13_AND4_U1_n31,
         SubCellInst_SboxInst_13_AND4_U1_n30,
         SubCellInst_SboxInst_13_AND4_U1_n29,
         SubCellInst_SboxInst_13_AND4_U1_n28,
         SubCellInst_SboxInst_13_AND4_U1_n27,
         SubCellInst_SboxInst_13_AND4_U1_n26,
         SubCellInst_SboxInst_13_AND4_U1_n25,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND2_U1_n36,
         SubCellInst_SboxInst_14_AND2_U1_n35,
         SubCellInst_SboxInst_14_AND2_U1_n34,
         SubCellInst_SboxInst_14_AND2_U1_n33,
         SubCellInst_SboxInst_14_AND2_U1_n32,
         SubCellInst_SboxInst_14_AND2_U1_n31,
         SubCellInst_SboxInst_14_AND2_U1_n30,
         SubCellInst_SboxInst_14_AND2_U1_n29,
         SubCellInst_SboxInst_14_AND2_U1_n28,
         SubCellInst_SboxInst_14_AND2_U1_n27,
         SubCellInst_SboxInst_14_AND2_U1_n26,
         SubCellInst_SboxInst_14_AND2_U1_n25,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND4_U1_n36,
         SubCellInst_SboxInst_14_AND4_U1_n35,
         SubCellInst_SboxInst_14_AND4_U1_n34,
         SubCellInst_SboxInst_14_AND4_U1_n33,
         SubCellInst_SboxInst_14_AND4_U1_n32,
         SubCellInst_SboxInst_14_AND4_U1_n31,
         SubCellInst_SboxInst_14_AND4_U1_n30,
         SubCellInst_SboxInst_14_AND4_U1_n29,
         SubCellInst_SboxInst_14_AND4_U1_n28,
         SubCellInst_SboxInst_14_AND4_U1_n27,
         SubCellInst_SboxInst_14_AND4_U1_n26,
         SubCellInst_SboxInst_14_AND4_U1_n25,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND2_U1_n36,
         SubCellInst_SboxInst_15_AND2_U1_n35,
         SubCellInst_SboxInst_15_AND2_U1_n34,
         SubCellInst_SboxInst_15_AND2_U1_n33,
         SubCellInst_SboxInst_15_AND2_U1_n32,
         SubCellInst_SboxInst_15_AND2_U1_n31,
         SubCellInst_SboxInst_15_AND2_U1_n30,
         SubCellInst_SboxInst_15_AND2_U1_n29,
         SubCellInst_SboxInst_15_AND2_U1_n28,
         SubCellInst_SboxInst_15_AND2_U1_n27,
         SubCellInst_SboxInst_15_AND2_U1_n26,
         SubCellInst_SboxInst_15_AND2_U1_n25,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND4_U1_n36,
         SubCellInst_SboxInst_15_AND4_U1_n35,
         SubCellInst_SboxInst_15_AND4_U1_n34,
         SubCellInst_SboxInst_15_AND4_U1_n33,
         SubCellInst_SboxInst_15_AND4_U1_n32,
         SubCellInst_SboxInst_15_AND4_U1_n31,
         SubCellInst_SboxInst_15_AND4_U1_n30,
         SubCellInst_SboxInst_15_AND4_U1_n29,
         SubCellInst_SboxInst_15_AND4_U1_n28,
         SubCellInst_SboxInst_15_AND4_U1_n27,
         SubCellInst_SboxInst_15_AND4_U1_n26,
         SubCellInst_SboxInst_15_AND4_U1_n25,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND4_U1_a_reg_2_;
  wire   [63:0] TweakeyGeneration_StateRegInput;
  wire   [63:0] TweakeyGeneration_key_Feedback;
  wire   [4:1] FSMUpdate;
  wire   [5:0] FSMSelected;
  wire   [5:4] FSM;
  wire   [63:0] StateRegInput;
  wire   [63:0] MCOutput;
  wire   [47:0] ShiftRowsOutput;
  wire   [63:32] AddRoundConstantOutput;
  wire   [63:60] SubCellOutput;
  wire   [2:0] SubCellInst_SboxInst_0_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_0_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_0_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_0_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_0_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_0_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_1_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_1_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_1_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_1_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_1_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_1_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_2_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_2_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_2_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_2_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_2_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_2_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_3_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_3_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_3_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_3_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_3_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_3_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_4_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_4_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_4_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_4_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_4_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_4_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_5_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_5_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_5_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_5_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_5_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_5_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_6_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_6_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_6_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_6_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_6_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_6_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_7_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_7_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_7_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_7_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_7_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_7_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_8_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_8_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_8_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_8_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_8_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_8_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_9_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_9_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_9_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_9_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_9_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_9_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_10_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_10_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_10_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_10_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_10_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_10_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_11_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_11_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_11_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_11_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_11_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_11_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_12_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_12_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_12_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_12_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_12_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_12_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_13_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_13_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_13_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_13_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_13_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_13_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_14_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_14_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_14_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_14_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_14_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_14_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_15_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_15_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_15_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_15_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_15_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_15_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_0_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_0_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_0_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_0_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_0_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_0_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_1_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_1_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_1_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_1_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_1_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_1_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_2_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_2_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_2_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_2_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_2_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_2_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_3_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_3_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_3_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_3_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_3_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_3_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_4_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_4_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_4_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_4_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_4_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_4_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_5_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_5_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_5_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_5_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_5_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_5_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_6_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_6_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_6_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_6_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_6_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_6_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_7_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_7_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_7_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_7_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_7_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_7_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_8_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_8_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_8_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_8_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_8_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_8_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_9_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_9_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_9_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_9_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_9_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_9_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_10_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_10_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_10_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_10_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_10_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_10_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_11_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_11_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_11_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_11_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_11_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_11_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_12_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_12_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_12_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_12_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_12_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_12_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_13_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_13_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_13_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_13_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_13_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_13_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_14_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_14_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_14_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_14_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_14_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_14_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_15_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_15_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_15_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_15_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_15_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_15_AND4_U1_mul;

  DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .D(FSMSelected[3]), .CK(
        clk_gated), .Q(FSMUpdate[4]), .QN(n16) );
  DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .D(FSMSelected[4]), .CK(
        clk_gated), .Q(FSM[4]), .QN(n14) );
  DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .D(FSMSelected[1]), .CK(
        clk_gated), .Q(FSM_1), .QN(n15) );
  DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .D(FSMSelected[0]), .CK(
        clk_gated), .Q(FSMUpdate[1]), .QN(n18) );
  DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .D(FSMSelected[5]), .CK(
        clk_gated), .Q(FSM[5]), .QN(n13) );
  DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .D(FSMSelected[2]), .CK(
        clk_gated), .Q(FSMUpdate[3]), .QN(n17) );
  INV_X1 U39 ( .A(rst), .ZN(n30) );
  NAND3_X1 U40 ( .A1(n16), .A2(n17), .A3(FSM_1), .ZN(n36) );
  NOR2_X1 U41 ( .A1(n18), .A2(n36), .ZN(n31) );
  OAI21_X1 U42 ( .B1(n13), .B2(n31), .A(n14), .ZN(n32) );
  OAI211_X1 U43 ( .C1(n13), .C2(n14), .A(n30), .B(n32), .ZN(FSMSelected[0]) );
  NOR2_X1 U44 ( .A1(rst), .A2(n18), .ZN(FSMSelected[1]) );
  NOR2_X1 U45 ( .A1(rst), .A2(n16), .ZN(FSMSelected[4]) );
  NOR2_X1 U46 ( .A1(rst), .A2(n17), .ZN(FSMSelected[3]) );
  NOR2_X1 U47 ( .A1(FSMSelected[4]), .A2(FSMSelected[3]), .ZN(n35) );
  NAND2_X1 U48 ( .A1(n14), .A2(FSM[5]), .ZN(n33) );
  OAI21_X1 U49 ( .B1(n18), .B2(n33), .A(n30), .ZN(n34) );
  AOI21_X1 U50 ( .B1(n35), .B2(n34), .A(n15), .ZN(FSMSelected[2]) );
  NAND2_X1 U51 ( .A1(FSMSelected[1]), .A2(FSM[5]), .ZN(n37) );
  OAI22_X1 U52 ( .A1(rst), .A2(n14), .B1(n37), .B2(n36), .ZN(FSMSelected[5])
         );
  NAND4_X1 U53 ( .A1(n15), .A2(n16), .A3(n17), .A4(FSM[5]), .ZN(n38) );
  NOR3_X1 U54 ( .A1(n14), .A2(n18), .A3(n38), .ZN(done) );
  INV_X1 SubCellInst_SboxInst_0_U1_U1 ( .A(Ciphertext_s0[2]), .ZN(
        SubCellInst_SboxInst_0_n3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[2]), 
        .B(Ciphertext_s0[3]), .Z(SubCellInst_SboxInst_0_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[2]), 
        .B(Ciphertext_s1[3]), .Z(new_AGEMA_signal_1170) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[2]), 
        .B(Ciphertext_s2[3]), .Z(new_AGEMA_signal_1171) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[0]), 
        .B(Ciphertext_s0[2]), .Z(SubCellInst_SboxInst_0_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[0]), 
        .B(Ciphertext_s1[2]), .Z(new_AGEMA_signal_1174) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[0]), 
        .B(Ciphertext_s2[2]), .Z(new_AGEMA_signal_1175) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_XX_2_), .Z(SubCellInst_SboxInst_0_Q0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        new_AGEMA_signal_1174), .Z(new_AGEMA_signal_1742) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        new_AGEMA_signal_1175), .Z(new_AGEMA_signal_1743) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_XX_1_), .Z(SubCellInst_SboxInst_0_Q1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        new_AGEMA_signal_1170), .Z(new_AGEMA_signal_1744) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        new_AGEMA_signal_1171), .Z(new_AGEMA_signal_1745) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_n3), .ZN(SubCellInst_SboxInst_0_Q4) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        Ciphertext_s1[2]), .Z(new_AGEMA_signal_1746) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        Ciphertext_s2[2]), .Z(new_AGEMA_signal_1747) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_XX_2_), .B(SubCellInst_SboxInst_0_n3), .Z(
        SubCellInst_SboxInst_0_Q6) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1174), 
        .B(Ciphertext_s1[2]), .Z(new_AGEMA_signal_1748) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1175), 
        .B(Ciphertext_s2[2]), .Z(new_AGEMA_signal_1749) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_0_Q1), .B(SubCellInst_SboxInst_0_Q6), .ZN(
        SubCellInst_SboxInst_0_L1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1744), 
        .B(new_AGEMA_signal_1748), .Z(new_AGEMA_signal_1936) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1745), 
        .B(new_AGEMA_signal_1749), .Z(new_AGEMA_signal_1937) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_n3), .Z(SubCellInst_SboxInst_0_L2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        Ciphertext_s1[2]), .Z(new_AGEMA_signal_1750) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        Ciphertext_s2[2]), .Z(new_AGEMA_signal_1751) );
  INV_X1 SubCellInst_SboxInst_1_U1_U1 ( .A(Ciphertext_s0[6]), .ZN(
        SubCellInst_SboxInst_1_n3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[6]), 
        .B(Ciphertext_s0[7]), .Z(SubCellInst_SboxInst_1_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[6]), 
        .B(Ciphertext_s1[7]), .Z(new_AGEMA_signal_1182) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[6]), 
        .B(Ciphertext_s2[7]), .Z(new_AGEMA_signal_1183) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[4]), 
        .B(Ciphertext_s0[6]), .Z(SubCellInst_SboxInst_1_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[4]), 
        .B(Ciphertext_s1[6]), .Z(new_AGEMA_signal_1186) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[4]), 
        .B(Ciphertext_s2[6]), .Z(new_AGEMA_signal_1187) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_XX_2_), .Z(SubCellInst_SboxInst_1_Q0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        new_AGEMA_signal_1186), .Z(new_AGEMA_signal_1754) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        new_AGEMA_signal_1187), .Z(new_AGEMA_signal_1755) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_XX_1_), .Z(SubCellInst_SboxInst_1_Q1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        new_AGEMA_signal_1182), .Z(new_AGEMA_signal_1756) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        new_AGEMA_signal_1183), .Z(new_AGEMA_signal_1757) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_n3), .ZN(SubCellInst_SboxInst_1_Q4) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        Ciphertext_s1[6]), .Z(new_AGEMA_signal_1758) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        Ciphertext_s2[6]), .Z(new_AGEMA_signal_1759) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_XX_2_), .B(SubCellInst_SboxInst_1_n3), .Z(
        SubCellInst_SboxInst_1_Q6) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1186), 
        .B(Ciphertext_s1[6]), .Z(new_AGEMA_signal_1760) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1187), 
        .B(Ciphertext_s2[6]), .Z(new_AGEMA_signal_1761) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_1_Q1), .B(SubCellInst_SboxInst_1_Q6), .ZN(
        SubCellInst_SboxInst_1_L1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1756), 
        .B(new_AGEMA_signal_1760), .Z(new_AGEMA_signal_1942) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1757), 
        .B(new_AGEMA_signal_1761), .Z(new_AGEMA_signal_1943) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_n3), .Z(SubCellInst_SboxInst_1_L2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        Ciphertext_s1[6]), .Z(new_AGEMA_signal_1762) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        Ciphertext_s2[6]), .Z(new_AGEMA_signal_1763) );
  INV_X1 SubCellInst_SboxInst_2_U1_U1 ( .A(Ciphertext_s0[10]), .ZN(
        SubCellInst_SboxInst_2_n3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[10]), 
        .B(Ciphertext_s0[11]), .Z(SubCellInst_SboxInst_2_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[10]), 
        .B(Ciphertext_s1[11]), .Z(new_AGEMA_signal_1194) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[10]), 
        .B(Ciphertext_s2[11]), .Z(new_AGEMA_signal_1195) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[8]), 
        .B(Ciphertext_s0[10]), .Z(SubCellInst_SboxInst_2_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[8]), 
        .B(Ciphertext_s1[10]), .Z(new_AGEMA_signal_1198) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[8]), 
        .B(Ciphertext_s2[10]), .Z(new_AGEMA_signal_1199) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_XX_2_), .Z(SubCellInst_SboxInst_2_Q0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        new_AGEMA_signal_1198), .Z(new_AGEMA_signal_1766) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        new_AGEMA_signal_1199), .Z(new_AGEMA_signal_1767) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_XX_1_), .Z(SubCellInst_SboxInst_2_Q1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        new_AGEMA_signal_1194), .Z(new_AGEMA_signal_1768) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        new_AGEMA_signal_1195), .Z(new_AGEMA_signal_1769) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_n3), .ZN(SubCellInst_SboxInst_2_Q4) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        Ciphertext_s1[10]), .Z(new_AGEMA_signal_1770) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        Ciphertext_s2[10]), .Z(new_AGEMA_signal_1771) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_XX_2_), .B(SubCellInst_SboxInst_2_n3), .Z(
        SubCellInst_SboxInst_2_Q6) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1198), 
        .B(Ciphertext_s1[10]), .Z(new_AGEMA_signal_1772) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1199), 
        .B(Ciphertext_s2[10]), .Z(new_AGEMA_signal_1773) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_2_Q1), .B(SubCellInst_SboxInst_2_Q6), .ZN(
        SubCellInst_SboxInst_2_L1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1768), 
        .B(new_AGEMA_signal_1772), .Z(new_AGEMA_signal_1948) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1769), 
        .B(new_AGEMA_signal_1773), .Z(new_AGEMA_signal_1949) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_n3), .Z(SubCellInst_SboxInst_2_L2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        Ciphertext_s1[10]), .Z(new_AGEMA_signal_1774) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        Ciphertext_s2[10]), .Z(new_AGEMA_signal_1775) );
  INV_X1 SubCellInst_SboxInst_3_U1_U1 ( .A(Ciphertext_s0[14]), .ZN(
        SubCellInst_SboxInst_3_n3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[14]), 
        .B(Ciphertext_s0[15]), .Z(SubCellInst_SboxInst_3_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[14]), 
        .B(Ciphertext_s1[15]), .Z(new_AGEMA_signal_1206) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[14]), 
        .B(Ciphertext_s2[15]), .Z(new_AGEMA_signal_1207) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[12]), 
        .B(Ciphertext_s0[14]), .Z(SubCellInst_SboxInst_3_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[12]), 
        .B(Ciphertext_s1[14]), .Z(new_AGEMA_signal_1210) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[12]), 
        .B(Ciphertext_s2[14]), .Z(new_AGEMA_signal_1211) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_XX_2_), .Z(SubCellInst_SboxInst_3_Q0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        new_AGEMA_signal_1210), .Z(new_AGEMA_signal_1778) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        new_AGEMA_signal_1211), .Z(new_AGEMA_signal_1779) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_XX_1_), .Z(SubCellInst_SboxInst_3_Q1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        new_AGEMA_signal_1206), .Z(new_AGEMA_signal_1780) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        new_AGEMA_signal_1207), .Z(new_AGEMA_signal_1781) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_n3), .ZN(SubCellInst_SboxInst_3_Q4) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        Ciphertext_s1[14]), .Z(new_AGEMA_signal_1782) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        Ciphertext_s2[14]), .Z(new_AGEMA_signal_1783) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_XX_2_), .B(SubCellInst_SboxInst_3_n3), .Z(
        SubCellInst_SboxInst_3_Q6) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1210), 
        .B(Ciphertext_s1[14]), .Z(new_AGEMA_signal_1784) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1211), 
        .B(Ciphertext_s2[14]), .Z(new_AGEMA_signal_1785) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_3_Q1), .B(SubCellInst_SboxInst_3_Q6), .ZN(
        SubCellInst_SboxInst_3_L1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1780), 
        .B(new_AGEMA_signal_1784), .Z(new_AGEMA_signal_1954) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1781), 
        .B(new_AGEMA_signal_1785), .Z(new_AGEMA_signal_1955) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_n3), .Z(SubCellInst_SboxInst_3_L2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        Ciphertext_s1[14]), .Z(new_AGEMA_signal_1786) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        Ciphertext_s2[14]), .Z(new_AGEMA_signal_1787) );
  INV_X1 SubCellInst_SboxInst_4_U1_U1 ( .A(Ciphertext_s0[18]), .ZN(
        SubCellInst_SboxInst_4_n3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[18]), 
        .B(Ciphertext_s0[19]), .Z(SubCellInst_SboxInst_4_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[18]), 
        .B(Ciphertext_s1[19]), .Z(new_AGEMA_signal_1218) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[18]), 
        .B(Ciphertext_s2[19]), .Z(new_AGEMA_signal_1219) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[16]), 
        .B(Ciphertext_s0[18]), .Z(SubCellInst_SboxInst_4_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[16]), 
        .B(Ciphertext_s1[18]), .Z(new_AGEMA_signal_1222) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[16]), 
        .B(Ciphertext_s2[18]), .Z(new_AGEMA_signal_1223) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_XX_2_), .Z(SubCellInst_SboxInst_4_Q0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        new_AGEMA_signal_1222), .Z(new_AGEMA_signal_1790) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        new_AGEMA_signal_1223), .Z(new_AGEMA_signal_1791) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_XX_1_), .Z(SubCellInst_SboxInst_4_Q1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        new_AGEMA_signal_1218), .Z(new_AGEMA_signal_1792) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        new_AGEMA_signal_1219), .Z(new_AGEMA_signal_1793) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_n3), .ZN(SubCellInst_SboxInst_4_Q4) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        Ciphertext_s1[18]), .Z(new_AGEMA_signal_1794) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        Ciphertext_s2[18]), .Z(new_AGEMA_signal_1795) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_XX_2_), .B(SubCellInst_SboxInst_4_n3), .Z(
        SubCellInst_SboxInst_4_Q6) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1222), 
        .B(Ciphertext_s1[18]), .Z(new_AGEMA_signal_1796) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1223), 
        .B(Ciphertext_s2[18]), .Z(new_AGEMA_signal_1797) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_4_Q1), .B(SubCellInst_SboxInst_4_Q6), .ZN(
        SubCellInst_SboxInst_4_L1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1792), 
        .B(new_AGEMA_signal_1796), .Z(new_AGEMA_signal_1960) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1793), 
        .B(new_AGEMA_signal_1797), .Z(new_AGEMA_signal_1961) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_n3), .Z(SubCellInst_SboxInst_4_L2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        Ciphertext_s1[18]), .Z(new_AGEMA_signal_1798) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        Ciphertext_s2[18]), .Z(new_AGEMA_signal_1799) );
  INV_X1 SubCellInst_SboxInst_5_U1_U1 ( .A(Ciphertext_s0[22]), .ZN(
        SubCellInst_SboxInst_5_n3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[22]), 
        .B(Ciphertext_s0[23]), .Z(SubCellInst_SboxInst_5_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[22]), 
        .B(Ciphertext_s1[23]), .Z(new_AGEMA_signal_1230) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[22]), 
        .B(Ciphertext_s2[23]), .Z(new_AGEMA_signal_1231) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[20]), 
        .B(Ciphertext_s0[22]), .Z(SubCellInst_SboxInst_5_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[20]), 
        .B(Ciphertext_s1[22]), .Z(new_AGEMA_signal_1234) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[20]), 
        .B(Ciphertext_s2[22]), .Z(new_AGEMA_signal_1235) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_XX_2_), .Z(SubCellInst_SboxInst_5_Q0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        new_AGEMA_signal_1234), .Z(new_AGEMA_signal_1802) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        new_AGEMA_signal_1235), .Z(new_AGEMA_signal_1803) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_XX_1_), .Z(SubCellInst_SboxInst_5_Q1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        new_AGEMA_signal_1230), .Z(new_AGEMA_signal_1804) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        new_AGEMA_signal_1231), .Z(new_AGEMA_signal_1805) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_n3), .ZN(SubCellInst_SboxInst_5_Q4) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        Ciphertext_s1[22]), .Z(new_AGEMA_signal_1806) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        Ciphertext_s2[22]), .Z(new_AGEMA_signal_1807) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_XX_2_), .B(SubCellInst_SboxInst_5_n3), .Z(
        SubCellInst_SboxInst_5_Q6) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1234), 
        .B(Ciphertext_s1[22]), .Z(new_AGEMA_signal_1808) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1235), 
        .B(Ciphertext_s2[22]), .Z(new_AGEMA_signal_1809) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_5_Q1), .B(SubCellInst_SboxInst_5_Q6), .ZN(
        SubCellInst_SboxInst_5_L1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1804), 
        .B(new_AGEMA_signal_1808), .Z(new_AGEMA_signal_1966) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1805), 
        .B(new_AGEMA_signal_1809), .Z(new_AGEMA_signal_1967) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_n3), .Z(SubCellInst_SboxInst_5_L2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        Ciphertext_s1[22]), .Z(new_AGEMA_signal_1810) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        Ciphertext_s2[22]), .Z(new_AGEMA_signal_1811) );
  INV_X1 SubCellInst_SboxInst_6_U1_U1 ( .A(Ciphertext_s0[26]), .ZN(
        SubCellInst_SboxInst_6_n3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[26]), 
        .B(Ciphertext_s0[27]), .Z(SubCellInst_SboxInst_6_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[26]), 
        .B(Ciphertext_s1[27]), .Z(new_AGEMA_signal_1242) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[26]), 
        .B(Ciphertext_s2[27]), .Z(new_AGEMA_signal_1243) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[24]), 
        .B(Ciphertext_s0[26]), .Z(SubCellInst_SboxInst_6_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[24]), 
        .B(Ciphertext_s1[26]), .Z(new_AGEMA_signal_1246) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[24]), 
        .B(Ciphertext_s2[26]), .Z(new_AGEMA_signal_1247) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_XX_2_), .Z(SubCellInst_SboxInst_6_Q0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        new_AGEMA_signal_1246), .Z(new_AGEMA_signal_1814) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        new_AGEMA_signal_1247), .Z(new_AGEMA_signal_1815) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_XX_1_), .Z(SubCellInst_SboxInst_6_Q1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        new_AGEMA_signal_1242), .Z(new_AGEMA_signal_1816) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        new_AGEMA_signal_1243), .Z(new_AGEMA_signal_1817) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_n3), .ZN(SubCellInst_SboxInst_6_Q4) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        Ciphertext_s1[26]), .Z(new_AGEMA_signal_1818) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        Ciphertext_s2[26]), .Z(new_AGEMA_signal_1819) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_XX_2_), .B(SubCellInst_SboxInst_6_n3), .Z(
        SubCellInst_SboxInst_6_Q6) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1246), 
        .B(Ciphertext_s1[26]), .Z(new_AGEMA_signal_1820) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1247), 
        .B(Ciphertext_s2[26]), .Z(new_AGEMA_signal_1821) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_6_Q1), .B(SubCellInst_SboxInst_6_Q6), .ZN(
        SubCellInst_SboxInst_6_L1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1816), 
        .B(new_AGEMA_signal_1820), .Z(new_AGEMA_signal_1972) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1817), 
        .B(new_AGEMA_signal_1821), .Z(new_AGEMA_signal_1973) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_n3), .Z(SubCellInst_SboxInst_6_L2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        Ciphertext_s1[26]), .Z(new_AGEMA_signal_1822) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        Ciphertext_s2[26]), .Z(new_AGEMA_signal_1823) );
  INV_X1 SubCellInst_SboxInst_7_U1_U1 ( .A(Ciphertext_s0[30]), .ZN(
        SubCellInst_SboxInst_7_n3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[30]), 
        .B(Ciphertext_s0[31]), .Z(SubCellInst_SboxInst_7_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[30]), 
        .B(Ciphertext_s1[31]), .Z(new_AGEMA_signal_1254) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[30]), 
        .B(Ciphertext_s2[31]), .Z(new_AGEMA_signal_1255) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[28]), 
        .B(Ciphertext_s0[30]), .Z(SubCellInst_SboxInst_7_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[28]), 
        .B(Ciphertext_s1[30]), .Z(new_AGEMA_signal_1258) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[28]), 
        .B(Ciphertext_s2[30]), .Z(new_AGEMA_signal_1259) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_XX_2_), .Z(SubCellInst_SboxInst_7_Q0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        new_AGEMA_signal_1258), .Z(new_AGEMA_signal_1826) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        new_AGEMA_signal_1259), .Z(new_AGEMA_signal_1827) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_XX_1_), .Z(SubCellInst_SboxInst_7_Q1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        new_AGEMA_signal_1254), .Z(new_AGEMA_signal_1828) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        new_AGEMA_signal_1255), .Z(new_AGEMA_signal_1829) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_n3), .ZN(SubCellInst_SboxInst_7_Q4) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        Ciphertext_s1[30]), .Z(new_AGEMA_signal_1830) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        Ciphertext_s2[30]), .Z(new_AGEMA_signal_1831) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_XX_2_), .B(SubCellInst_SboxInst_7_n3), .Z(
        SubCellInst_SboxInst_7_Q6) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1258), 
        .B(Ciphertext_s1[30]), .Z(new_AGEMA_signal_1832) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1259), 
        .B(Ciphertext_s2[30]), .Z(new_AGEMA_signal_1833) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_7_Q1), .B(SubCellInst_SboxInst_7_Q6), .ZN(
        SubCellInst_SboxInst_7_L1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1828), 
        .B(new_AGEMA_signal_1832), .Z(new_AGEMA_signal_1978) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1829), 
        .B(new_AGEMA_signal_1833), .Z(new_AGEMA_signal_1979) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_n3), .Z(SubCellInst_SboxInst_7_L2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        Ciphertext_s1[30]), .Z(new_AGEMA_signal_1834) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        Ciphertext_s2[30]), .Z(new_AGEMA_signal_1835) );
  INV_X1 SubCellInst_SboxInst_8_U1_U1 ( .A(Ciphertext_s0[34]), .ZN(
        SubCellInst_SboxInst_8_n3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[34]), 
        .B(Ciphertext_s0[35]), .Z(SubCellInst_SboxInst_8_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[34]), 
        .B(Ciphertext_s1[35]), .Z(new_AGEMA_signal_1266) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[34]), 
        .B(Ciphertext_s2[35]), .Z(new_AGEMA_signal_1267) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[32]), 
        .B(Ciphertext_s0[34]), .Z(SubCellInst_SboxInst_8_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[32]), 
        .B(Ciphertext_s1[34]), .Z(new_AGEMA_signal_1270) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[32]), 
        .B(Ciphertext_s2[34]), .Z(new_AGEMA_signal_1271) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_XX_2_), .Z(SubCellInst_SboxInst_8_Q0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        new_AGEMA_signal_1270), .Z(new_AGEMA_signal_1838) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        new_AGEMA_signal_1271), .Z(new_AGEMA_signal_1839) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_XX_1_), .Z(SubCellInst_SboxInst_8_Q1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        new_AGEMA_signal_1266), .Z(new_AGEMA_signal_1840) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        new_AGEMA_signal_1267), .Z(new_AGEMA_signal_1841) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_n3), .ZN(SubCellInst_SboxInst_8_Q4) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        Ciphertext_s1[34]), .Z(new_AGEMA_signal_1842) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        Ciphertext_s2[34]), .Z(new_AGEMA_signal_1843) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_XX_2_), .B(SubCellInst_SboxInst_8_n3), .Z(
        SubCellInst_SboxInst_8_Q6) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1270), 
        .B(Ciphertext_s1[34]), .Z(new_AGEMA_signal_1844) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1271), 
        .B(Ciphertext_s2[34]), .Z(new_AGEMA_signal_1845) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_8_Q1), .B(SubCellInst_SboxInst_8_Q6), .ZN(
        SubCellInst_SboxInst_8_L1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1840), 
        .B(new_AGEMA_signal_1844), .Z(new_AGEMA_signal_1984) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1841), 
        .B(new_AGEMA_signal_1845), .Z(new_AGEMA_signal_1985) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_n3), .Z(SubCellInst_SboxInst_8_L2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        Ciphertext_s1[34]), .Z(new_AGEMA_signal_1846) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        Ciphertext_s2[34]), .Z(new_AGEMA_signal_1847) );
  INV_X1 SubCellInst_SboxInst_9_U1_U1 ( .A(Ciphertext_s0[38]), .ZN(
        SubCellInst_SboxInst_9_n3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[38]), 
        .B(Ciphertext_s0[39]), .Z(SubCellInst_SboxInst_9_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[38]), 
        .B(Ciphertext_s1[39]), .Z(new_AGEMA_signal_1278) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[38]), 
        .B(Ciphertext_s2[39]), .Z(new_AGEMA_signal_1279) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[36]), 
        .B(Ciphertext_s0[38]), .Z(SubCellInst_SboxInst_9_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[36]), 
        .B(Ciphertext_s1[38]), .Z(new_AGEMA_signal_1282) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[36]), 
        .B(Ciphertext_s2[38]), .Z(new_AGEMA_signal_1283) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_XX_2_), .Z(SubCellInst_SboxInst_9_Q0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        new_AGEMA_signal_1282), .Z(new_AGEMA_signal_1850) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        new_AGEMA_signal_1283), .Z(new_AGEMA_signal_1851) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_XX_1_), .Z(SubCellInst_SboxInst_9_Q1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        new_AGEMA_signal_1278), .Z(new_AGEMA_signal_1852) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        new_AGEMA_signal_1279), .Z(new_AGEMA_signal_1853) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_n3), .ZN(SubCellInst_SboxInst_9_Q4) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        Ciphertext_s1[38]), .Z(new_AGEMA_signal_1854) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        Ciphertext_s2[38]), .Z(new_AGEMA_signal_1855) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_XX_2_), .B(SubCellInst_SboxInst_9_n3), .Z(
        SubCellInst_SboxInst_9_Q6) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1282), 
        .B(Ciphertext_s1[38]), .Z(new_AGEMA_signal_1856) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1283), 
        .B(Ciphertext_s2[38]), .Z(new_AGEMA_signal_1857) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_9_Q1), .B(SubCellInst_SboxInst_9_Q6), .ZN(
        SubCellInst_SboxInst_9_L1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1852), 
        .B(new_AGEMA_signal_1856), .Z(new_AGEMA_signal_1990) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1853), 
        .B(new_AGEMA_signal_1857), .Z(new_AGEMA_signal_1991) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_n3), .Z(SubCellInst_SboxInst_9_L2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        Ciphertext_s1[38]), .Z(new_AGEMA_signal_1858) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        Ciphertext_s2[38]), .Z(new_AGEMA_signal_1859) );
  INV_X1 SubCellInst_SboxInst_10_U1_U1 ( .A(Ciphertext_s0[42]), .ZN(
        SubCellInst_SboxInst_10_n3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[42]), 
        .B(Ciphertext_s0[43]), .Z(SubCellInst_SboxInst_10_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[42]), 
        .B(Ciphertext_s1[43]), .Z(new_AGEMA_signal_1290) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[42]), 
        .B(Ciphertext_s2[43]), .Z(new_AGEMA_signal_1291) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[40]), 
        .B(Ciphertext_s0[42]), .Z(SubCellInst_SboxInst_10_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[40]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1294) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[40]), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_1295) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_XX_2_), .Z(SubCellInst_SboxInst_10_Q0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(new_AGEMA_signal_1294), .Z(new_AGEMA_signal_1862) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(new_AGEMA_signal_1295), .Z(new_AGEMA_signal_1863) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_XX_1_), .Z(SubCellInst_SboxInst_10_Q1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(new_AGEMA_signal_1290), .Z(new_AGEMA_signal_1864) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(new_AGEMA_signal_1291), .Z(new_AGEMA_signal_1865) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_Q4) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1866) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_1867) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_XX_2_), .B(SubCellInst_SboxInst_10_n3), .Z(
        SubCellInst_SboxInst_10_Q6) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1294), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1868) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1295), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_1869) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_10_Q1), .B(SubCellInst_SboxInst_10_Q6), .ZN(
        SubCellInst_SboxInst_10_L1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1864), 
        .B(new_AGEMA_signal_1868), .Z(new_AGEMA_signal_1996) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1865), 
        .B(new_AGEMA_signal_1869), .Z(new_AGEMA_signal_1997) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_n3), .Z(SubCellInst_SboxInst_10_L2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1870) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_1871) );
  INV_X1 SubCellInst_SboxInst_11_U1_U1 ( .A(Ciphertext_s0[46]), .ZN(
        SubCellInst_SboxInst_11_n3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[46]), 
        .B(Ciphertext_s0[47]), .Z(SubCellInst_SboxInst_11_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[46]), 
        .B(Ciphertext_s1[47]), .Z(new_AGEMA_signal_1302) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[46]), 
        .B(Ciphertext_s2[47]), .Z(new_AGEMA_signal_1303) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[44]), 
        .B(Ciphertext_s0[46]), .Z(SubCellInst_SboxInst_11_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[44]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1306) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[44]), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_1307) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_XX_2_), .Z(SubCellInst_SboxInst_11_Q0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(new_AGEMA_signal_1306), .Z(new_AGEMA_signal_1874) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(new_AGEMA_signal_1307), .Z(new_AGEMA_signal_1875) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_XX_1_), .Z(SubCellInst_SboxInst_11_Q1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(new_AGEMA_signal_1302), .Z(new_AGEMA_signal_1876) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(new_AGEMA_signal_1303), .Z(new_AGEMA_signal_1877) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_Q4) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1878) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_1879) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_XX_2_), .B(SubCellInst_SboxInst_11_n3), .Z(
        SubCellInst_SboxInst_11_Q6) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1306), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1880) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1307), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_1881) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_11_Q1), .B(SubCellInst_SboxInst_11_Q6), .ZN(
        SubCellInst_SboxInst_11_L1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1876), 
        .B(new_AGEMA_signal_1880), .Z(new_AGEMA_signal_2002) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1877), 
        .B(new_AGEMA_signal_1881), .Z(new_AGEMA_signal_2003) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_n3), .Z(SubCellInst_SboxInst_11_L2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1882) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_1883) );
  INV_X1 SubCellInst_SboxInst_12_U1_U1 ( .A(Ciphertext_s0[50]), .ZN(
        SubCellInst_SboxInst_12_n3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[50]), 
        .B(Ciphertext_s0[51]), .Z(SubCellInst_SboxInst_12_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[50]), 
        .B(Ciphertext_s1[51]), .Z(new_AGEMA_signal_1314) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[50]), 
        .B(Ciphertext_s2[51]), .Z(new_AGEMA_signal_1315) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[48]), 
        .B(Ciphertext_s0[50]), .Z(SubCellInst_SboxInst_12_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[48]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1318) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[48]), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_1319) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_XX_2_), .Z(SubCellInst_SboxInst_12_Q0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(new_AGEMA_signal_1318), .Z(new_AGEMA_signal_1886) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(new_AGEMA_signal_1319), .Z(new_AGEMA_signal_1887) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_XX_1_), .Z(SubCellInst_SboxInst_12_Q1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(new_AGEMA_signal_1314), .Z(new_AGEMA_signal_1888) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(new_AGEMA_signal_1315), .Z(new_AGEMA_signal_1889) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_Q4) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1890) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_1891) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_XX_2_), .B(SubCellInst_SboxInst_12_n3), .Z(
        SubCellInst_SboxInst_12_Q6) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1318), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1892) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1319), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_1893) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_12_Q1), .B(SubCellInst_SboxInst_12_Q6), .ZN(
        SubCellInst_SboxInst_12_L1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1888), 
        .B(new_AGEMA_signal_1892), .Z(new_AGEMA_signal_2008) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1889), 
        .B(new_AGEMA_signal_1893), .Z(new_AGEMA_signal_2009) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_n3), .Z(SubCellInst_SboxInst_12_L2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1894) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_1895) );
  INV_X1 SubCellInst_SboxInst_13_U1_U1 ( .A(Ciphertext_s0[54]), .ZN(
        SubCellInst_SboxInst_13_n3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[54]), 
        .B(Ciphertext_s0[55]), .Z(SubCellInst_SboxInst_13_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[54]), 
        .B(Ciphertext_s1[55]), .Z(new_AGEMA_signal_1326) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[54]), 
        .B(Ciphertext_s2[55]), .Z(new_AGEMA_signal_1327) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[52]), 
        .B(Ciphertext_s0[54]), .Z(SubCellInst_SboxInst_13_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[52]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1330) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[52]), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_1331) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_XX_2_), .Z(SubCellInst_SboxInst_13_Q0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(new_AGEMA_signal_1330), .Z(new_AGEMA_signal_1898) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(new_AGEMA_signal_1331), .Z(new_AGEMA_signal_1899) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_XX_1_), .Z(SubCellInst_SboxInst_13_Q1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(new_AGEMA_signal_1326), .Z(new_AGEMA_signal_1900) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(new_AGEMA_signal_1327), .Z(new_AGEMA_signal_1901) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_Q4) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1902) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_1903) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_XX_2_), .B(SubCellInst_SboxInst_13_n3), .Z(
        SubCellInst_SboxInst_13_Q6) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1330), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1904) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1331), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_1905) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_13_Q1), .B(SubCellInst_SboxInst_13_Q6), .ZN(
        SubCellInst_SboxInst_13_L1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1900), 
        .B(new_AGEMA_signal_1904), .Z(new_AGEMA_signal_2014) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1901), 
        .B(new_AGEMA_signal_1905), .Z(new_AGEMA_signal_2015) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_n3), .Z(SubCellInst_SboxInst_13_L2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1906) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_1907) );
  INV_X1 SubCellInst_SboxInst_14_U1_U1 ( .A(Ciphertext_s0[58]), .ZN(
        SubCellInst_SboxInst_14_n3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[58]), 
        .B(Ciphertext_s0[59]), .Z(SubCellInst_SboxInst_14_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[58]), 
        .B(Ciphertext_s1[59]), .Z(new_AGEMA_signal_1338) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[58]), 
        .B(Ciphertext_s2[59]), .Z(new_AGEMA_signal_1339) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[56]), 
        .B(Ciphertext_s0[58]), .Z(SubCellInst_SboxInst_14_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[56]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1342) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[56]), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_1343) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_XX_2_), .Z(SubCellInst_SboxInst_14_Q0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(new_AGEMA_signal_1342), .Z(new_AGEMA_signal_1910) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(new_AGEMA_signal_1343), .Z(new_AGEMA_signal_1911) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_XX_1_), .Z(SubCellInst_SboxInst_14_Q1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(new_AGEMA_signal_1338), .Z(new_AGEMA_signal_1912) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(new_AGEMA_signal_1339), .Z(new_AGEMA_signal_1913) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_Q4) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1914) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_1915) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_XX_2_), .B(SubCellInst_SboxInst_14_n3), .Z(
        SubCellInst_SboxInst_14_Q6) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1342), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1916) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1343), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_1917) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_14_Q1), .B(SubCellInst_SboxInst_14_Q6), .ZN(
        SubCellInst_SboxInst_14_L1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1912), 
        .B(new_AGEMA_signal_1916), .Z(new_AGEMA_signal_2020) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1913), 
        .B(new_AGEMA_signal_1917), .Z(new_AGEMA_signal_2021) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_n3), .Z(SubCellInst_SboxInst_14_L2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1918) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_1919) );
  INV_X1 SubCellInst_SboxInst_15_U1_U1 ( .A(Ciphertext_s0[62]), .ZN(
        SubCellInst_SboxInst_15_n3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[62]), 
        .B(Ciphertext_s0[63]), .Z(SubCellInst_SboxInst_15_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[62]), 
        .B(Ciphertext_s1[63]), .Z(new_AGEMA_signal_1350) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[62]), 
        .B(Ciphertext_s2[63]), .Z(new_AGEMA_signal_1351) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[60]), 
        .B(Ciphertext_s0[62]), .Z(SubCellInst_SboxInst_15_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[60]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1354) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[60]), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_1355) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_XX_2_), .Z(SubCellInst_SboxInst_15_Q0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(new_AGEMA_signal_1354), .Z(new_AGEMA_signal_1922) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(new_AGEMA_signal_1355), .Z(new_AGEMA_signal_1923) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_XX_1_), .Z(SubCellInst_SboxInst_15_Q1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(new_AGEMA_signal_1350), .Z(new_AGEMA_signal_1924) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(new_AGEMA_signal_1351), .Z(new_AGEMA_signal_1925) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_Q4) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1926) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_1927) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_XX_2_), .B(SubCellInst_SboxInst_15_n3), .Z(
        SubCellInst_SboxInst_15_Q6) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1354), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1928) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1355), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_1929) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_15_Q1), .B(SubCellInst_SboxInst_15_Q6), .ZN(
        SubCellInst_SboxInst_15_L1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1924), 
        .B(new_AGEMA_signal_1928), .Z(new_AGEMA_signal_2026) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1925), 
        .B(new_AGEMA_signal_1929), .Z(new_AGEMA_signal_2027) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_n3), .Z(SubCellInst_SboxInst_15_L2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1930) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_1931) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[0]), .B(Key_s0[0]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[0]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1356), .B(Key_s1[0]), .S(rst), .Z(
        new_AGEMA_signal_1360) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1357), .B(Key_s2[0]), .S(rst), .Z(
        new_AGEMA_signal_1361) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[1]), .B(Key_s0[1]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[1]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1362), .B(Key_s1[1]), .S(rst), .Z(
        new_AGEMA_signal_1366) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1363), .B(Key_s2[1]), .S(rst), .Z(
        new_AGEMA_signal_1367) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[2]), .B(Key_s0[2]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[2]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1368), .B(Key_s1[2]), .S(rst), .Z(
        new_AGEMA_signal_1372) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1369), .B(Key_s2[2]), .S(rst), .Z(
        new_AGEMA_signal_1373) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[3]), .B(Key_s0[3]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[3]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1374), .B(Key_s1[3]), .S(rst), .Z(
        new_AGEMA_signal_1378) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1375), .B(Key_s2[3]), .S(rst), .Z(
        new_AGEMA_signal_1379) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[4]), .B(Key_s0[4]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[4]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1380), .B(Key_s1[4]), .S(rst), .Z(
        new_AGEMA_signal_1384) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1381), .B(Key_s2[4]), .S(rst), .Z(
        new_AGEMA_signal_1385) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[5]), .B(Key_s0[5]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[5]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1386), .B(Key_s1[5]), .S(rst), .Z(
        new_AGEMA_signal_1390) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1387), .B(Key_s2[5]), .S(rst), .Z(
        new_AGEMA_signal_1391) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[6]), .B(Key_s0[6]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[6]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1392), .B(Key_s1[6]), .S(rst), .Z(
        new_AGEMA_signal_1396) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1393), .B(Key_s2[6]), .S(rst), .Z(
        new_AGEMA_signal_1397) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[7]), .B(Key_s0[7]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[7]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1398), .B(Key_s1[7]), .S(rst), .Z(
        new_AGEMA_signal_1402) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1399), .B(Key_s2[7]), .S(rst), .Z(
        new_AGEMA_signal_1403) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[8]), .B(Key_s0[8]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[8]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1404), .B(Key_s1[8]), .S(rst), .Z(
        new_AGEMA_signal_1408) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1405), .B(Key_s2[8]), .S(rst), .Z(
        new_AGEMA_signal_1409) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[9]), .B(Key_s0[9]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[9]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1410), .B(Key_s1[9]), .S(rst), .Z(
        new_AGEMA_signal_1414) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1411), .B(Key_s2[9]), .S(rst), .Z(
        new_AGEMA_signal_1415) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[10]), .B(Key_s0[10]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[10]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1416), .B(Key_s1[10]), .S(rst), .Z(
        new_AGEMA_signal_1420) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1417), .B(Key_s2[10]), .S(rst), .Z(
        new_AGEMA_signal_1421) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[11]), .B(Key_s0[11]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[11]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1422), .B(Key_s1[11]), .S(rst), .Z(
        new_AGEMA_signal_1426) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1423), .B(Key_s2[11]), .S(rst), .Z(
        new_AGEMA_signal_1427) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[12]), .B(Key_s0[12]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[12]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1428), .B(Key_s1[12]), .S(rst), .Z(
        new_AGEMA_signal_1432) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1429), .B(Key_s2[12]), .S(rst), .Z(
        new_AGEMA_signal_1433) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[13]), .B(Key_s0[13]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[13]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1434), .B(Key_s1[13]), .S(rst), .Z(
        new_AGEMA_signal_1438) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1435), .B(Key_s2[13]), .S(rst), .Z(
        new_AGEMA_signal_1439) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[14]), .B(Key_s0[14]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[14]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1440), .B(Key_s1[14]), .S(rst), .Z(
        new_AGEMA_signal_1444) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1441), .B(Key_s2[14]), .S(rst), .Z(
        new_AGEMA_signal_1445) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[15]), .B(Key_s0[15]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[15]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1446), .B(Key_s1[15]), .S(rst), .Z(
        new_AGEMA_signal_1450) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1447), .B(Key_s2[15]), .S(rst), .Z(
        new_AGEMA_signal_1451) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[16]), .B(Key_s0[16]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[16]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1452), .B(Key_s1[16]), .S(rst), .Z(
        new_AGEMA_signal_1456) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1453), .B(Key_s2[16]), .S(rst), .Z(
        new_AGEMA_signal_1457) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[17]), .B(Key_s0[17]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[17]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1458), .B(Key_s1[17]), .S(rst), .Z(
        new_AGEMA_signal_1462) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1459), .B(Key_s2[17]), .S(rst), .Z(
        new_AGEMA_signal_1463) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[18]), .B(Key_s0[18]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[18]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1464), .B(Key_s1[18]), .S(rst), .Z(
        new_AGEMA_signal_1468) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1465), .B(Key_s2[18]), .S(rst), .Z(
        new_AGEMA_signal_1469) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[19]), .B(Key_s0[19]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[19]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1470), .B(Key_s1[19]), .S(rst), .Z(
        new_AGEMA_signal_1474) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1471), .B(Key_s2[19]), .S(rst), .Z(
        new_AGEMA_signal_1475) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[20]), .B(Key_s0[20]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[20]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1476), .B(Key_s1[20]), .S(rst), .Z(
        new_AGEMA_signal_1480) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1477), .B(Key_s2[20]), .S(rst), .Z(
        new_AGEMA_signal_1481) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[21]), .B(Key_s0[21]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[21]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1482), .B(Key_s1[21]), .S(rst), .Z(
        new_AGEMA_signal_1486) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1483), .B(Key_s2[21]), .S(rst), .Z(
        new_AGEMA_signal_1487) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[22]), .B(Key_s0[22]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[22]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1488), .B(Key_s1[22]), .S(rst), .Z(
        new_AGEMA_signal_1492) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1489), .B(Key_s2[22]), .S(rst), .Z(
        new_AGEMA_signal_1493) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[23]), .B(Key_s0[23]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[23]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1494), .B(Key_s1[23]), .S(rst), .Z(
        new_AGEMA_signal_1498) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1495), .B(Key_s2[23]), .S(rst), .Z(
        new_AGEMA_signal_1499) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[24]), .B(Key_s0[24]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[24]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1500), .B(Key_s1[24]), .S(rst), .Z(
        new_AGEMA_signal_1504) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1501), .B(Key_s2[24]), .S(rst), .Z(
        new_AGEMA_signal_1505) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[25]), .B(Key_s0[25]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[25]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1506), .B(Key_s1[25]), .S(rst), .Z(
        new_AGEMA_signal_1510) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1507), .B(Key_s2[25]), .S(rst), .Z(
        new_AGEMA_signal_1511) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[26]), .B(Key_s0[26]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[26]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1512), .B(Key_s1[26]), .S(rst), .Z(
        new_AGEMA_signal_1516) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1513), .B(Key_s2[26]), .S(rst), .Z(
        new_AGEMA_signal_1517) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[27]), .B(Key_s0[27]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[27]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1518), .B(Key_s1[27]), .S(rst), .Z(
        new_AGEMA_signal_1522) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1519), .B(Key_s2[27]), .S(rst), .Z(
        new_AGEMA_signal_1523) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[28]), .B(Key_s0[28]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[28]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1524), .B(Key_s1[28]), .S(rst), .Z(
        new_AGEMA_signal_1528) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1525), .B(Key_s2[28]), .S(rst), .Z(
        new_AGEMA_signal_1529) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[29]), .B(Key_s0[29]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[29]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1530), .B(Key_s1[29]), .S(rst), .Z(
        new_AGEMA_signal_1534) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1531), .B(Key_s2[29]), .S(rst), .Z(
        new_AGEMA_signal_1535) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[30]), .B(Key_s0[30]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[30]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1536), .B(Key_s1[30]), .S(rst), .Z(
        new_AGEMA_signal_1540) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1537), .B(Key_s2[30]), .S(rst), .Z(
        new_AGEMA_signal_1541) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[31]), .B(Key_s0[31]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[31]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1542), .B(Key_s1[31]), .S(rst), .Z(
        new_AGEMA_signal_1546) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1543), .B(Key_s2[31]), .S(rst), .Z(
        new_AGEMA_signal_1547) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[32]), .B(Key_s0[32]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[32]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1548), .B(Key_s1[32]), .S(rst), .Z(
        new_AGEMA_signal_1552) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1549), .B(Key_s2[32]), .S(rst), .Z(
        new_AGEMA_signal_1553) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[33]), .B(Key_s0[33]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[33]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1554), .B(Key_s1[33]), .S(rst), .Z(
        new_AGEMA_signal_1558) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1555), .B(Key_s2[33]), .S(rst), .Z(
        new_AGEMA_signal_1559) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[34]), .B(Key_s0[34]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[34]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1560), .B(Key_s1[34]), .S(rst), .Z(
        new_AGEMA_signal_1564) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1561), .B(Key_s2[34]), .S(rst), .Z(
        new_AGEMA_signal_1565) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[35]), .B(Key_s0[35]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[35]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1566), .B(Key_s1[35]), .S(rst), .Z(
        new_AGEMA_signal_1570) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1567), .B(Key_s2[35]), .S(rst), .Z(
        new_AGEMA_signal_1571) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[36]), .B(Key_s0[36]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[36]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1572), .B(Key_s1[36]), .S(rst), .Z(
        new_AGEMA_signal_1576) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1573), .B(Key_s2[36]), .S(rst), .Z(
        new_AGEMA_signal_1577) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[37]), .B(Key_s0[37]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[37]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1578), .B(Key_s1[37]), .S(rst), .Z(
        new_AGEMA_signal_1582) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1579), .B(Key_s2[37]), .S(rst), .Z(
        new_AGEMA_signal_1583) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[38]), .B(Key_s0[38]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[38]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1584), .B(Key_s1[38]), .S(rst), .Z(
        new_AGEMA_signal_1588) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1585), .B(Key_s2[38]), .S(rst), .Z(
        new_AGEMA_signal_1589) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[39]), .B(Key_s0[39]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[39]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1590), .B(Key_s1[39]), .S(rst), .Z(
        new_AGEMA_signal_1594) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1591), .B(Key_s2[39]), .S(rst), .Z(
        new_AGEMA_signal_1595) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[40]), .B(Key_s0[40]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[40]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1596), .B(Key_s1[40]), .S(rst), .Z(
        new_AGEMA_signal_1600) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1597), .B(Key_s2[40]), .S(rst), .Z(
        new_AGEMA_signal_1601) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[41]), .B(Key_s0[41]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[41]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1602), .B(Key_s1[41]), .S(rst), .Z(
        new_AGEMA_signal_1606) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1603), .B(Key_s2[41]), .S(rst), .Z(
        new_AGEMA_signal_1607) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[42]), .B(Key_s0[42]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[42]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1608), .B(Key_s1[42]), .S(rst), .Z(
        new_AGEMA_signal_1612) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1609), .B(Key_s2[42]), .S(rst), .Z(
        new_AGEMA_signal_1613) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[43]), .B(Key_s0[43]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[43]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1614), .B(Key_s1[43]), .S(rst), .Z(
        new_AGEMA_signal_1618) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1615), .B(Key_s2[43]), .S(rst), .Z(
        new_AGEMA_signal_1619) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[44]), .B(Key_s0[44]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[44]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1620), .B(Key_s1[44]), .S(rst), .Z(
        new_AGEMA_signal_1624) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1621), .B(Key_s2[44]), .S(rst), .Z(
        new_AGEMA_signal_1625) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[45]), .B(Key_s0[45]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[45]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1626), .B(Key_s1[45]), .S(rst), .Z(
        new_AGEMA_signal_1630) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1627), .B(Key_s2[45]), .S(rst), .Z(
        new_AGEMA_signal_1631) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[46]), .B(Key_s0[46]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[46]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1632), .B(Key_s1[46]), .S(rst), .Z(
        new_AGEMA_signal_1636) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1633), .B(Key_s2[46]), .S(rst), .Z(
        new_AGEMA_signal_1637) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[47]), .B(Key_s0[47]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[47]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1638), .B(Key_s1[47]), .S(rst), .Z(
        new_AGEMA_signal_1642) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1639), .B(Key_s2[47]), .S(rst), .Z(
        new_AGEMA_signal_1643) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[48]), .B(Key_s0[48]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[48]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1644), .B(Key_s1[48]), .S(rst), .Z(
        new_AGEMA_signal_1648) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1645), .B(Key_s2[48]), .S(rst), .Z(
        new_AGEMA_signal_1649) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[49]), .B(Key_s0[49]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[49]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1650), .B(Key_s1[49]), .S(rst), .Z(
        new_AGEMA_signal_1654) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1651), .B(Key_s2[49]), .S(rst), .Z(
        new_AGEMA_signal_1655) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[50]), .B(Key_s0[50]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[50]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1656), .B(Key_s1[50]), .S(rst), .Z(
        new_AGEMA_signal_1660) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1657), .B(Key_s2[50]), .S(rst), .Z(
        new_AGEMA_signal_1661) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[51]), .B(Key_s0[51]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[51]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1662), .B(Key_s1[51]), .S(rst), .Z(
        new_AGEMA_signal_1666) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1663), .B(Key_s2[51]), .S(rst), .Z(
        new_AGEMA_signal_1667) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[52]), .B(Key_s0[52]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[52]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1668), .B(Key_s1[52]), .S(rst), .Z(
        new_AGEMA_signal_1672) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1669), .B(Key_s2[52]), .S(rst), .Z(
        new_AGEMA_signal_1673) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[53]), .B(Key_s0[53]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[53]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1674), .B(Key_s1[53]), .S(rst), .Z(
        new_AGEMA_signal_1678) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1675), .B(Key_s2[53]), .S(rst), .Z(
        new_AGEMA_signal_1679) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[54]), .B(Key_s0[54]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[54]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1680), .B(Key_s1[54]), .S(rst), .Z(
        new_AGEMA_signal_1684) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1681), .B(Key_s2[54]), .S(rst), .Z(
        new_AGEMA_signal_1685) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[55]), .B(Key_s0[55]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[55]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1686), .B(Key_s1[55]), .S(rst), .Z(
        new_AGEMA_signal_1690) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1687), .B(Key_s2[55]), .S(rst), .Z(
        new_AGEMA_signal_1691) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[56]), .B(Key_s0[56]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[56]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1692), .B(Key_s1[56]), .S(rst), .Z(
        new_AGEMA_signal_1696) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1693), .B(Key_s2[56]), .S(rst), .Z(
        new_AGEMA_signal_1697) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[57]), .B(Key_s0[57]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[57]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1698), .B(Key_s1[57]), .S(rst), .Z(
        new_AGEMA_signal_1702) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1699), .B(Key_s2[57]), .S(rst), .Z(
        new_AGEMA_signal_1703) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[58]), .B(Key_s0[58]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[58]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1704), .B(Key_s1[58]), .S(rst), .Z(
        new_AGEMA_signal_1708) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1705), .B(Key_s2[58]), .S(rst), .Z(
        new_AGEMA_signal_1709) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[59]), .B(Key_s0[59]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[59]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1710), .B(Key_s1[59]), .S(rst), .Z(
        new_AGEMA_signal_1714) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1711), .B(Key_s2[59]), .S(rst), .Z(
        new_AGEMA_signal_1715) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[60]), .B(Key_s0[60]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[60]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1716), .B(Key_s1[60]), .S(rst), .Z(
        new_AGEMA_signal_1720) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1717), .B(Key_s2[60]), .S(rst), .Z(
        new_AGEMA_signal_1721) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[61]), .B(Key_s0[61]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[61]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1722), .B(Key_s1[61]), .S(rst), .Z(
        new_AGEMA_signal_1726) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1723), .B(Key_s2[61]), .S(rst), .Z(
        new_AGEMA_signal_1727) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[62]), .B(Key_s0[62]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[62]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1728), .B(Key_s1[62]), .S(rst), .Z(
        new_AGEMA_signal_1732) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1729), .B(Key_s2[62]), .S(rst), .Z(
        new_AGEMA_signal_1733) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[63]), .B(Key_s0[63]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[63]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1734), .B(Key_s1[63]), .S(rst), .Z(
        new_AGEMA_signal_1738) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1735), .B(Key_s2[63]), .S(rst), .Z(
        new_AGEMA_signal_1739) );
  NOR2_X1 ClockGatingInst_U9 ( .A1(rst), .A2(ClockGatingInst_n9), .ZN(
        ClockGatingInst_n4) );
  NOR2_X1 ClockGatingInst_U8 ( .A1(rst), .A2(ClockGatingInst_n8), .ZN(
        ClockGatingInst_n3) );
  NOR2_X1 ClockGatingInst_U7 ( .A1(rst), .A2(ClockGatingInst_n7), .ZN(
        ClockGatingInst_n2) );
  NOR2_X1 ClockGatingInst_U6 ( .A1(rst), .A2(ClockGatingInst_n6), .ZN(
        ClockGatingInst_n1) );
  NAND2_X1 ClockGatingInst_U5 ( .A1(ClockGatingInst_n10), .A2(
        ClockGatingInst_n11), .ZN(ClockGatingInst_N7) );
  AND2_X1 ClockGatingInst_U4 ( .A1(ClockGatingInst_LatchedEnable), .A2(clk), 
        .ZN(clk_gated) );
  INV_X1 ClockGatingInst_U3 ( .A(rst), .ZN(ClockGatingInst_n11) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_2_ ( .D(ClockGatingInst_n1), .CK(
        clk), .Q(), .QN(ClockGatingInst_n7) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_3_ ( .D(ClockGatingInst_n2), .CK(
        clk), .Q(), .QN(ClockGatingInst_n8) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_4_ ( .D(ClockGatingInst_n3), .CK(
        clk), .Q(), .QN(ClockGatingInst_n9) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_5_ ( .D(ClockGatingInst_n4), .CK(
        clk), .Q(ClockGatingInst_ShiftRegister_5_), .QN(ClockGatingInst_n10)
         );
  DLL_X1 ClockGatingInst_LatchedEnable_reg ( .D(ClockGatingInst_N7), .GN(clk), 
        .Q(ClockGatingInst_LatchedEnable) );
  DLL_X1 ClockGatingInst_Synch_reg ( .D(ClockGatingInst_ShiftRegister_5_), 
        .GN(clk), .Q(Synch) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_1_ ( .D(ClockGatingInst_N7), .CK(
        clk), .Q(), .QN(ClockGatingInst_n6) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_0_U1 ( .A(MCOutput[2]), .B(
        Plaintext_s0[2]), .S(rst), .Z(StateRegInput[2]) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2666), .B(
        Plaintext_s1[2]), .S(rst), .Z(new_AGEMA_signal_2680) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2667), .B(
        Plaintext_s2[2]), .S(rst), .Z(new_AGEMA_signal_2681) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_0_U1 ( .A(MCOutput[3]), .B(
        Plaintext_s0[3]), .S(rst), .Z(StateRegInput[3]) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2786), .B(
        Plaintext_s1[3]), .S(rst), .Z(new_AGEMA_signal_2800) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2787), .B(
        Plaintext_s2[3]), .S(rst), .Z(new_AGEMA_signal_2801) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_0_U1 ( .A(MCOutput[6]), .B(
        Plaintext_s0[6]), .S(rst), .Z(StateRegInput[6]) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2670), .B(
        Plaintext_s1[6]), .S(rst), .Z(new_AGEMA_signal_2684) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2671), .B(
        Plaintext_s2[6]), .S(rst), .Z(new_AGEMA_signal_2685) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_0_U1 ( .A(MCOutput[7]), .B(
        Plaintext_s0[7]), .S(rst), .Z(StateRegInput[7]) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2790), .B(
        Plaintext_s1[7]), .S(rst), .Z(new_AGEMA_signal_2804) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2791), .B(
        Plaintext_s2[7]), .S(rst), .Z(new_AGEMA_signal_2805) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_0_U1 ( .A(MCOutput[10]), .B(
        Plaintext_s0[10]), .S(rst), .Z(StateRegInput[10]) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2674), .B(
        Plaintext_s1[10]), .S(rst), .Z(new_AGEMA_signal_2688) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2675), .B(
        Plaintext_s2[10]), .S(rst), .Z(new_AGEMA_signal_2689) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_0_U1 ( .A(MCOutput[11]), .B(
        Plaintext_s0[11]), .S(rst), .Z(StateRegInput[11]) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2794), .B(
        Plaintext_s1[11]), .S(rst), .Z(new_AGEMA_signal_2808) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2795), .B(
        Plaintext_s2[11]), .S(rst), .Z(new_AGEMA_signal_2809) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_0_U1 ( .A(MCOutput[14]), .B(
        Plaintext_s0[14]), .S(rst), .Z(StateRegInput[14]) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2902), .B(
        Plaintext_s1[14]), .S(rst), .Z(new_AGEMA_signal_2920) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2903), .B(
        Plaintext_s2[14]), .S(rst), .Z(new_AGEMA_signal_2921) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_0_U1 ( .A(MCOutput[15]), .B(
        Plaintext_s0[15]), .S(rst), .Z(StateRegInput[15]) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2990), .B(
        Plaintext_s1[15]), .S(rst), .Z(new_AGEMA_signal_3006) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2991), .B(
        Plaintext_s2[15]), .S(rst), .Z(new_AGEMA_signal_3007) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_0_U1 ( .A(MCOutput[18]), .B(
        Plaintext_s0[18]), .S(rst), .Z(StateRegInput[18]) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2654), .B(
        Plaintext_s1[18]), .S(rst), .Z(new_AGEMA_signal_2692) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2655), .B(
        Plaintext_s2[18]), .S(rst), .Z(new_AGEMA_signal_2693) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_0_U1 ( .A(MCOutput[19]), .B(
        Plaintext_s0[19]), .S(rst), .Z(StateRegInput[19]) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2772), .B(
        Plaintext_s1[19]), .S(rst), .Z(new_AGEMA_signal_2812) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2773), .B(
        Plaintext_s2[19]), .S(rst), .Z(new_AGEMA_signal_2813) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_0_U1 ( .A(MCOutput[22]), .B(
        Plaintext_s0[22]), .S(rst), .Z(StateRegInput[22]) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2658), .B(
        Plaintext_s1[22]), .S(rst), .Z(new_AGEMA_signal_2696) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2659), .B(
        Plaintext_s2[22]), .S(rst), .Z(new_AGEMA_signal_2697) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_0_U1 ( .A(MCOutput[23]), .B(
        Plaintext_s0[23]), .S(rst), .Z(StateRegInput[23]) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2776), .B(
        Plaintext_s1[23]), .S(rst), .Z(new_AGEMA_signal_2816) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2777), .B(
        Plaintext_s2[23]), .S(rst), .Z(new_AGEMA_signal_2817) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_0_U1 ( .A(MCOutput[26]), .B(
        Plaintext_s0[26]), .S(rst), .Z(StateRegInput[26]) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2882), .B(
        Plaintext_s1[26]), .S(rst), .Z(new_AGEMA_signal_2932) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2883), .B(
        Plaintext_s2[26]), .S(rst), .Z(new_AGEMA_signal_2933) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_0_U1 ( .A(MCOutput[27]), .B(
        Plaintext_s0[27]), .S(rst), .Z(StateRegInput[27]) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2978), .B(
        Plaintext_s1[27]), .S(rst), .Z(new_AGEMA_signal_3018) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2979), .B(
        Plaintext_s2[27]), .S(rst), .Z(new_AGEMA_signal_3019) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_0_U1 ( .A(MCOutput[30]), .B(
        Plaintext_s0[30]), .S(rst), .Z(StateRegInput[30]) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2662), .B(
        Plaintext_s1[30]), .S(rst), .Z(new_AGEMA_signal_2700) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2663), .B(
        Plaintext_s2[30]), .S(rst), .Z(new_AGEMA_signal_2701) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_0_U1 ( .A(MCOutput[31]), .B(
        Plaintext_s0[31]), .S(rst), .Z(StateRegInput[31]) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2782), .B(
        Plaintext_s1[31]), .S(rst), .Z(new_AGEMA_signal_2820) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2783), .B(
        Plaintext_s2[31]), .S(rst), .Z(new_AGEMA_signal_2821) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_0_U1 ( .A(MCOutput[34]), .B(
        Plaintext_s0[34]), .S(rst), .Z(StateRegInput[34]) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2456), .B(
        Plaintext_s1[34]), .S(rst), .Z(new_AGEMA_signal_2478) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2457), .B(
        Plaintext_s2[34]), .S(rst), .Z(new_AGEMA_signal_2479) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_0_U1 ( .A(MCOutput[35]), .B(
        Plaintext_s0[35]), .S(rst), .Z(StateRegInput[35]) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2544), .B(
        Plaintext_s1[35]), .S(rst), .Z(new_AGEMA_signal_2584) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2545), .B(
        Plaintext_s2[35]), .S(rst), .Z(new_AGEMA_signal_2585) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_0_U1 ( .A(MCOutput[38]), .B(
        Plaintext_s0[38]), .S(rst), .Z(StateRegInput[38]) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2460), .B(
        Plaintext_s1[38]), .S(rst), .Z(new_AGEMA_signal_2482) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2461), .B(
        Plaintext_s2[38]), .S(rst), .Z(new_AGEMA_signal_2483) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_0_U1 ( .A(MCOutput[39]), .B(
        Plaintext_s0[39]), .S(rst), .Z(StateRegInput[39]) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2548), .B(
        Plaintext_s1[39]), .S(rst), .Z(new_AGEMA_signal_2588) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2549), .B(
        Plaintext_s2[39]), .S(rst), .Z(new_AGEMA_signal_2589) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_0_U1 ( .A(MCOutput[42]), .B(
        Plaintext_s0[42]), .S(rst), .Z(StateRegInput[42]) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2464), .B(
        Plaintext_s1[42]), .S(rst), .Z(new_AGEMA_signal_2486) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2465), .B(
        Plaintext_s2[42]), .S(rst), .Z(new_AGEMA_signal_2487) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_0_U1 ( .A(MCOutput[43]), .B(
        Plaintext_s0[43]), .S(rst), .Z(StateRegInput[43]) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2552), .B(
        Plaintext_s1[43]), .S(rst), .Z(new_AGEMA_signal_2592) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2553), .B(
        Plaintext_s2[43]), .S(rst), .Z(new_AGEMA_signal_2593) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_0_U1 ( .A(MCOutput[46]), .B(
        Plaintext_s0[46]), .S(rst), .Z(StateRegInput[46]) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2632), .B(
        Plaintext_s1[46]), .S(rst), .Z(new_AGEMA_signal_2716) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2633), .B(
        Plaintext_s2[46]), .S(rst), .Z(new_AGEMA_signal_2717) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_0_U1 ( .A(MCOutput[47]), .B(
        Plaintext_s0[47]), .S(rst), .Z(StateRegInput[47]) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2752), .B(
        Plaintext_s1[47]), .S(rst), .Z(new_AGEMA_signal_2836) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2753), .B(
        Plaintext_s2[47]), .S(rst), .Z(new_AGEMA_signal_2837) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_0_U1 ( .A(MCOutput[50]), .B(
        Plaintext_s0[50]), .S(rst), .Z(StateRegInput[50]) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2638), .B(
        Plaintext_s1[50]), .S(rst), .Z(new_AGEMA_signal_2720) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2639), .B(
        Plaintext_s2[50]), .S(rst), .Z(new_AGEMA_signal_2721) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_0_U1 ( .A(MCOutput[51]), .B(
        Plaintext_s0[51]), .S(rst), .Z(StateRegInput[51]) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2756), .B(
        Plaintext_s1[51]), .S(rst), .Z(new_AGEMA_signal_2840) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2757), .B(
        Plaintext_s2[51]), .S(rst), .Z(new_AGEMA_signal_2841) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_0_U1 ( .A(MCOutput[54]), .B(
        Plaintext_s0[54]), .S(rst), .Z(StateRegInput[54]) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2642), .B(
        Plaintext_s1[54]), .S(rst), .Z(new_AGEMA_signal_2724) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2643), .B(
        Plaintext_s2[54]), .S(rst), .Z(new_AGEMA_signal_2725) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_0_U1 ( .A(MCOutput[55]), .B(
        Plaintext_s0[55]), .S(rst), .Z(StateRegInput[55]) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2762), .B(
        Plaintext_s1[55]), .S(rst), .Z(new_AGEMA_signal_2844) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2763), .B(
        Plaintext_s2[55]), .S(rst), .Z(new_AGEMA_signal_2845) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_0_U1 ( .A(MCOutput[58]), .B(
        Plaintext_s0[58]), .S(rst), .Z(StateRegInput[58]) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2648), .B(
        Plaintext_s1[58]), .S(rst), .Z(new_AGEMA_signal_2728) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2649), .B(
        Plaintext_s2[58]), .S(rst), .Z(new_AGEMA_signal_2729) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_0_U1 ( .A(MCOutput[59]), .B(
        Plaintext_s0[59]), .S(rst), .Z(StateRegInput[59]) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2766), .B(
        Plaintext_s1[59]), .S(rst), .Z(new_AGEMA_signal_2848) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2767), .B(
        Plaintext_s2[59]), .S(rst), .Z(new_AGEMA_signal_2849) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_0_U1 ( .A(MCOutput[62]), .B(
        Plaintext_s0[62]), .S(rst), .Z(StateRegInput[62]) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2870), .B(
        Plaintext_s1[62]), .S(rst), .Z(new_AGEMA_signal_2956) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2871), .B(
        Plaintext_s2[62]), .S(rst), .Z(new_AGEMA_signal_2957) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_0_U1 ( .A(MCOutput[63]), .B(
        Plaintext_s0[63]), .S(rst), .Z(StateRegInput[63]) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2970), .B(
        Plaintext_s1[63]), .S(rst), .Z(new_AGEMA_signal_3042) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2971), .B(
        Plaintext_s2[63]), .S(rst), .Z(new_AGEMA_signal_3043) );
  INV_X1 SubCellInst_SboxInst_0_U3_U1 ( .A(SubCellInst_SboxInst_0_YY_1_), .ZN(
        ShiftRowsOutput[7]) );
  INV_X1 SubCellInst_SboxInst_0_U2_U1 ( .A(SubCellInst_SboxInst_0_YY_0_), .ZN(
        ShiftRowsOutput[6]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U37 ( .A(new_AGEMA_signal_1744), .B(
        Fresh[2]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U36 ( .A(Fresh[1]), .B(
        SubCellInst_SboxInst_0_Q1), .Z(
        SubCellInst_SboxInst_0_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U35 ( .A(new_AGEMA_signal_1745), .B(
        Fresh[2]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U34 ( .A(Fresh[0]), .B(
        SubCellInst_SboxInst_0_Q1), .Z(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U33 ( .A(Fresh[1]), .B(
        new_AGEMA_signal_1745), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U32 ( .A(new_AGEMA_signal_1744), .B(
        Fresh[0]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U25 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U24 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U23 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U22 ( .A(Fresh[2]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U21 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U19 ( .A(Fresh[1]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U17 ( .A(Fresh[0]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U16 ( .A1(new_AGEMA_signal_1745), 
        .A2(Ciphertext_s2[2]), .ZN(SubCellInst_SboxInst_0_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U15 ( .A1(new_AGEMA_signal_1744), 
        .A2(Ciphertext_s1[2]), .ZN(SubCellInst_SboxInst_0_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_0_Q1), 
        .A2(SubCellInst_SboxInst_0_n3), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_n33), .Z(new_AGEMA_signal_1933) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n32), .B(
        SubCellInst_SboxInst_0_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_n30), .Z(new_AGEMA_signal_1932) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n29), .B(
        SubCellInst_SboxInst_0_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_n27), .Z(SubCellInst_SboxInst_0_T0) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n26), .B(
        SubCellInst_SboxInst_0_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_Q0), .B(SubCellInst_SboxInst_0_T0), .Z(
        SubCellInst_SboxInst_0_Q2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1742), 
        .B(new_AGEMA_signal_1932), .Z(new_AGEMA_signal_2028) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1743), 
        .B(new_AGEMA_signal_1933), .Z(new_AGEMA_signal_2029) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U37 ( .A(new_AGEMA_signal_1746), .B(
        Fresh[5]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U36 ( .A(Fresh[4]), .B(
        SubCellInst_SboxInst_0_Q4), .Z(
        SubCellInst_SboxInst_0_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U35 ( .A(new_AGEMA_signal_1747), .B(
        Fresh[5]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U34 ( .A(Fresh[3]), .B(
        SubCellInst_SboxInst_0_Q4), .Z(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U33 ( .A(Fresh[4]), .B(
        new_AGEMA_signal_1747), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U32 ( .A(new_AGEMA_signal_1746), .B(
        Fresh[3]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U25 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U24 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U23 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U22 ( .A(Fresh[5]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U21 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U19 ( .A(Fresh[4]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U17 ( .A(Fresh[3]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U16 ( .A1(new_AGEMA_signal_1747), 
        .A2(Ciphertext_s2[2]), .ZN(SubCellInst_SboxInst_0_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U15 ( .A1(new_AGEMA_signal_1746), 
        .A2(Ciphertext_s1[2]), .ZN(SubCellInst_SboxInst_0_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_0_Q4), 
        .A2(SubCellInst_SboxInst_0_n3), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_n33), .Z(new_AGEMA_signal_1935) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n32), .B(
        SubCellInst_SboxInst_0_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_n30), .Z(new_AGEMA_signal_1934) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n29), .B(
        SubCellInst_SboxInst_0_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_n27), .Z(SubCellInst_SboxInst_0_T2) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n26), .B(
        SubCellInst_SboxInst_0_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L1), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_Q7) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1936), 
        .B(new_AGEMA_signal_1934), .Z(new_AGEMA_signal_2030) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1937), 
        .B(new_AGEMA_signal_1935), .Z(new_AGEMA_signal_2031) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_XX_2_), .B(SubCellInst_SboxInst_0_T0), .Z(
        SubCellInst_SboxInst_0_L3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1174), 
        .B(new_AGEMA_signal_1932), .Z(new_AGEMA_signal_2032) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1175), 
        .B(new_AGEMA_signal_1933), .Z(new_AGEMA_signal_2033) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L3), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2032), 
        .B(new_AGEMA_signal_1934), .Z(new_AGEMA_signal_2284) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2033), 
        .B(new_AGEMA_signal_1935), .Z(new_AGEMA_signal_2285) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_XX_1_), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1170), 
        .B(new_AGEMA_signal_1934), .Z(new_AGEMA_signal_2156) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1171), 
        .B(new_AGEMA_signal_1935), .Z(new_AGEMA_signal_2157) );
  INV_X1 SubCellInst_SboxInst_1_U3_U1 ( .A(SubCellInst_SboxInst_1_YY_1_), .ZN(
        ShiftRowsOutput[11]) );
  INV_X1 SubCellInst_SboxInst_1_U2_U1 ( .A(SubCellInst_SboxInst_1_YY_0_), .ZN(
        ShiftRowsOutput[10]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U37 ( .A(new_AGEMA_signal_1756), .B(
        Fresh[8]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U36 ( .A(Fresh[7]), .B(
        SubCellInst_SboxInst_1_Q1), .Z(
        SubCellInst_SboxInst_1_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U35 ( .A(new_AGEMA_signal_1757), .B(
        Fresh[8]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U34 ( .A(Fresh[6]), .B(
        SubCellInst_SboxInst_1_Q1), .Z(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U33 ( .A(Fresh[7]), .B(
        new_AGEMA_signal_1757), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U32 ( .A(new_AGEMA_signal_1756), .B(
        Fresh[6]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U25 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U24 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U23 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U22 ( .A(Fresh[8]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U21 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U19 ( .A(Fresh[7]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U17 ( .A(Fresh[6]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U16 ( .A1(new_AGEMA_signal_1757), 
        .A2(Ciphertext_s2[6]), .ZN(SubCellInst_SboxInst_1_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U15 ( .A1(new_AGEMA_signal_1756), 
        .A2(Ciphertext_s1[6]), .ZN(SubCellInst_SboxInst_1_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_1_Q1), 
        .A2(SubCellInst_SboxInst_1_n3), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_n33), .Z(new_AGEMA_signal_1939) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n32), .B(
        SubCellInst_SboxInst_1_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_n30), .Z(new_AGEMA_signal_1938) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n29), .B(
        SubCellInst_SboxInst_1_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_n27), .Z(SubCellInst_SboxInst_1_T0) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n26), .B(
        SubCellInst_SboxInst_1_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_Q0), .B(SubCellInst_SboxInst_1_T0), .Z(
        SubCellInst_SboxInst_1_Q2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1754), 
        .B(new_AGEMA_signal_1938), .Z(new_AGEMA_signal_2036) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1755), 
        .B(new_AGEMA_signal_1939), .Z(new_AGEMA_signal_2037) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U37 ( .A(new_AGEMA_signal_1758), .B(
        Fresh[11]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U36 ( .A(Fresh[10]), .B(
        SubCellInst_SboxInst_1_Q4), .Z(
        SubCellInst_SboxInst_1_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U35 ( .A(new_AGEMA_signal_1759), .B(
        Fresh[11]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U34 ( .A(Fresh[9]), .B(
        SubCellInst_SboxInst_1_Q4), .Z(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U33 ( .A(Fresh[10]), .B(
        new_AGEMA_signal_1759), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U32 ( .A(new_AGEMA_signal_1758), .B(
        Fresh[9]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U25 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U24 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U23 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U22 ( .A(Fresh[11]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U21 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U19 ( .A(Fresh[10]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U17 ( .A(Fresh[9]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U16 ( .A1(new_AGEMA_signal_1759), 
        .A2(Ciphertext_s2[6]), .ZN(SubCellInst_SboxInst_1_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U15 ( .A1(new_AGEMA_signal_1758), 
        .A2(Ciphertext_s1[6]), .ZN(SubCellInst_SboxInst_1_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_1_Q4), 
        .A2(SubCellInst_SboxInst_1_n3), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_n33), .Z(new_AGEMA_signal_1941) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n32), .B(
        SubCellInst_SboxInst_1_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_n30), .Z(new_AGEMA_signal_1940) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n29), .B(
        SubCellInst_SboxInst_1_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_n27), .Z(SubCellInst_SboxInst_1_T2) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n26), .B(
        SubCellInst_SboxInst_1_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L1), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_Q7) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1942), 
        .B(new_AGEMA_signal_1940), .Z(new_AGEMA_signal_2038) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1943), 
        .B(new_AGEMA_signal_1941), .Z(new_AGEMA_signal_2039) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_XX_2_), .B(SubCellInst_SboxInst_1_T0), .Z(
        SubCellInst_SboxInst_1_L3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1186), 
        .B(new_AGEMA_signal_1938), .Z(new_AGEMA_signal_2040) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1187), 
        .B(new_AGEMA_signal_1939), .Z(new_AGEMA_signal_2041) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L3), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2040), 
        .B(new_AGEMA_signal_1940), .Z(new_AGEMA_signal_2288) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2041), 
        .B(new_AGEMA_signal_1941), .Z(new_AGEMA_signal_2289) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_XX_1_), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1182), 
        .B(new_AGEMA_signal_1940), .Z(new_AGEMA_signal_2164) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1183), 
        .B(new_AGEMA_signal_1941), .Z(new_AGEMA_signal_2165) );
  INV_X1 SubCellInst_SboxInst_2_U3_U1 ( .A(SubCellInst_SboxInst_2_YY_1_), .ZN(
        ShiftRowsOutput[15]) );
  INV_X1 SubCellInst_SboxInst_2_U2_U1 ( .A(SubCellInst_SboxInst_2_YY_0_), .ZN(
        ShiftRowsOutput[14]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U37 ( .A(new_AGEMA_signal_1768), .B(
        Fresh[14]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U36 ( .A(Fresh[13]), .B(
        SubCellInst_SboxInst_2_Q1), .Z(
        SubCellInst_SboxInst_2_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U35 ( .A(new_AGEMA_signal_1769), .B(
        Fresh[14]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U34 ( .A(Fresh[12]), .B(
        SubCellInst_SboxInst_2_Q1), .Z(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U33 ( .A(Fresh[13]), .B(
        new_AGEMA_signal_1769), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U32 ( .A(new_AGEMA_signal_1768), .B(
        Fresh[12]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U25 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U24 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U23 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U22 ( .A(Fresh[14]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U21 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U19 ( .A(Fresh[13]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U17 ( .A(Fresh[12]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U16 ( .A1(new_AGEMA_signal_1769), 
        .A2(Ciphertext_s2[10]), .ZN(SubCellInst_SboxInst_2_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U15 ( .A1(new_AGEMA_signal_1768), 
        .A2(Ciphertext_s1[10]), .ZN(SubCellInst_SboxInst_2_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_2_Q1), 
        .A2(SubCellInst_SboxInst_2_n3), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_n33), .Z(new_AGEMA_signal_1945) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n32), .B(
        SubCellInst_SboxInst_2_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_n30), .Z(new_AGEMA_signal_1944) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n29), .B(
        SubCellInst_SboxInst_2_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_n27), .Z(SubCellInst_SboxInst_2_T0) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n26), .B(
        SubCellInst_SboxInst_2_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_Q0), .B(SubCellInst_SboxInst_2_T0), .Z(
        SubCellInst_SboxInst_2_Q2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1766), 
        .B(new_AGEMA_signal_1944), .Z(new_AGEMA_signal_2044) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1767), 
        .B(new_AGEMA_signal_1945), .Z(new_AGEMA_signal_2045) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U37 ( .A(new_AGEMA_signal_1770), .B(
        Fresh[17]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U36 ( .A(Fresh[16]), .B(
        SubCellInst_SboxInst_2_Q4), .Z(
        SubCellInst_SboxInst_2_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U35 ( .A(new_AGEMA_signal_1771), .B(
        Fresh[17]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U34 ( .A(Fresh[15]), .B(
        SubCellInst_SboxInst_2_Q4), .Z(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U33 ( .A(Fresh[16]), .B(
        new_AGEMA_signal_1771), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U32 ( .A(new_AGEMA_signal_1770), .B(
        Fresh[15]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U25 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U24 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U23 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U22 ( .A(Fresh[17]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U21 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U19 ( .A(Fresh[16]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U17 ( .A(Fresh[15]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U16 ( .A1(new_AGEMA_signal_1771), 
        .A2(Ciphertext_s2[10]), .ZN(SubCellInst_SboxInst_2_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U15 ( .A1(new_AGEMA_signal_1770), 
        .A2(Ciphertext_s1[10]), .ZN(SubCellInst_SboxInst_2_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_2_Q4), 
        .A2(SubCellInst_SboxInst_2_n3), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_n33), .Z(new_AGEMA_signal_1947) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n32), .B(
        SubCellInst_SboxInst_2_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_n30), .Z(new_AGEMA_signal_1946) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n29), .B(
        SubCellInst_SboxInst_2_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_n27), .Z(SubCellInst_SboxInst_2_T2) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n26), .B(
        SubCellInst_SboxInst_2_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L1), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_Q7) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1948), 
        .B(new_AGEMA_signal_1946), .Z(new_AGEMA_signal_2046) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1949), 
        .B(new_AGEMA_signal_1947), .Z(new_AGEMA_signal_2047) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_XX_2_), .B(SubCellInst_SboxInst_2_T0), .Z(
        SubCellInst_SboxInst_2_L3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1198), 
        .B(new_AGEMA_signal_1944), .Z(new_AGEMA_signal_2048) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1199), 
        .B(new_AGEMA_signal_1945), .Z(new_AGEMA_signal_2049) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L3), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2048), 
        .B(new_AGEMA_signal_1946), .Z(new_AGEMA_signal_2292) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2049), 
        .B(new_AGEMA_signal_1947), .Z(new_AGEMA_signal_2293) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_XX_1_), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1194), 
        .B(new_AGEMA_signal_1946), .Z(new_AGEMA_signal_2172) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1195), 
        .B(new_AGEMA_signal_1947), .Z(new_AGEMA_signal_2173) );
  INV_X1 SubCellInst_SboxInst_3_U3_U1 ( .A(SubCellInst_SboxInst_3_YY_1_), .ZN(
        ShiftRowsOutput[3]) );
  INV_X1 SubCellInst_SboxInst_3_U2_U1 ( .A(SubCellInst_SboxInst_3_YY_0_), .ZN(
        ShiftRowsOutput[2]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U37 ( .A(new_AGEMA_signal_1780), .B(
        Fresh[20]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U36 ( .A(Fresh[19]), .B(
        SubCellInst_SboxInst_3_Q1), .Z(
        SubCellInst_SboxInst_3_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U35 ( .A(new_AGEMA_signal_1781), .B(
        Fresh[20]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U34 ( .A(Fresh[18]), .B(
        SubCellInst_SboxInst_3_Q1), .Z(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U33 ( .A(Fresh[19]), .B(
        new_AGEMA_signal_1781), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U32 ( .A(new_AGEMA_signal_1780), .B(
        Fresh[18]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U25 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U24 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U23 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U22 ( .A(Fresh[20]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U21 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U19 ( .A(Fresh[19]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U17 ( .A(Fresh[18]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U16 ( .A1(new_AGEMA_signal_1781), 
        .A2(Ciphertext_s2[14]), .ZN(SubCellInst_SboxInst_3_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U15 ( .A1(new_AGEMA_signal_1780), 
        .A2(Ciphertext_s1[14]), .ZN(SubCellInst_SboxInst_3_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_3_Q1), 
        .A2(SubCellInst_SboxInst_3_n3), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_n33), .Z(new_AGEMA_signal_1951) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n32), .B(
        SubCellInst_SboxInst_3_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_n30), .Z(new_AGEMA_signal_1950) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n29), .B(
        SubCellInst_SboxInst_3_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_n27), .Z(SubCellInst_SboxInst_3_T0) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n26), .B(
        SubCellInst_SboxInst_3_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_Q0), .B(SubCellInst_SboxInst_3_T0), .Z(
        SubCellInst_SboxInst_3_Q2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1778), 
        .B(new_AGEMA_signal_1950), .Z(new_AGEMA_signal_2052) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1779), 
        .B(new_AGEMA_signal_1951), .Z(new_AGEMA_signal_2053) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U37 ( .A(new_AGEMA_signal_1782), .B(
        Fresh[23]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U36 ( .A(Fresh[22]), .B(
        SubCellInst_SboxInst_3_Q4), .Z(
        SubCellInst_SboxInst_3_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U35 ( .A(new_AGEMA_signal_1783), .B(
        Fresh[23]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U34 ( .A(Fresh[21]), .B(
        SubCellInst_SboxInst_3_Q4), .Z(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U33 ( .A(Fresh[22]), .B(
        new_AGEMA_signal_1783), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U32 ( .A(new_AGEMA_signal_1782), .B(
        Fresh[21]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U25 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U24 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U23 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U22 ( .A(Fresh[23]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U21 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U19 ( .A(Fresh[22]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U17 ( .A(Fresh[21]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U16 ( .A1(new_AGEMA_signal_1783), 
        .A2(Ciphertext_s2[14]), .ZN(SubCellInst_SboxInst_3_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U15 ( .A1(new_AGEMA_signal_1782), 
        .A2(Ciphertext_s1[14]), .ZN(SubCellInst_SboxInst_3_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_3_Q4), 
        .A2(SubCellInst_SboxInst_3_n3), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_n33), .Z(new_AGEMA_signal_1953) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n32), .B(
        SubCellInst_SboxInst_3_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_n30), .Z(new_AGEMA_signal_1952) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n29), .B(
        SubCellInst_SboxInst_3_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_n27), .Z(SubCellInst_SboxInst_3_T2) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n26), .B(
        SubCellInst_SboxInst_3_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L1), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_Q7) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1954), 
        .B(new_AGEMA_signal_1952), .Z(new_AGEMA_signal_2054) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1955), 
        .B(new_AGEMA_signal_1953), .Z(new_AGEMA_signal_2055) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_XX_2_), .B(SubCellInst_SboxInst_3_T0), .Z(
        SubCellInst_SboxInst_3_L3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1210), 
        .B(new_AGEMA_signal_1950), .Z(new_AGEMA_signal_2056) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1211), 
        .B(new_AGEMA_signal_1951), .Z(new_AGEMA_signal_2057) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L3), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2056), 
        .B(new_AGEMA_signal_1952), .Z(new_AGEMA_signal_2296) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2057), 
        .B(new_AGEMA_signal_1953), .Z(new_AGEMA_signal_2297) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_XX_1_), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1206), 
        .B(new_AGEMA_signal_1952), .Z(new_AGEMA_signal_2180) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1207), 
        .B(new_AGEMA_signal_1953), .Z(new_AGEMA_signal_2181) );
  INV_X1 SubCellInst_SboxInst_4_U3_U1 ( .A(SubCellInst_SboxInst_4_YY_1_), .ZN(
        ShiftRowsOutput[27]) );
  INV_X1 SubCellInst_SboxInst_4_U2_U1 ( .A(SubCellInst_SboxInst_4_YY_0_), .ZN(
        ShiftRowsOutput[26]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U37 ( .A(new_AGEMA_signal_1792), .B(
        Fresh[26]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U36 ( .A(Fresh[25]), .B(
        SubCellInst_SboxInst_4_Q1), .Z(
        SubCellInst_SboxInst_4_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U35 ( .A(new_AGEMA_signal_1793), .B(
        Fresh[26]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U34 ( .A(Fresh[24]), .B(
        SubCellInst_SboxInst_4_Q1), .Z(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U33 ( .A(Fresh[25]), .B(
        new_AGEMA_signal_1793), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U32 ( .A(new_AGEMA_signal_1792), .B(
        Fresh[24]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U25 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U24 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U23 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U22 ( .A(Fresh[26]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U21 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U19 ( .A(Fresh[25]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U17 ( .A(Fresh[24]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U16 ( .A1(new_AGEMA_signal_1793), 
        .A2(Ciphertext_s2[18]), .ZN(SubCellInst_SboxInst_4_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U15 ( .A1(new_AGEMA_signal_1792), 
        .A2(Ciphertext_s1[18]), .ZN(SubCellInst_SboxInst_4_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_4_Q1), 
        .A2(SubCellInst_SboxInst_4_n3), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_n33), .Z(new_AGEMA_signal_1957) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n32), .B(
        SubCellInst_SboxInst_4_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_n30), .Z(new_AGEMA_signal_1956) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n29), .B(
        SubCellInst_SboxInst_4_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_n27), .Z(SubCellInst_SboxInst_4_T0) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n26), .B(
        SubCellInst_SboxInst_4_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_Q0), .B(SubCellInst_SboxInst_4_T0), .Z(
        SubCellInst_SboxInst_4_Q2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1790), 
        .B(new_AGEMA_signal_1956), .Z(new_AGEMA_signal_2060) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1791), 
        .B(new_AGEMA_signal_1957), .Z(new_AGEMA_signal_2061) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U37 ( .A(new_AGEMA_signal_1794), .B(
        Fresh[29]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U36 ( .A(Fresh[28]), .B(
        SubCellInst_SboxInst_4_Q4), .Z(
        SubCellInst_SboxInst_4_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U35 ( .A(new_AGEMA_signal_1795), .B(
        Fresh[29]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U34 ( .A(Fresh[27]), .B(
        SubCellInst_SboxInst_4_Q4), .Z(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U33 ( .A(Fresh[28]), .B(
        new_AGEMA_signal_1795), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U32 ( .A(new_AGEMA_signal_1794), .B(
        Fresh[27]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U25 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U24 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U23 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U22 ( .A(Fresh[29]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U21 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U19 ( .A(Fresh[28]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U17 ( .A(Fresh[27]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U16 ( .A1(new_AGEMA_signal_1795), 
        .A2(Ciphertext_s2[18]), .ZN(SubCellInst_SboxInst_4_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U15 ( .A1(new_AGEMA_signal_1794), 
        .A2(Ciphertext_s1[18]), .ZN(SubCellInst_SboxInst_4_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_4_Q4), 
        .A2(SubCellInst_SboxInst_4_n3), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_n33), .Z(new_AGEMA_signal_1959) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n32), .B(
        SubCellInst_SboxInst_4_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_n30), .Z(new_AGEMA_signal_1958) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n29), .B(
        SubCellInst_SboxInst_4_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_n27), .Z(SubCellInst_SboxInst_4_T2) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n26), .B(
        SubCellInst_SboxInst_4_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L1), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_Q7) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1960), 
        .B(new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2062) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1961), 
        .B(new_AGEMA_signal_1959), .Z(new_AGEMA_signal_2063) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_XX_2_), .B(SubCellInst_SboxInst_4_T0), .Z(
        SubCellInst_SboxInst_4_L3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1222), 
        .B(new_AGEMA_signal_1956), .Z(new_AGEMA_signal_2064) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1223), 
        .B(new_AGEMA_signal_1957), .Z(new_AGEMA_signal_2065) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L3), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2064), 
        .B(new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2300) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2065), 
        .B(new_AGEMA_signal_1959), .Z(new_AGEMA_signal_2301) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_XX_1_), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1218), 
        .B(new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2188) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1219), 
        .B(new_AGEMA_signal_1959), .Z(new_AGEMA_signal_2189) );
  INV_X1 SubCellInst_SboxInst_5_U3_U1 ( .A(SubCellInst_SboxInst_5_YY_1_), .ZN(
        ShiftRowsOutput[31]) );
  INV_X1 SubCellInst_SboxInst_5_U2_U1 ( .A(SubCellInst_SboxInst_5_YY_0_), .ZN(
        ShiftRowsOutput[30]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U37 ( .A(new_AGEMA_signal_1804), .B(
        Fresh[32]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U36 ( .A(Fresh[31]), .B(
        SubCellInst_SboxInst_5_Q1), .Z(
        SubCellInst_SboxInst_5_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U35 ( .A(new_AGEMA_signal_1805), .B(
        Fresh[32]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U34 ( .A(Fresh[30]), .B(
        SubCellInst_SboxInst_5_Q1), .Z(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U33 ( .A(Fresh[31]), .B(
        new_AGEMA_signal_1805), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U32 ( .A(new_AGEMA_signal_1804), .B(
        Fresh[30]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U25 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U24 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U23 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U22 ( .A(Fresh[32]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U21 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U19 ( .A(Fresh[31]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U17 ( .A(Fresh[30]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U16 ( .A1(new_AGEMA_signal_1805), 
        .A2(Ciphertext_s2[22]), .ZN(SubCellInst_SboxInst_5_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U15 ( .A1(new_AGEMA_signal_1804), 
        .A2(Ciphertext_s1[22]), .ZN(SubCellInst_SboxInst_5_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_5_Q1), 
        .A2(SubCellInst_SboxInst_5_n3), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_n33), .Z(new_AGEMA_signal_1963) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n32), .B(
        SubCellInst_SboxInst_5_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_n30), .Z(new_AGEMA_signal_1962) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n29), .B(
        SubCellInst_SboxInst_5_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_n27), .Z(SubCellInst_SboxInst_5_T0) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n26), .B(
        SubCellInst_SboxInst_5_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_Q0), .B(SubCellInst_SboxInst_5_T0), .Z(
        SubCellInst_SboxInst_5_Q2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1802), 
        .B(new_AGEMA_signal_1962), .Z(new_AGEMA_signal_2068) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1803), 
        .B(new_AGEMA_signal_1963), .Z(new_AGEMA_signal_2069) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U37 ( .A(new_AGEMA_signal_1806), .B(
        Fresh[35]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U36 ( .A(Fresh[34]), .B(
        SubCellInst_SboxInst_5_Q4), .Z(
        SubCellInst_SboxInst_5_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U35 ( .A(new_AGEMA_signal_1807), .B(
        Fresh[35]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U34 ( .A(Fresh[33]), .B(
        SubCellInst_SboxInst_5_Q4), .Z(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U33 ( .A(Fresh[34]), .B(
        new_AGEMA_signal_1807), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U32 ( .A(new_AGEMA_signal_1806), .B(
        Fresh[33]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U25 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U24 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U23 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U22 ( .A(Fresh[35]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U21 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U19 ( .A(Fresh[34]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U17 ( .A(Fresh[33]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U16 ( .A1(new_AGEMA_signal_1807), 
        .A2(Ciphertext_s2[22]), .ZN(SubCellInst_SboxInst_5_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U15 ( .A1(new_AGEMA_signal_1806), 
        .A2(Ciphertext_s1[22]), .ZN(SubCellInst_SboxInst_5_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_5_Q4), 
        .A2(SubCellInst_SboxInst_5_n3), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_n33), .Z(new_AGEMA_signal_1965) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n32), .B(
        SubCellInst_SboxInst_5_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_n30), .Z(new_AGEMA_signal_1964) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n29), .B(
        SubCellInst_SboxInst_5_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_n27), .Z(SubCellInst_SboxInst_5_T2) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n26), .B(
        SubCellInst_SboxInst_5_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L1), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_Q7) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1966), 
        .B(new_AGEMA_signal_1964), .Z(new_AGEMA_signal_2070) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1967), 
        .B(new_AGEMA_signal_1965), .Z(new_AGEMA_signal_2071) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_XX_2_), .B(SubCellInst_SboxInst_5_T0), .Z(
        SubCellInst_SboxInst_5_L3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1234), 
        .B(new_AGEMA_signal_1962), .Z(new_AGEMA_signal_2072) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1235), 
        .B(new_AGEMA_signal_1963), .Z(new_AGEMA_signal_2073) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L3), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2072), 
        .B(new_AGEMA_signal_1964), .Z(new_AGEMA_signal_2304) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2073), 
        .B(new_AGEMA_signal_1965), .Z(new_AGEMA_signal_2305) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_XX_1_), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1230), 
        .B(new_AGEMA_signal_1964), .Z(new_AGEMA_signal_2196) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1231), 
        .B(new_AGEMA_signal_1965), .Z(new_AGEMA_signal_2197) );
  INV_X1 SubCellInst_SboxInst_6_U3_U1 ( .A(SubCellInst_SboxInst_6_YY_1_), .ZN(
        ShiftRowsOutput[19]) );
  INV_X1 SubCellInst_SboxInst_6_U2_U1 ( .A(SubCellInst_SboxInst_6_YY_0_), .ZN(
        ShiftRowsOutput[18]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U37 ( .A(new_AGEMA_signal_1816), .B(
        Fresh[38]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U36 ( .A(Fresh[37]), .B(
        SubCellInst_SboxInst_6_Q1), .Z(
        SubCellInst_SboxInst_6_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U35 ( .A(new_AGEMA_signal_1817), .B(
        Fresh[38]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U34 ( .A(Fresh[36]), .B(
        SubCellInst_SboxInst_6_Q1), .Z(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U33 ( .A(Fresh[37]), .B(
        new_AGEMA_signal_1817), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U32 ( .A(new_AGEMA_signal_1816), .B(
        Fresh[36]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U25 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U24 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U23 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U22 ( .A(Fresh[38]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U21 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U19 ( .A(Fresh[37]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U17 ( .A(Fresh[36]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U16 ( .A1(new_AGEMA_signal_1817), 
        .A2(Ciphertext_s2[26]), .ZN(SubCellInst_SboxInst_6_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U15 ( .A1(new_AGEMA_signal_1816), 
        .A2(Ciphertext_s1[26]), .ZN(SubCellInst_SboxInst_6_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_6_Q1), 
        .A2(SubCellInst_SboxInst_6_n3), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_n33), .Z(new_AGEMA_signal_1969) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n32), .B(
        SubCellInst_SboxInst_6_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_n30), .Z(new_AGEMA_signal_1968) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n29), .B(
        SubCellInst_SboxInst_6_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_n27), .Z(SubCellInst_SboxInst_6_T0) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n26), .B(
        SubCellInst_SboxInst_6_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_Q0), .B(SubCellInst_SboxInst_6_T0), .Z(
        SubCellInst_SboxInst_6_Q2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1814), 
        .B(new_AGEMA_signal_1968), .Z(new_AGEMA_signal_2076) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1815), 
        .B(new_AGEMA_signal_1969), .Z(new_AGEMA_signal_2077) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U37 ( .A(new_AGEMA_signal_1818), .B(
        Fresh[41]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U36 ( .A(Fresh[40]), .B(
        SubCellInst_SboxInst_6_Q4), .Z(
        SubCellInst_SboxInst_6_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U35 ( .A(new_AGEMA_signal_1819), .B(
        Fresh[41]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U34 ( .A(Fresh[39]), .B(
        SubCellInst_SboxInst_6_Q4), .Z(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U33 ( .A(Fresh[40]), .B(
        new_AGEMA_signal_1819), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U32 ( .A(new_AGEMA_signal_1818), .B(
        Fresh[39]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U25 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U24 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U23 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U22 ( .A(Fresh[41]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U21 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U19 ( .A(Fresh[40]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U17 ( .A(Fresh[39]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U16 ( .A1(new_AGEMA_signal_1819), 
        .A2(Ciphertext_s2[26]), .ZN(SubCellInst_SboxInst_6_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U15 ( .A1(new_AGEMA_signal_1818), 
        .A2(Ciphertext_s1[26]), .ZN(SubCellInst_SboxInst_6_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_6_Q4), 
        .A2(SubCellInst_SboxInst_6_n3), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_n33), .Z(new_AGEMA_signal_1971) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n32), .B(
        SubCellInst_SboxInst_6_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_n30), .Z(new_AGEMA_signal_1970) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n29), .B(
        SubCellInst_SboxInst_6_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_n27), .Z(SubCellInst_SboxInst_6_T2) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n26), .B(
        SubCellInst_SboxInst_6_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L1), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_Q7) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1972), 
        .B(new_AGEMA_signal_1970), .Z(new_AGEMA_signal_2078) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1973), 
        .B(new_AGEMA_signal_1971), .Z(new_AGEMA_signal_2079) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_XX_2_), .B(SubCellInst_SboxInst_6_T0), .Z(
        SubCellInst_SboxInst_6_L3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1246), 
        .B(new_AGEMA_signal_1968), .Z(new_AGEMA_signal_2080) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1247), 
        .B(new_AGEMA_signal_1969), .Z(new_AGEMA_signal_2081) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L3), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2080), 
        .B(new_AGEMA_signal_1970), .Z(new_AGEMA_signal_2308) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2081), 
        .B(new_AGEMA_signal_1971), .Z(new_AGEMA_signal_2309) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_XX_1_), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1242), 
        .B(new_AGEMA_signal_1970), .Z(new_AGEMA_signal_2204) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1243), 
        .B(new_AGEMA_signal_1971), .Z(new_AGEMA_signal_2205) );
  INV_X1 SubCellInst_SboxInst_7_U3_U1 ( .A(SubCellInst_SboxInst_7_YY_1_), .ZN(
        ShiftRowsOutput[23]) );
  INV_X1 SubCellInst_SboxInst_7_U2_U1 ( .A(SubCellInst_SboxInst_7_YY_0_), .ZN(
        ShiftRowsOutput[22]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U37 ( .A(new_AGEMA_signal_1828), .B(
        Fresh[44]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U36 ( .A(Fresh[43]), .B(
        SubCellInst_SboxInst_7_Q1), .Z(
        SubCellInst_SboxInst_7_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U35 ( .A(new_AGEMA_signal_1829), .B(
        Fresh[44]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U34 ( .A(Fresh[42]), .B(
        SubCellInst_SboxInst_7_Q1), .Z(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U33 ( .A(Fresh[43]), .B(
        new_AGEMA_signal_1829), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U32 ( .A(new_AGEMA_signal_1828), .B(
        Fresh[42]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U25 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U24 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U23 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U22 ( .A(Fresh[44]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U21 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U19 ( .A(Fresh[43]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U17 ( .A(Fresh[42]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U16 ( .A1(new_AGEMA_signal_1829), 
        .A2(Ciphertext_s2[30]), .ZN(SubCellInst_SboxInst_7_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U15 ( .A1(new_AGEMA_signal_1828), 
        .A2(Ciphertext_s1[30]), .ZN(SubCellInst_SboxInst_7_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_7_Q1), 
        .A2(SubCellInst_SboxInst_7_n3), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_n33), .Z(new_AGEMA_signal_1975) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n32), .B(
        SubCellInst_SboxInst_7_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_n30), .Z(new_AGEMA_signal_1974) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n29), .B(
        SubCellInst_SboxInst_7_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_n27), .Z(SubCellInst_SboxInst_7_T0) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n26), .B(
        SubCellInst_SboxInst_7_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_Q0), .B(SubCellInst_SboxInst_7_T0), .Z(
        SubCellInst_SboxInst_7_Q2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1826), 
        .B(new_AGEMA_signal_1974), .Z(new_AGEMA_signal_2084) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1827), 
        .B(new_AGEMA_signal_1975), .Z(new_AGEMA_signal_2085) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U37 ( .A(new_AGEMA_signal_1830), .B(
        Fresh[47]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U36 ( .A(Fresh[46]), .B(
        SubCellInst_SboxInst_7_Q4), .Z(
        SubCellInst_SboxInst_7_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U35 ( .A(new_AGEMA_signal_1831), .B(
        Fresh[47]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U34 ( .A(Fresh[45]), .B(
        SubCellInst_SboxInst_7_Q4), .Z(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U33 ( .A(Fresh[46]), .B(
        new_AGEMA_signal_1831), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U32 ( .A(new_AGEMA_signal_1830), .B(
        Fresh[45]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U25 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U24 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U23 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U22 ( .A(Fresh[47]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U21 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U19 ( .A(Fresh[46]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U17 ( .A(Fresh[45]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U16 ( .A1(new_AGEMA_signal_1831), 
        .A2(Ciphertext_s2[30]), .ZN(SubCellInst_SboxInst_7_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U15 ( .A1(new_AGEMA_signal_1830), 
        .A2(Ciphertext_s1[30]), .ZN(SubCellInst_SboxInst_7_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_7_Q4), 
        .A2(SubCellInst_SboxInst_7_n3), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_n33), .Z(new_AGEMA_signal_1977) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n32), .B(
        SubCellInst_SboxInst_7_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_n30), .Z(new_AGEMA_signal_1976) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n29), .B(
        SubCellInst_SboxInst_7_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_n27), .Z(SubCellInst_SboxInst_7_T2) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n26), .B(
        SubCellInst_SboxInst_7_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L1), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_Q7) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1978), 
        .B(new_AGEMA_signal_1976), .Z(new_AGEMA_signal_2086) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1979), 
        .B(new_AGEMA_signal_1977), .Z(new_AGEMA_signal_2087) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_XX_2_), .B(SubCellInst_SboxInst_7_T0), .Z(
        SubCellInst_SboxInst_7_L3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1258), 
        .B(new_AGEMA_signal_1974), .Z(new_AGEMA_signal_2088) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1259), 
        .B(new_AGEMA_signal_1975), .Z(new_AGEMA_signal_2089) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L3), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2088), 
        .B(new_AGEMA_signal_1976), .Z(new_AGEMA_signal_2312) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2089), 
        .B(new_AGEMA_signal_1977), .Z(new_AGEMA_signal_2313) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_XX_1_), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1254), 
        .B(new_AGEMA_signal_1976), .Z(new_AGEMA_signal_2212) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1255), 
        .B(new_AGEMA_signal_1977), .Z(new_AGEMA_signal_2213) );
  INV_X1 SubCellInst_SboxInst_8_U3_U1 ( .A(SubCellInst_SboxInst_8_YY_1_), .ZN(
        AddRoundConstantOutput[35]) );
  INV_X1 SubCellInst_SboxInst_8_U2_U1 ( .A(SubCellInst_SboxInst_8_YY_0_), .ZN(
        AddRoundConstantOutput[34]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U37 ( .A(new_AGEMA_signal_1840), .B(
        Fresh[50]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U36 ( .A(Fresh[49]), .B(
        SubCellInst_SboxInst_8_Q1), .Z(
        SubCellInst_SboxInst_8_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U35 ( .A(new_AGEMA_signal_1841), .B(
        Fresh[50]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U34 ( .A(Fresh[48]), .B(
        SubCellInst_SboxInst_8_Q1), .Z(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U33 ( .A(Fresh[49]), .B(
        new_AGEMA_signal_1841), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U32 ( .A(new_AGEMA_signal_1840), .B(
        Fresh[48]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U25 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U24 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U23 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U22 ( .A(Fresh[50]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U21 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U19 ( .A(Fresh[49]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U17 ( .A(Fresh[48]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U16 ( .A1(new_AGEMA_signal_1841), 
        .A2(Ciphertext_s2[34]), .ZN(SubCellInst_SboxInst_8_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U15 ( .A1(new_AGEMA_signal_1840), 
        .A2(Ciphertext_s1[34]), .ZN(SubCellInst_SboxInst_8_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_8_Q1), 
        .A2(SubCellInst_SboxInst_8_n3), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_n33), .Z(new_AGEMA_signal_1981) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n32), .B(
        SubCellInst_SboxInst_8_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_n30), .Z(new_AGEMA_signal_1980) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n29), .B(
        SubCellInst_SboxInst_8_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_n27), .Z(SubCellInst_SboxInst_8_T0) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n26), .B(
        SubCellInst_SboxInst_8_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_Q0), .B(SubCellInst_SboxInst_8_T0), .Z(
        SubCellInst_SboxInst_8_Q2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1838), 
        .B(new_AGEMA_signal_1980), .Z(new_AGEMA_signal_2092) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1839), 
        .B(new_AGEMA_signal_1981), .Z(new_AGEMA_signal_2093) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U37 ( .A(new_AGEMA_signal_1842), .B(
        Fresh[53]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U36 ( .A(Fresh[52]), .B(
        SubCellInst_SboxInst_8_Q4), .Z(
        SubCellInst_SboxInst_8_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U35 ( .A(new_AGEMA_signal_1843), .B(
        Fresh[53]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U34 ( .A(Fresh[51]), .B(
        SubCellInst_SboxInst_8_Q4), .Z(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U33 ( .A(Fresh[52]), .B(
        new_AGEMA_signal_1843), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U32 ( .A(new_AGEMA_signal_1842), .B(
        Fresh[51]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U25 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U24 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U23 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U22 ( .A(Fresh[53]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U21 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U19 ( .A(Fresh[52]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U17 ( .A(Fresh[51]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U16 ( .A1(new_AGEMA_signal_1843), 
        .A2(Ciphertext_s2[34]), .ZN(SubCellInst_SboxInst_8_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U15 ( .A1(new_AGEMA_signal_1842), 
        .A2(Ciphertext_s1[34]), .ZN(SubCellInst_SboxInst_8_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_8_Q4), 
        .A2(SubCellInst_SboxInst_8_n3), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_n33), .Z(new_AGEMA_signal_1983) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n32), .B(
        SubCellInst_SboxInst_8_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_n30), .Z(new_AGEMA_signal_1982) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n29), .B(
        SubCellInst_SboxInst_8_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_n27), .Z(SubCellInst_SboxInst_8_T2) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n26), .B(
        SubCellInst_SboxInst_8_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L1), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_Q7) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1984), 
        .B(new_AGEMA_signal_1982), .Z(new_AGEMA_signal_2094) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1985), 
        .B(new_AGEMA_signal_1983), .Z(new_AGEMA_signal_2095) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_XX_2_), .B(SubCellInst_SboxInst_8_T0), .Z(
        SubCellInst_SboxInst_8_L3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1270), 
        .B(new_AGEMA_signal_1980), .Z(new_AGEMA_signal_2096) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1271), 
        .B(new_AGEMA_signal_1981), .Z(new_AGEMA_signal_2097) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L3), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2096), 
        .B(new_AGEMA_signal_1982), .Z(new_AGEMA_signal_2316) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2097), 
        .B(new_AGEMA_signal_1983), .Z(new_AGEMA_signal_2317) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_XX_1_), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1266), 
        .B(new_AGEMA_signal_1982), .Z(new_AGEMA_signal_2220) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1267), 
        .B(new_AGEMA_signal_1983), .Z(new_AGEMA_signal_2221) );
  INV_X1 SubCellInst_SboxInst_9_U3_U1 ( .A(SubCellInst_SboxInst_9_YY_1_), .ZN(
        AddRoundConstantOutput[39]) );
  INV_X1 SubCellInst_SboxInst_9_U2_U1 ( .A(SubCellInst_SboxInst_9_YY_0_), .ZN(
        AddRoundConstantOutput[38]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U37 ( .A(new_AGEMA_signal_1852), .B(
        Fresh[56]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U36 ( .A(Fresh[55]), .B(
        SubCellInst_SboxInst_9_Q1), .Z(
        SubCellInst_SboxInst_9_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U35 ( .A(new_AGEMA_signal_1853), .B(
        Fresh[56]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U34 ( .A(Fresh[54]), .B(
        SubCellInst_SboxInst_9_Q1), .Z(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U33 ( .A(Fresh[55]), .B(
        new_AGEMA_signal_1853), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U32 ( .A(new_AGEMA_signal_1852), .B(
        Fresh[54]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U25 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U24 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U23 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U22 ( .A(Fresh[56]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U21 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U19 ( .A(Fresh[55]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U17 ( .A(Fresh[54]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U16 ( .A1(new_AGEMA_signal_1853), 
        .A2(Ciphertext_s2[38]), .ZN(SubCellInst_SboxInst_9_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U15 ( .A1(new_AGEMA_signal_1852), 
        .A2(Ciphertext_s1[38]), .ZN(SubCellInst_SboxInst_9_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_9_Q1), 
        .A2(SubCellInst_SboxInst_9_n3), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_n33), .Z(new_AGEMA_signal_1987) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n32), .B(
        SubCellInst_SboxInst_9_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_n30), .Z(new_AGEMA_signal_1986) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n29), .B(
        SubCellInst_SboxInst_9_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_n27), .Z(SubCellInst_SboxInst_9_T0) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n26), .B(
        SubCellInst_SboxInst_9_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_Q0), .B(SubCellInst_SboxInst_9_T0), .Z(
        SubCellInst_SboxInst_9_Q2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1850), 
        .B(new_AGEMA_signal_1986), .Z(new_AGEMA_signal_2100) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1851), 
        .B(new_AGEMA_signal_1987), .Z(new_AGEMA_signal_2101) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U37 ( .A(new_AGEMA_signal_1854), .B(
        Fresh[59]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U36 ( .A(Fresh[58]), .B(
        SubCellInst_SboxInst_9_Q4), .Z(
        SubCellInst_SboxInst_9_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U35 ( .A(new_AGEMA_signal_1855), .B(
        Fresh[59]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U34 ( .A(Fresh[57]), .B(
        SubCellInst_SboxInst_9_Q4), .Z(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U33 ( .A(Fresh[58]), .B(
        new_AGEMA_signal_1855), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U32 ( .A(new_AGEMA_signal_1854), .B(
        Fresh[57]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U25 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U24 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U23 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U22 ( .A(Fresh[59]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U21 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U19 ( .A(Fresh[58]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U17 ( .A(Fresh[57]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U16 ( .A1(new_AGEMA_signal_1855), 
        .A2(Ciphertext_s2[38]), .ZN(SubCellInst_SboxInst_9_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U15 ( .A1(new_AGEMA_signal_1854), 
        .A2(Ciphertext_s1[38]), .ZN(SubCellInst_SboxInst_9_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_9_Q4), 
        .A2(SubCellInst_SboxInst_9_n3), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_n33), .Z(new_AGEMA_signal_1989) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n32), .B(
        SubCellInst_SboxInst_9_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_n30), .Z(new_AGEMA_signal_1988) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n29), .B(
        SubCellInst_SboxInst_9_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_n27), .Z(SubCellInst_SboxInst_9_T2) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n26), .B(
        SubCellInst_SboxInst_9_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L1), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_Q7) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1990), 
        .B(new_AGEMA_signal_1988), .Z(new_AGEMA_signal_2102) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1991), 
        .B(new_AGEMA_signal_1989), .Z(new_AGEMA_signal_2103) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_XX_2_), .B(SubCellInst_SboxInst_9_T0), .Z(
        SubCellInst_SboxInst_9_L3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1282), 
        .B(new_AGEMA_signal_1986), .Z(new_AGEMA_signal_2104) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1283), 
        .B(new_AGEMA_signal_1987), .Z(new_AGEMA_signal_2105) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L3), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2104), 
        .B(new_AGEMA_signal_1988), .Z(new_AGEMA_signal_2320) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2105), 
        .B(new_AGEMA_signal_1989), .Z(new_AGEMA_signal_2321) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_XX_1_), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1278), 
        .B(new_AGEMA_signal_1988), .Z(new_AGEMA_signal_2228) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1279), 
        .B(new_AGEMA_signal_1989), .Z(new_AGEMA_signal_2229) );
  INV_X1 SubCellInst_SboxInst_10_U3_U1 ( .A(SubCellInst_SboxInst_10_YY_1_), 
        .ZN(AddRoundConstantOutput[43]) );
  INV_X1 SubCellInst_SboxInst_10_U2_U1 ( .A(SubCellInst_SboxInst_10_YY_0_), 
        .ZN(AddRoundConstantOutput[42]) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U37 ( .A(new_AGEMA_signal_1864), .B(
        Fresh[62]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U36 ( .A(Fresh[61]), .B(
        SubCellInst_SboxInst_10_Q1), .Z(
        SubCellInst_SboxInst_10_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U35 ( .A(new_AGEMA_signal_1865), .B(
        Fresh[62]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U34 ( .A(Fresh[60]), .B(
        SubCellInst_SboxInst_10_Q1), .Z(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U33 ( .A(Fresh[61]), .B(
        new_AGEMA_signal_1865), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U32 ( .A(new_AGEMA_signal_1864), .B(
        Fresh[60]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U25 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U24 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U23 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U22 ( .A(Fresh[62]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U21 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U19 ( .A(Fresh[61]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U17 ( .A(Fresh[60]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U16 ( .A1(new_AGEMA_signal_1865), 
        .A2(Ciphertext_s2[42]), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U15 ( .A1(new_AGEMA_signal_1864), 
        .A2(Ciphertext_s1[42]), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_10_Q1), .A2(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_n33), .Z(new_AGEMA_signal_1993) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n32), .B(
        SubCellInst_SboxInst_10_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_n30), .Z(new_AGEMA_signal_1992) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n29), .B(
        SubCellInst_SboxInst_10_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_n27), .Z(SubCellInst_SboxInst_10_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n26), .B(
        SubCellInst_SboxInst_10_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_Q0), .B(SubCellInst_SboxInst_10_T0), .Z(
        SubCellInst_SboxInst_10_Q2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1862), 
        .B(new_AGEMA_signal_1992), .Z(new_AGEMA_signal_2108) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1863), 
        .B(new_AGEMA_signal_1993), .Z(new_AGEMA_signal_2109) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U37 ( .A(new_AGEMA_signal_1866), .B(
        Fresh[65]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U36 ( .A(Fresh[64]), .B(
        SubCellInst_SboxInst_10_Q4), .Z(
        SubCellInst_SboxInst_10_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U35 ( .A(new_AGEMA_signal_1867), .B(
        Fresh[65]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U34 ( .A(Fresh[63]), .B(
        SubCellInst_SboxInst_10_Q4), .Z(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U33 ( .A(Fresh[64]), .B(
        new_AGEMA_signal_1867), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U32 ( .A(new_AGEMA_signal_1866), .B(
        Fresh[63]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U25 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U24 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U23 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U22 ( .A(Fresh[65]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U21 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U19 ( .A(Fresh[64]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U17 ( .A(Fresh[63]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U16 ( .A1(new_AGEMA_signal_1867), 
        .A2(Ciphertext_s2[42]), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U15 ( .A1(new_AGEMA_signal_1866), 
        .A2(Ciphertext_s1[42]), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_10_Q4), .A2(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_n33), .Z(new_AGEMA_signal_1995) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n32), .B(
        SubCellInst_SboxInst_10_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_n30), .Z(new_AGEMA_signal_1994) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n29), .B(
        SubCellInst_SboxInst_10_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_n27), .Z(SubCellInst_SboxInst_10_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n26), .B(
        SubCellInst_SboxInst_10_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L1), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_Q7) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1996), 
        .B(new_AGEMA_signal_1994), .Z(new_AGEMA_signal_2110) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1997), 
        .B(new_AGEMA_signal_1995), .Z(new_AGEMA_signal_2111) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_XX_2_), .B(SubCellInst_SboxInst_10_T0), .Z(
        SubCellInst_SboxInst_10_L3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1294), .B(new_AGEMA_signal_1992), .Z(new_AGEMA_signal_2112) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1295), .B(new_AGEMA_signal_1993), .Z(new_AGEMA_signal_2113) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L3), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2112), .B(new_AGEMA_signal_1994), .Z(new_AGEMA_signal_2324) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2113), .B(new_AGEMA_signal_1995), .Z(new_AGEMA_signal_2325) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_XX_1_), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1290), .B(new_AGEMA_signal_1994), .Z(new_AGEMA_signal_2236) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1291), .B(new_AGEMA_signal_1995), .Z(new_AGEMA_signal_2237) );
  INV_X1 SubCellInst_SboxInst_11_U3_U1 ( .A(SubCellInst_SboxInst_11_YY_1_), 
        .ZN(SubCellOutput_47) );
  INV_X1 SubCellInst_SboxInst_11_U2_U1 ( .A(SubCellInst_SboxInst_11_YY_0_), 
        .ZN(SubCellOutput_46) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U37 ( .A(new_AGEMA_signal_1876), .B(
        Fresh[68]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U36 ( .A(Fresh[67]), .B(
        SubCellInst_SboxInst_11_Q1), .Z(
        SubCellInst_SboxInst_11_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U35 ( .A(new_AGEMA_signal_1877), .B(
        Fresh[68]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U34 ( .A(Fresh[66]), .B(
        SubCellInst_SboxInst_11_Q1), .Z(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U33 ( .A(Fresh[67]), .B(
        new_AGEMA_signal_1877), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U32 ( .A(new_AGEMA_signal_1876), .B(
        Fresh[66]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U25 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U24 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U23 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U22 ( .A(Fresh[68]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U21 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U19 ( .A(Fresh[67]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U17 ( .A(Fresh[66]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U16 ( .A1(new_AGEMA_signal_1877), 
        .A2(Ciphertext_s2[46]), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U15 ( .A1(new_AGEMA_signal_1876), 
        .A2(Ciphertext_s1[46]), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_11_Q1), .A2(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_n33), .Z(new_AGEMA_signal_1999) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n32), .B(
        SubCellInst_SboxInst_11_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_n30), .Z(new_AGEMA_signal_1998) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n29), .B(
        SubCellInst_SboxInst_11_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_n27), .Z(SubCellInst_SboxInst_11_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n26), .B(
        SubCellInst_SboxInst_11_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_Q0), .B(SubCellInst_SboxInst_11_T0), .Z(
        SubCellInst_SboxInst_11_Q2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1874), 
        .B(new_AGEMA_signal_1998), .Z(new_AGEMA_signal_2116) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1875), 
        .B(new_AGEMA_signal_1999), .Z(new_AGEMA_signal_2117) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U37 ( .A(new_AGEMA_signal_1878), .B(
        Fresh[71]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U36 ( .A(Fresh[70]), .B(
        SubCellInst_SboxInst_11_Q4), .Z(
        SubCellInst_SboxInst_11_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U35 ( .A(new_AGEMA_signal_1879), .B(
        Fresh[71]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U34 ( .A(Fresh[69]), .B(
        SubCellInst_SboxInst_11_Q4), .Z(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U33 ( .A(Fresh[70]), .B(
        new_AGEMA_signal_1879), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U32 ( .A(new_AGEMA_signal_1878), .B(
        Fresh[69]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U25 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U24 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U23 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U22 ( .A(Fresh[71]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U21 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U19 ( .A(Fresh[70]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U17 ( .A(Fresh[69]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U16 ( .A1(new_AGEMA_signal_1879), 
        .A2(Ciphertext_s2[46]), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U15 ( .A1(new_AGEMA_signal_1878), 
        .A2(Ciphertext_s1[46]), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_11_Q4), .A2(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_n33), .Z(new_AGEMA_signal_2001) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n32), .B(
        SubCellInst_SboxInst_11_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_n30), .Z(new_AGEMA_signal_2000) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n29), .B(
        SubCellInst_SboxInst_11_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_n27), .Z(SubCellInst_SboxInst_11_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n26), .B(
        SubCellInst_SboxInst_11_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L1), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_Q7) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2002), 
        .B(new_AGEMA_signal_2000), .Z(new_AGEMA_signal_2118) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2003), 
        .B(new_AGEMA_signal_2001), .Z(new_AGEMA_signal_2119) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_XX_2_), .B(SubCellInst_SboxInst_11_T0), .Z(
        SubCellInst_SboxInst_11_L3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1306), .B(new_AGEMA_signal_1998), .Z(new_AGEMA_signal_2120) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1307), .B(new_AGEMA_signal_1999), .Z(new_AGEMA_signal_2121) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L3), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2120), .B(new_AGEMA_signal_2000), .Z(new_AGEMA_signal_2328) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2121), .B(new_AGEMA_signal_2001), .Z(new_AGEMA_signal_2329) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_XX_1_), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1302), .B(new_AGEMA_signal_2000), .Z(new_AGEMA_signal_2244) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1303), .B(new_AGEMA_signal_2001), .Z(new_AGEMA_signal_2245) );
  INV_X1 SubCellInst_SboxInst_12_U3_U1 ( .A(SubCellInst_SboxInst_12_YY_1_), 
        .ZN(AddRoundConstantOutput[51]) );
  INV_X1 SubCellInst_SboxInst_12_U2_U1 ( .A(SubCellInst_SboxInst_12_YY_0_), 
        .ZN(AddRoundConstantOutput[50]) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U37 ( .A(new_AGEMA_signal_1888), .B(
        Fresh[74]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U36 ( .A(Fresh[73]), .B(
        SubCellInst_SboxInst_12_Q1), .Z(
        SubCellInst_SboxInst_12_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U35 ( .A(new_AGEMA_signal_1889), .B(
        Fresh[74]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U34 ( .A(Fresh[72]), .B(
        SubCellInst_SboxInst_12_Q1), .Z(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U33 ( .A(Fresh[73]), .B(
        new_AGEMA_signal_1889), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U32 ( .A(new_AGEMA_signal_1888), .B(
        Fresh[72]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U25 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U24 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U23 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U22 ( .A(Fresh[74]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U21 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U19 ( .A(Fresh[73]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U17 ( .A(Fresh[72]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U16 ( .A1(new_AGEMA_signal_1889), 
        .A2(Ciphertext_s2[50]), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U15 ( .A1(new_AGEMA_signal_1888), 
        .A2(Ciphertext_s1[50]), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_12_Q1), .A2(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_n33), .Z(new_AGEMA_signal_2005) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n32), .B(
        SubCellInst_SboxInst_12_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_n30), .Z(new_AGEMA_signal_2004) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n29), .B(
        SubCellInst_SboxInst_12_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_n27), .Z(SubCellInst_SboxInst_12_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n26), .B(
        SubCellInst_SboxInst_12_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_Q0), .B(SubCellInst_SboxInst_12_T0), .Z(
        SubCellInst_SboxInst_12_Q2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1886), 
        .B(new_AGEMA_signal_2004), .Z(new_AGEMA_signal_2124) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1887), 
        .B(new_AGEMA_signal_2005), .Z(new_AGEMA_signal_2125) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U37 ( .A(new_AGEMA_signal_1890), .B(
        Fresh[77]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U36 ( .A(Fresh[76]), .B(
        SubCellInst_SboxInst_12_Q4), .Z(
        SubCellInst_SboxInst_12_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U35 ( .A(new_AGEMA_signal_1891), .B(
        Fresh[77]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U34 ( .A(Fresh[75]), .B(
        SubCellInst_SboxInst_12_Q4), .Z(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U33 ( .A(Fresh[76]), .B(
        new_AGEMA_signal_1891), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U32 ( .A(new_AGEMA_signal_1890), .B(
        Fresh[75]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U25 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U24 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U23 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U22 ( .A(Fresh[77]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U21 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U19 ( .A(Fresh[76]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U17 ( .A(Fresh[75]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U16 ( .A1(new_AGEMA_signal_1891), 
        .A2(Ciphertext_s2[50]), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U15 ( .A1(new_AGEMA_signal_1890), 
        .A2(Ciphertext_s1[50]), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_12_Q4), .A2(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_n33), .Z(new_AGEMA_signal_2007) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n32), .B(
        SubCellInst_SboxInst_12_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_n30), .Z(new_AGEMA_signal_2006) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n29), .B(
        SubCellInst_SboxInst_12_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_n27), .Z(SubCellInst_SboxInst_12_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n26), .B(
        SubCellInst_SboxInst_12_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L1), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_Q7) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2008), 
        .B(new_AGEMA_signal_2006), .Z(new_AGEMA_signal_2126) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2009), 
        .B(new_AGEMA_signal_2007), .Z(new_AGEMA_signal_2127) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_XX_2_), .B(SubCellInst_SboxInst_12_T0), .Z(
        SubCellInst_SboxInst_12_L3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1318), .B(new_AGEMA_signal_2004), .Z(new_AGEMA_signal_2128) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1319), .B(new_AGEMA_signal_2005), .Z(new_AGEMA_signal_2129) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L3), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2128), .B(new_AGEMA_signal_2006), .Z(new_AGEMA_signal_2332) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2129), .B(new_AGEMA_signal_2007), .Z(new_AGEMA_signal_2333) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_XX_1_), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1314), .B(new_AGEMA_signal_2006), .Z(new_AGEMA_signal_2252) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1315), .B(new_AGEMA_signal_2007), .Z(new_AGEMA_signal_2253) );
  INV_X1 SubCellInst_SboxInst_13_U3_U1 ( .A(SubCellInst_SboxInst_13_YY_1_), 
        .ZN(AddRoundConstantOutput[55]) );
  INV_X1 SubCellInst_SboxInst_13_U2_U1 ( .A(SubCellInst_SboxInst_13_YY_0_), 
        .ZN(AddRoundConstantOutput[54]) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U37 ( .A(new_AGEMA_signal_1900), .B(
        Fresh[80]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U36 ( .A(Fresh[79]), .B(
        SubCellInst_SboxInst_13_Q1), .Z(
        SubCellInst_SboxInst_13_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U35 ( .A(new_AGEMA_signal_1901), .B(
        Fresh[80]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U34 ( .A(Fresh[78]), .B(
        SubCellInst_SboxInst_13_Q1), .Z(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U33 ( .A(Fresh[79]), .B(
        new_AGEMA_signal_1901), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U32 ( .A(new_AGEMA_signal_1900), .B(
        Fresh[78]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U25 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U24 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U23 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U22 ( .A(Fresh[80]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U21 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U19 ( .A(Fresh[79]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U17 ( .A(Fresh[78]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U16 ( .A1(new_AGEMA_signal_1901), 
        .A2(Ciphertext_s2[54]), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U15 ( .A1(new_AGEMA_signal_1900), 
        .A2(Ciphertext_s1[54]), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_13_Q1), .A2(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_n33), .Z(new_AGEMA_signal_2011) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n32), .B(
        SubCellInst_SboxInst_13_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_n30), .Z(new_AGEMA_signal_2010) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n29), .B(
        SubCellInst_SboxInst_13_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_n27), .Z(SubCellInst_SboxInst_13_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n26), .B(
        SubCellInst_SboxInst_13_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_Q0), .B(SubCellInst_SboxInst_13_T0), .Z(
        SubCellInst_SboxInst_13_Q2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1898), 
        .B(new_AGEMA_signal_2010), .Z(new_AGEMA_signal_2132) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1899), 
        .B(new_AGEMA_signal_2011), .Z(new_AGEMA_signal_2133) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U37 ( .A(new_AGEMA_signal_1902), .B(
        Fresh[83]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U36 ( .A(Fresh[82]), .B(
        SubCellInst_SboxInst_13_Q4), .Z(
        SubCellInst_SboxInst_13_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U35 ( .A(new_AGEMA_signal_1903), .B(
        Fresh[83]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U34 ( .A(Fresh[81]), .B(
        SubCellInst_SboxInst_13_Q4), .Z(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U33 ( .A(Fresh[82]), .B(
        new_AGEMA_signal_1903), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U32 ( .A(new_AGEMA_signal_1902), .B(
        Fresh[81]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U25 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U24 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U23 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U22 ( .A(Fresh[83]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U21 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U19 ( .A(Fresh[82]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U17 ( .A(Fresh[81]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U16 ( .A1(new_AGEMA_signal_1903), 
        .A2(Ciphertext_s2[54]), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U15 ( .A1(new_AGEMA_signal_1902), 
        .A2(Ciphertext_s1[54]), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_13_Q4), .A2(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_n33), .Z(new_AGEMA_signal_2013) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n32), .B(
        SubCellInst_SboxInst_13_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_n30), .Z(new_AGEMA_signal_2012) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n29), .B(
        SubCellInst_SboxInst_13_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_n27), .Z(SubCellInst_SboxInst_13_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n26), .B(
        SubCellInst_SboxInst_13_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L1), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_Q7) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2014), 
        .B(new_AGEMA_signal_2012), .Z(new_AGEMA_signal_2134) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2015), 
        .B(new_AGEMA_signal_2013), .Z(new_AGEMA_signal_2135) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_XX_2_), .B(SubCellInst_SboxInst_13_T0), .Z(
        SubCellInst_SboxInst_13_L3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1330), .B(new_AGEMA_signal_2010), .Z(new_AGEMA_signal_2136) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1331), .B(new_AGEMA_signal_2011), .Z(new_AGEMA_signal_2137) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L3), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2136), .B(new_AGEMA_signal_2012), .Z(new_AGEMA_signal_2336) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2137), .B(new_AGEMA_signal_2013), .Z(new_AGEMA_signal_2337) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_XX_1_), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1326), .B(new_AGEMA_signal_2012), .Z(new_AGEMA_signal_2260) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1327), .B(new_AGEMA_signal_2013), .Z(new_AGEMA_signal_2261) );
  INV_X1 SubCellInst_SboxInst_14_U3_U1 ( .A(SubCellInst_SboxInst_14_YY_1_), 
        .ZN(AddRoundConstantOutput[59]) );
  INV_X1 SubCellInst_SboxInst_14_U2_U1 ( .A(SubCellInst_SboxInst_14_YY_0_), 
        .ZN(AddRoundConstantOutput[58]) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U37 ( .A(new_AGEMA_signal_1912), .B(
        Fresh[86]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U36 ( .A(Fresh[85]), .B(
        SubCellInst_SboxInst_14_Q1), .Z(
        SubCellInst_SboxInst_14_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U35 ( .A(new_AGEMA_signal_1913), .B(
        Fresh[86]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U34 ( .A(Fresh[84]), .B(
        SubCellInst_SboxInst_14_Q1), .Z(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U33 ( .A(Fresh[85]), .B(
        new_AGEMA_signal_1913), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U32 ( .A(new_AGEMA_signal_1912), .B(
        Fresh[84]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U25 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U24 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U23 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U22 ( .A(Fresh[86]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U21 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U19 ( .A(Fresh[85]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U17 ( .A(Fresh[84]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U16 ( .A1(new_AGEMA_signal_1913), 
        .A2(Ciphertext_s2[58]), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U15 ( .A1(new_AGEMA_signal_1912), 
        .A2(Ciphertext_s1[58]), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_14_Q1), .A2(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_n33), .Z(new_AGEMA_signal_2017) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n32), .B(
        SubCellInst_SboxInst_14_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_n30), .Z(new_AGEMA_signal_2016) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n29), .B(
        SubCellInst_SboxInst_14_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_n27), .Z(SubCellInst_SboxInst_14_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n26), .B(
        SubCellInst_SboxInst_14_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_Q0), .B(SubCellInst_SboxInst_14_T0), .Z(
        SubCellInst_SboxInst_14_Q2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1910), 
        .B(new_AGEMA_signal_2016), .Z(new_AGEMA_signal_2140) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1911), 
        .B(new_AGEMA_signal_2017), .Z(new_AGEMA_signal_2141) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U37 ( .A(new_AGEMA_signal_1914), .B(
        Fresh[89]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U36 ( .A(Fresh[88]), .B(
        SubCellInst_SboxInst_14_Q4), .Z(
        SubCellInst_SboxInst_14_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U35 ( .A(new_AGEMA_signal_1915), .B(
        Fresh[89]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U34 ( .A(Fresh[87]), .B(
        SubCellInst_SboxInst_14_Q4), .Z(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U33 ( .A(Fresh[88]), .B(
        new_AGEMA_signal_1915), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U32 ( .A(new_AGEMA_signal_1914), .B(
        Fresh[87]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U25 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U24 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U23 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U22 ( .A(Fresh[89]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U21 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U19 ( .A(Fresh[88]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U17 ( .A(Fresh[87]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U16 ( .A1(new_AGEMA_signal_1915), 
        .A2(Ciphertext_s2[58]), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U15 ( .A1(new_AGEMA_signal_1914), 
        .A2(Ciphertext_s1[58]), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_14_Q4), .A2(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_n33), .Z(new_AGEMA_signal_2019) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n32), .B(
        SubCellInst_SboxInst_14_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_n30), .Z(new_AGEMA_signal_2018) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n29), .B(
        SubCellInst_SboxInst_14_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_n27), .Z(SubCellInst_SboxInst_14_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n26), .B(
        SubCellInst_SboxInst_14_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L1), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_Q7) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2020), 
        .B(new_AGEMA_signal_2018), .Z(new_AGEMA_signal_2142) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2021), 
        .B(new_AGEMA_signal_2019), .Z(new_AGEMA_signal_2143) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_XX_2_), .B(SubCellInst_SboxInst_14_T0), .Z(
        SubCellInst_SboxInst_14_L3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1342), .B(new_AGEMA_signal_2016), .Z(new_AGEMA_signal_2144) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1343), .B(new_AGEMA_signal_2017), .Z(new_AGEMA_signal_2145) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L3), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2144), .B(new_AGEMA_signal_2018), .Z(new_AGEMA_signal_2340) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2145), .B(new_AGEMA_signal_2019), .Z(new_AGEMA_signal_2341) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_XX_1_), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1338), .B(new_AGEMA_signal_2018), .Z(new_AGEMA_signal_2268) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1339), .B(new_AGEMA_signal_2019), .Z(new_AGEMA_signal_2269) );
  INV_X1 SubCellInst_SboxInst_15_U3_U1 ( .A(SubCellInst_SboxInst_15_YY_1_), 
        .ZN(SubCellOutput[63]) );
  INV_X1 SubCellInst_SboxInst_15_U2_U1 ( .A(SubCellInst_SboxInst_15_YY_0_), 
        .ZN(SubCellOutput[62]) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U37 ( .A(new_AGEMA_signal_1924), .B(
        Fresh[92]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U36 ( .A(Fresh[91]), .B(
        SubCellInst_SboxInst_15_Q1), .Z(
        SubCellInst_SboxInst_15_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U35 ( .A(new_AGEMA_signal_1925), .B(
        Fresh[92]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U34 ( .A(Fresh[90]), .B(
        SubCellInst_SboxInst_15_Q1), .Z(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U33 ( .A(Fresh[91]), .B(
        new_AGEMA_signal_1925), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U32 ( .A(new_AGEMA_signal_1924), .B(
        Fresh[90]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U25 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U24 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U23 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U22 ( .A(Fresh[92]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U21 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U19 ( .A(Fresh[91]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U17 ( .A(Fresh[90]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U16 ( .A1(new_AGEMA_signal_1925), 
        .A2(Ciphertext_s2[62]), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U15 ( .A1(new_AGEMA_signal_1924), 
        .A2(Ciphertext_s1[62]), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_15_Q1), .A2(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_n33), .Z(new_AGEMA_signal_2023) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n32), .B(
        SubCellInst_SboxInst_15_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_n30), .Z(new_AGEMA_signal_2022) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n29), .B(
        SubCellInst_SboxInst_15_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_n27), .Z(SubCellInst_SboxInst_15_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n26), .B(
        SubCellInst_SboxInst_15_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_Q0), .B(SubCellInst_SboxInst_15_T0), .Z(
        SubCellInst_SboxInst_15_Q2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1922), 
        .B(new_AGEMA_signal_2022), .Z(new_AGEMA_signal_2148) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1923), 
        .B(new_AGEMA_signal_2023), .Z(new_AGEMA_signal_2149) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U37 ( .A(new_AGEMA_signal_1926), .B(
        Fresh[95]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U36 ( .A(Fresh[94]), .B(
        SubCellInst_SboxInst_15_Q4), .Z(
        SubCellInst_SboxInst_15_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U35 ( .A(new_AGEMA_signal_1927), .B(
        Fresh[95]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U34 ( .A(Fresh[93]), .B(
        SubCellInst_SboxInst_15_Q4), .Z(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U33 ( .A(Fresh[94]), .B(
        new_AGEMA_signal_1927), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U32 ( .A(new_AGEMA_signal_1926), .B(
        Fresh[93]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U25 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U24 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U23 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U22 ( .A(Fresh[95]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U21 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U19 ( .A(Fresh[94]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U17 ( .A(Fresh[93]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U16 ( .A1(new_AGEMA_signal_1927), 
        .A2(Ciphertext_s2[62]), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U15 ( .A1(new_AGEMA_signal_1926), 
        .A2(Ciphertext_s1[62]), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_15_Q4), .A2(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_n33), .Z(new_AGEMA_signal_2025) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n32), .B(
        SubCellInst_SboxInst_15_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_n30), .Z(new_AGEMA_signal_2024) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n29), .B(
        SubCellInst_SboxInst_15_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_n27), .Z(SubCellInst_SboxInst_15_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n26), .B(
        SubCellInst_SboxInst_15_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L1), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_Q7) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2026), 
        .B(new_AGEMA_signal_2024), .Z(new_AGEMA_signal_2150) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2027), 
        .B(new_AGEMA_signal_2025), .Z(new_AGEMA_signal_2151) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_XX_2_), .B(SubCellInst_SboxInst_15_T0), .Z(
        SubCellInst_SboxInst_15_L3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1354), .B(new_AGEMA_signal_2022), .Z(new_AGEMA_signal_2152) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1355), .B(new_AGEMA_signal_2023), .Z(new_AGEMA_signal_2153) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L3), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2152), .B(new_AGEMA_signal_2024), .Z(new_AGEMA_signal_2344) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2153), .B(new_AGEMA_signal_2025), .Z(new_AGEMA_signal_2345) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_XX_1_), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1350), .B(new_AGEMA_signal_2024), .Z(new_AGEMA_signal_2276) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1351), .B(new_AGEMA_signal_2025), .Z(new_AGEMA_signal_2277) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_2_n1), .B(FSMUpdate[3]), .ZN(
        AddRoundConstantOutput[62]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2348), .B(1'b0), .Z(new_AGEMA_signal_2436) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2349), .B(1'b0), .Z(new_AGEMA_signal_2437) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[62]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_2_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2276), .Z(new_AGEMA_signal_2348) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2277), .Z(new_AGEMA_signal_2349) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_3_n1), .B(FSMUpdate[4]), .ZN(
        AddRoundConstantOutput[63]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2438), .B(1'b0), .Z(new_AGEMA_signal_2522) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2439), .B(1'b0), .Z(new_AGEMA_signal_2523) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[63]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_3_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2344), .Z(new_AGEMA_signal_2438) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2345), .Z(new_AGEMA_signal_2439) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_2_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[46]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2350), .B(1'b0), .Z(new_AGEMA_signal_2440) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2351), .B(1'b0), .Z(new_AGEMA_signal_2441) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_46), .ZN(AddConstXOR_AddConstXOR_XORInst_1_2_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2244), .Z(new_AGEMA_signal_2350) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2245), .Z(new_AGEMA_signal_2351) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_3_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[47]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2442), .B(1'b0), .Z(new_AGEMA_signal_2526) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2443), .B(1'b0), .Z(new_AGEMA_signal_2527) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_47), .ZN(AddConstXOR_AddConstXOR_XORInst_1_3_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2328), .Z(new_AGEMA_signal_2442) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2329), .Z(new_AGEMA_signal_2443) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_2_n1), .B(
        TweakeyGeneration_key_Feedback[2]), .ZN(ShiftRowsOutput[46]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2352), .B(new_AGEMA_signal_1368), .Z(
        new_AGEMA_signal_2444) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2353), .B(new_AGEMA_signal_1369), .Z(
        new_AGEMA_signal_2445) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[34]), .ZN(AddRoundTweakeyXOR_XORInst_0_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2220), .Z(new_AGEMA_signal_2352) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2221), .Z(new_AGEMA_signal_2353) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_3_n1), .B(
        TweakeyGeneration_key_Feedback[3]), .ZN(ShiftRowsOutput[47]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2446), .B(new_AGEMA_signal_1374), .Z(
        new_AGEMA_signal_2530) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2447), .B(new_AGEMA_signal_1375), .Z(
        new_AGEMA_signal_2531) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[35]), .ZN(AddRoundTweakeyXOR_XORInst_0_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2316), .Z(new_AGEMA_signal_2446) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2317), .Z(new_AGEMA_signal_2447) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_2_n1), .B(
        TweakeyGeneration_key_Feedback[6]), .ZN(ShiftRowsOutput[34]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2354), .B(new_AGEMA_signal_1392), .Z(
        new_AGEMA_signal_2448) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2355), .B(new_AGEMA_signal_1393), .Z(
        new_AGEMA_signal_2449) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[38]), .ZN(AddRoundTweakeyXOR_XORInst_1_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2228), .Z(new_AGEMA_signal_2354) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2229), .Z(new_AGEMA_signal_2355) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_3_n1), .B(
        TweakeyGeneration_key_Feedback[7]), .ZN(ShiftRowsOutput[35]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2450), .B(new_AGEMA_signal_1398), .Z(
        new_AGEMA_signal_2534) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2451), .B(new_AGEMA_signal_1399), .Z(
        new_AGEMA_signal_2535) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[39]), .ZN(AddRoundTweakeyXOR_XORInst_1_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2320), .Z(new_AGEMA_signal_2450) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2321), .Z(new_AGEMA_signal_2451) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_2_n1), .B(
        TweakeyGeneration_key_Feedback[10]), .ZN(ShiftRowsOutput[38]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2356), .B(new_AGEMA_signal_1416), .Z(
        new_AGEMA_signal_2452) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2357), .B(new_AGEMA_signal_1417), .Z(
        new_AGEMA_signal_2453) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[42]), .ZN(AddRoundTweakeyXOR_XORInst_2_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2236), .Z(new_AGEMA_signal_2356) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2237), .Z(new_AGEMA_signal_2357) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_3_n1), .B(
        TweakeyGeneration_key_Feedback[11]), .ZN(ShiftRowsOutput[39]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2454), .B(new_AGEMA_signal_1422), .Z(
        new_AGEMA_signal_2538) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2455), .B(new_AGEMA_signal_1423), .Z(
        new_AGEMA_signal_2539) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[43]), .ZN(AddRoundTweakeyXOR_XORInst_2_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2324), .Z(new_AGEMA_signal_2454) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2325), .Z(new_AGEMA_signal_2455) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_2_n1), .B(
        TweakeyGeneration_key_Feedback[14]), .ZN(ShiftRowsOutput[42]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2540), .B(new_AGEMA_signal_1440), .Z(
        new_AGEMA_signal_2616) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2541), .B(new_AGEMA_signal_1441), .Z(
        new_AGEMA_signal_2617) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[46]), .ZN(AddRoundTweakeyXOR_XORInst_3_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2440), .Z(new_AGEMA_signal_2540) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2441), .Z(new_AGEMA_signal_2541) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_3_n1), .B(
        TweakeyGeneration_key_Feedback[15]), .ZN(ShiftRowsOutput[43]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2618), .B(new_AGEMA_signal_1446), .Z(
        new_AGEMA_signal_2742) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2619), .B(new_AGEMA_signal_1447), .Z(
        new_AGEMA_signal_2743) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[47]), .ZN(AddRoundTweakeyXOR_XORInst_3_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2526), .Z(new_AGEMA_signal_2618) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2527), .Z(new_AGEMA_signal_2619) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_2_n1), .B(
        TweakeyGeneration_key_Feedback[18]), .ZN(MCOutput[34]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2358), .B(new_AGEMA_signal_1464), .Z(
        new_AGEMA_signal_2456) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2359), .B(new_AGEMA_signal_1465), .Z(
        new_AGEMA_signal_2457) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[50]), .ZN(AddRoundTweakeyXOR_XORInst_4_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2252), .Z(new_AGEMA_signal_2358) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2253), .Z(new_AGEMA_signal_2359) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_3_n1), .B(
        TweakeyGeneration_key_Feedback[19]), .ZN(MCOutput[35]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2458), .B(new_AGEMA_signal_1470), .Z(
        new_AGEMA_signal_2544) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2459), .B(new_AGEMA_signal_1471), .Z(
        new_AGEMA_signal_2545) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[51]), .ZN(AddRoundTweakeyXOR_XORInst_4_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2332), .Z(new_AGEMA_signal_2458) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2333), .Z(new_AGEMA_signal_2459) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_2_n1), .B(
        TweakeyGeneration_key_Feedback[22]), .ZN(MCOutput[38]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2360), .B(new_AGEMA_signal_1488), .Z(
        new_AGEMA_signal_2460) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2361), .B(new_AGEMA_signal_1489), .Z(
        new_AGEMA_signal_2461) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[54]), .ZN(AddRoundTweakeyXOR_XORInst_5_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2260), .Z(new_AGEMA_signal_2360) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2261), .Z(new_AGEMA_signal_2361) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_3_n1), .B(
        TweakeyGeneration_key_Feedback[23]), .ZN(MCOutput[39]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2462), .B(new_AGEMA_signal_1494), .Z(
        new_AGEMA_signal_2548) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2463), .B(new_AGEMA_signal_1495), .Z(
        new_AGEMA_signal_2549) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[55]), .ZN(AddRoundTweakeyXOR_XORInst_5_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2336), .Z(new_AGEMA_signal_2462) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2337), .Z(new_AGEMA_signal_2463) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_2_n1), .B(
        TweakeyGeneration_key_Feedback[26]), .ZN(MCOutput[42]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2362), .B(new_AGEMA_signal_1512), .Z(
        new_AGEMA_signal_2464) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2363), .B(new_AGEMA_signal_1513), .Z(
        new_AGEMA_signal_2465) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[58]), .ZN(AddRoundTweakeyXOR_XORInst_6_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2268), .Z(new_AGEMA_signal_2362) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2269), .Z(new_AGEMA_signal_2363) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_3_n1), .B(
        TweakeyGeneration_key_Feedback[27]), .ZN(MCOutput[43]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2466), .B(new_AGEMA_signal_1518), .Z(
        new_AGEMA_signal_2552) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2467), .B(new_AGEMA_signal_1519), .Z(
        new_AGEMA_signal_2553) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[59]), .ZN(AddRoundTweakeyXOR_XORInst_6_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2340), .Z(new_AGEMA_signal_2466) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2341), .Z(new_AGEMA_signal_2467) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_2_n1), .B(
        TweakeyGeneration_key_Feedback[30]), .ZN(MCOutput[46]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2554), .B(new_AGEMA_signal_1536), .Z(
        new_AGEMA_signal_2632) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2555), .B(new_AGEMA_signal_1537), .Z(
        new_AGEMA_signal_2633) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[62]), .ZN(AddRoundTweakeyXOR_XORInst_7_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2436), .Z(new_AGEMA_signal_2554) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2437), .Z(new_AGEMA_signal_2555) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_3_n1), .B(
        TweakeyGeneration_key_Feedback[31]), .ZN(MCOutput[47]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2634), .B(new_AGEMA_signal_1542), .Z(
        new_AGEMA_signal_2752) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2635), .B(new_AGEMA_signal_1543), .Z(
        new_AGEMA_signal_2753) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[63]), .ZN(AddRoundTweakeyXOR_XORInst_7_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2522), .Z(new_AGEMA_signal_2634) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2523), .Z(new_AGEMA_signal_2635) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_2_n2), 
        .B(MCInst_MCR0_XORInst_0_2_n1), .ZN(MCOutput[50]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2558), .B(
        new_AGEMA_signal_2364), .Z(new_AGEMA_signal_2638) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2559), .B(
        new_AGEMA_signal_2365), .Z(new_AGEMA_signal_2639) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[18]), .B(
        ShiftRowsOutput[2]), .ZN(MCInst_MCR0_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2204), .B(
        new_AGEMA_signal_2180), .Z(new_AGEMA_signal_2364) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2205), .B(
        new_AGEMA_signal_2181), .Z(new_AGEMA_signal_2365) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[34]), 
        .Z(MCInst_MCR0_XORInst_0_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2456), .Z(new_AGEMA_signal_2558) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2457), .Z(new_AGEMA_signal_2559) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_3_n2), 
        .B(MCInst_MCR0_XORInst_0_3_n1), .ZN(MCOutput[51]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2640), .B(
        new_AGEMA_signal_2468), .Z(new_AGEMA_signal_2756) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2641), .B(
        new_AGEMA_signal_2469), .Z(new_AGEMA_signal_2757) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[19]), .B(
        ShiftRowsOutput[3]), .ZN(MCInst_MCR0_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2308), .B(
        new_AGEMA_signal_2296), .Z(new_AGEMA_signal_2468) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2309), .B(
        new_AGEMA_signal_2297), .Z(new_AGEMA_signal_2469) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[35]), 
        .Z(MCInst_MCR0_XORInst_0_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2544), .Z(new_AGEMA_signal_2640) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2545), .Z(new_AGEMA_signal_2641) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_2_n2), 
        .B(MCInst_MCR0_XORInst_1_2_n1), .ZN(MCOutput[54]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2562), .B(
        new_AGEMA_signal_2366), .Z(new_AGEMA_signal_2642) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2563), .B(
        new_AGEMA_signal_2367), .Z(new_AGEMA_signal_2643) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[22]), .B(
        ShiftRowsOutput[6]), .ZN(MCInst_MCR0_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2212), .B(
        new_AGEMA_signal_2156), .Z(new_AGEMA_signal_2366) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2213), .B(
        new_AGEMA_signal_2157), .Z(new_AGEMA_signal_2367) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[38]), 
        .Z(MCInst_MCR0_XORInst_1_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2460), .Z(new_AGEMA_signal_2562) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2461), .Z(new_AGEMA_signal_2563) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_3_n2), 
        .B(MCInst_MCR0_XORInst_1_3_n1), .ZN(MCOutput[55]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2644), .B(
        new_AGEMA_signal_2470), .Z(new_AGEMA_signal_2762) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2645), .B(
        new_AGEMA_signal_2471), .Z(new_AGEMA_signal_2763) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[23]), .B(
        ShiftRowsOutput[7]), .ZN(MCInst_MCR0_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2312), .B(
        new_AGEMA_signal_2284), .Z(new_AGEMA_signal_2470) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2313), .B(
        new_AGEMA_signal_2285), .Z(new_AGEMA_signal_2471) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[39]), 
        .Z(MCInst_MCR0_XORInst_1_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2548), .Z(new_AGEMA_signal_2644) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2549), .Z(new_AGEMA_signal_2645) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_2_n2), 
        .B(MCInst_MCR0_XORInst_2_2_n1), .ZN(MCOutput[58]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2566), .B(
        new_AGEMA_signal_2368), .Z(new_AGEMA_signal_2648) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2567), .B(
        new_AGEMA_signal_2369), .Z(new_AGEMA_signal_2649) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[26]), .B(
        ShiftRowsOutput[10]), .ZN(MCInst_MCR0_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2188), .B(
        new_AGEMA_signal_2164), .Z(new_AGEMA_signal_2368) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2189), .B(
        new_AGEMA_signal_2165), .Z(new_AGEMA_signal_2369) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[42]), 
        .Z(MCInst_MCR0_XORInst_2_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2464), .Z(new_AGEMA_signal_2566) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2465), .Z(new_AGEMA_signal_2567) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_3_n2), 
        .B(MCInst_MCR0_XORInst_2_3_n1), .ZN(MCOutput[59]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2650), .B(
        new_AGEMA_signal_2472), .Z(new_AGEMA_signal_2766) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2651), .B(
        new_AGEMA_signal_2473), .Z(new_AGEMA_signal_2767) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[27]), .B(
        ShiftRowsOutput[11]), .ZN(MCInst_MCR0_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2300), .B(
        new_AGEMA_signal_2288), .Z(new_AGEMA_signal_2472) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2301), .B(
        new_AGEMA_signal_2289), .Z(new_AGEMA_signal_2473) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[43]), 
        .Z(MCInst_MCR0_XORInst_2_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2552), .Z(new_AGEMA_signal_2650) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2553), .Z(new_AGEMA_signal_2651) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_2_n2), 
        .B(MCInst_MCR0_XORInst_3_2_n1), .ZN(MCOutput[62]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2768), .B(
        new_AGEMA_signal_2370), .Z(new_AGEMA_signal_2870) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2769), .B(
        new_AGEMA_signal_2371), .Z(new_AGEMA_signal_2871) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[30]), .B(
        ShiftRowsOutput[14]), .ZN(MCInst_MCR0_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2196), .B(
        new_AGEMA_signal_2172), .Z(new_AGEMA_signal_2370) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2197), .B(
        new_AGEMA_signal_2173), .Z(new_AGEMA_signal_2371) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[46]), 
        .Z(MCInst_MCR0_XORInst_3_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2632), .Z(new_AGEMA_signal_2768) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2633), .Z(new_AGEMA_signal_2769) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_3_n2), 
        .B(MCInst_MCR0_XORInst_3_3_n1), .ZN(MCOutput[63]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2872), .B(
        new_AGEMA_signal_2474), .Z(new_AGEMA_signal_2970) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2873), .B(
        new_AGEMA_signal_2475), .Z(new_AGEMA_signal_2971) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[31]), .B(
        ShiftRowsOutput[15]), .ZN(MCInst_MCR0_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2304), .B(
        new_AGEMA_signal_2292), .Z(new_AGEMA_signal_2474) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2305), .B(
        new_AGEMA_signal_2293), .Z(new_AGEMA_signal_2475) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[47]), 
        .Z(MCInst_MCR0_XORInst_3_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2752), .Z(new_AGEMA_signal_2872) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2753), .Z(new_AGEMA_signal_2873) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_2_n1), 
        .B(ShiftRowsOutput[18]), .ZN(MCOutput[18]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2570), .B(
        new_AGEMA_signal_2204), .Z(new_AGEMA_signal_2654) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2571), .B(
        new_AGEMA_signal_2205), .Z(new_AGEMA_signal_2655) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[34]), .ZN(MCInst_MCR2_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2448), .Z(new_AGEMA_signal_2570) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2449), .Z(new_AGEMA_signal_2571) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_3_n1), 
        .B(ShiftRowsOutput[19]), .ZN(MCOutput[19]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2656), .B(
        new_AGEMA_signal_2308), .Z(new_AGEMA_signal_2772) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2657), .B(
        new_AGEMA_signal_2309), .Z(new_AGEMA_signal_2773) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[35]), .ZN(MCInst_MCR2_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2534), .Z(new_AGEMA_signal_2656) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2535), .Z(new_AGEMA_signal_2657) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_2_n1), 
        .B(ShiftRowsOutput[22]), .ZN(MCOutput[22]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2572), .B(
        new_AGEMA_signal_2212), .Z(new_AGEMA_signal_2658) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2573), .B(
        new_AGEMA_signal_2213), .Z(new_AGEMA_signal_2659) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[38]), .ZN(MCInst_MCR2_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2452), .Z(new_AGEMA_signal_2572) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2453), .Z(new_AGEMA_signal_2573) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_3_n1), 
        .B(ShiftRowsOutput[23]), .ZN(MCOutput[23]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2660), .B(
        new_AGEMA_signal_2312), .Z(new_AGEMA_signal_2776) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2661), .B(
        new_AGEMA_signal_2313), .Z(new_AGEMA_signal_2777) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[39]), .ZN(MCInst_MCR2_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2538), .Z(new_AGEMA_signal_2660) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2539), .Z(new_AGEMA_signal_2661) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_2_n1), 
        .B(ShiftRowsOutput[26]), .ZN(MCOutput[26]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2778), .B(
        new_AGEMA_signal_2188), .Z(new_AGEMA_signal_2882) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2779), .B(
        new_AGEMA_signal_2189), .Z(new_AGEMA_signal_2883) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[42]), .ZN(MCInst_MCR2_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2616), .Z(new_AGEMA_signal_2778) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2617), .Z(new_AGEMA_signal_2779) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_3_n1), 
        .B(ShiftRowsOutput[27]), .ZN(MCOutput[27]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2884), .B(
        new_AGEMA_signal_2300), .Z(new_AGEMA_signal_2978) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2885), .B(
        new_AGEMA_signal_2301), .Z(new_AGEMA_signal_2979) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[43]), .ZN(MCInst_MCR2_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2742), .Z(new_AGEMA_signal_2884) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2743), .Z(new_AGEMA_signal_2885) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_2_n1), 
        .B(ShiftRowsOutput[30]), .ZN(MCOutput[30]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2574), .B(
        new_AGEMA_signal_2196), .Z(new_AGEMA_signal_2662) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2575), .B(
        new_AGEMA_signal_2197), .Z(new_AGEMA_signal_2663) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[46]), .ZN(MCInst_MCR2_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2444), .Z(new_AGEMA_signal_2574) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2445), .Z(new_AGEMA_signal_2575) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_3_n1), 
        .B(ShiftRowsOutput[31]), .ZN(MCOutput[31]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2664), .B(
        new_AGEMA_signal_2304), .Z(new_AGEMA_signal_2782) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2665), .B(
        new_AGEMA_signal_2305), .Z(new_AGEMA_signal_2783) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[47]), .ZN(MCInst_MCR2_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2530), .Z(new_AGEMA_signal_2664) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2531), .Z(new_AGEMA_signal_2665) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_2_n1), 
        .B(ShiftRowsOutput[18]), .ZN(MCOutput[2]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2576), .B(
        new_AGEMA_signal_2204), .Z(new_AGEMA_signal_2666) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2577), .B(
        new_AGEMA_signal_2205), .Z(new_AGEMA_signal_2667) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[34]), 
        .ZN(MCInst_MCR3_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2456), .Z(new_AGEMA_signal_2576) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2457), .Z(new_AGEMA_signal_2577) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_3_n1), 
        .B(ShiftRowsOutput[19]), .ZN(MCOutput[3]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2668), .B(
        new_AGEMA_signal_2308), .Z(new_AGEMA_signal_2786) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2669), .B(
        new_AGEMA_signal_2309), .Z(new_AGEMA_signal_2787) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[35]), 
        .ZN(MCInst_MCR3_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2544), .Z(new_AGEMA_signal_2668) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2545), .Z(new_AGEMA_signal_2669) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_2_n1), 
        .B(ShiftRowsOutput[22]), .ZN(MCOutput[6]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2578), .B(
        new_AGEMA_signal_2212), .Z(new_AGEMA_signal_2670) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2579), .B(
        new_AGEMA_signal_2213), .Z(new_AGEMA_signal_2671) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[38]), 
        .ZN(MCInst_MCR3_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2460), .Z(new_AGEMA_signal_2578) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2461), .Z(new_AGEMA_signal_2579) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_3_n1), 
        .B(ShiftRowsOutput[23]), .ZN(MCOutput[7]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2672), .B(
        new_AGEMA_signal_2312), .Z(new_AGEMA_signal_2790) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2673), .B(
        new_AGEMA_signal_2313), .Z(new_AGEMA_signal_2791) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[39]), 
        .ZN(MCInst_MCR3_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2548), .Z(new_AGEMA_signal_2672) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2549), .Z(new_AGEMA_signal_2673) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_2_n1), 
        .B(ShiftRowsOutput[26]), .ZN(MCOutput[10]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2580), .B(
        new_AGEMA_signal_2188), .Z(new_AGEMA_signal_2674) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2581), .B(
        new_AGEMA_signal_2189), .Z(new_AGEMA_signal_2675) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[42]), 
        .ZN(MCInst_MCR3_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2464), .Z(new_AGEMA_signal_2580) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2465), .Z(new_AGEMA_signal_2581) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_3_n1), 
        .B(ShiftRowsOutput[27]), .ZN(MCOutput[11]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2676), .B(
        new_AGEMA_signal_2300), .Z(new_AGEMA_signal_2794) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2677), .B(
        new_AGEMA_signal_2301), .Z(new_AGEMA_signal_2795) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[43]), 
        .ZN(MCInst_MCR3_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2552), .Z(new_AGEMA_signal_2676) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2553), .Z(new_AGEMA_signal_2677) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_2_n1), 
        .B(ShiftRowsOutput[30]), .ZN(MCOutput[14]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2796), .B(
        new_AGEMA_signal_2196), .Z(new_AGEMA_signal_2902) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2797), .B(
        new_AGEMA_signal_2197), .Z(new_AGEMA_signal_2903) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[46]), 
        .ZN(MCInst_MCR3_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2632), .Z(new_AGEMA_signal_2796) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2633), .Z(new_AGEMA_signal_2797) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_3_n1), 
        .B(ShiftRowsOutput[31]), .ZN(MCOutput[15]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2904), .B(
        new_AGEMA_signal_2304), .Z(new_AGEMA_signal_2990) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2905), .B(
        new_AGEMA_signal_2305), .Z(new_AGEMA_signal_2991) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[47]), 
        .ZN(MCInst_MCR3_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2752), .Z(new_AGEMA_signal_2904) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2753), .Z(new_AGEMA_signal_2905) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_0_U1 ( .A(MCOutput[0]), .B(
        Plaintext_s0[0]), .S(rst), .Z(StateRegInput[0]) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2890), .B(
        Plaintext_s1[0]), .S(rst), .Z(new_AGEMA_signal_2908) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2891), .B(
        Plaintext_s2[0]), .S(rst), .Z(new_AGEMA_signal_2909) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_0_U1 ( .A(MCOutput[1]), .B(
        Plaintext_s0[1]), .S(rst), .Z(StateRegInput[1]) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2982), .B(
        Plaintext_s1[1]), .S(rst), .Z(new_AGEMA_signal_2994) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2983), .B(
        Plaintext_s2[1]), .S(rst), .Z(new_AGEMA_signal_2995) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_0_U1 ( .A(MCOutput[4]), .B(
        Plaintext_s0[4]), .S(rst), .Z(StateRegInput[4]) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2894), .B(
        Plaintext_s1[4]), .S(rst), .Z(new_AGEMA_signal_2912) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2895), .B(
        Plaintext_s2[4]), .S(rst), .Z(new_AGEMA_signal_2913) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_0_U1 ( .A(MCOutput[5]), .B(
        Plaintext_s0[5]), .S(rst), .Z(StateRegInput[5]) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2984), .B(
        Plaintext_s1[5]), .S(rst), .Z(new_AGEMA_signal_2998) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2985), .B(
        Plaintext_s2[5]), .S(rst), .Z(new_AGEMA_signal_2999) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_0_U1 ( .A(MCOutput[8]), .B(
        Plaintext_s0[8]), .S(rst), .Z(StateRegInput[8]) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2898), .B(
        Plaintext_s1[8]), .S(rst), .Z(new_AGEMA_signal_2916) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2899), .B(
        Plaintext_s2[8]), .S(rst), .Z(new_AGEMA_signal_2917) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_0_U1 ( .A(MCOutput[9]), .B(
        Plaintext_s0[9]), .S(rst), .Z(StateRegInput[9]) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2986), .B(
        Plaintext_s1[9]), .S(rst), .Z(new_AGEMA_signal_3002) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2987), .B(
        Plaintext_s2[9]), .S(rst), .Z(new_AGEMA_signal_3003) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_0_U1 ( .A(MCOutput[12]), .B(
        Plaintext_s0[12]), .S(rst), .Z(StateRegInput[12]) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3052), .B(
        Plaintext_s1[12]), .S(rst), .Z(new_AGEMA_signal_3058) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3053), .B(
        Plaintext_s2[12]), .S(rst), .Z(new_AGEMA_signal_3059) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_0_U1 ( .A(MCOutput[13]), .B(
        Plaintext_s0[13]), .S(rst), .Z(StateRegInput[13]) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3072), .B(
        Plaintext_s1[13]), .S(rst), .Z(new_AGEMA_signal_3076) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3073), .B(
        Plaintext_s2[13]), .S(rst), .Z(new_AGEMA_signal_3077) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_0_U1 ( .A(MCOutput[16]), .B(
        Plaintext_s0[16]), .S(rst), .Z(StateRegInput[16]) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2874), .B(
        Plaintext_s1[16]), .S(rst), .Z(new_AGEMA_signal_2924) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2875), .B(
        Plaintext_s2[16]), .S(rst), .Z(new_AGEMA_signal_2925) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_0_U1 ( .A(MCOutput[17]), .B(
        Plaintext_s0[17]), .S(rst), .Z(StateRegInput[17]) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2972), .B(
        Plaintext_s1[17]), .S(rst), .Z(new_AGEMA_signal_3010) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2973), .B(
        Plaintext_s2[17]), .S(rst), .Z(new_AGEMA_signal_3011) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_0_U1 ( .A(MCOutput[20]), .B(
        Plaintext_s0[20]), .S(rst), .Z(StateRegInput[20]) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2878), .B(
        Plaintext_s1[20]), .S(rst), .Z(new_AGEMA_signal_2928) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2879), .B(
        Plaintext_s2[20]), .S(rst), .Z(new_AGEMA_signal_2929) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_0_U1 ( .A(MCOutput[21]), .B(
        Plaintext_s0[21]), .S(rst), .Z(StateRegInput[21]) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2974), .B(
        Plaintext_s1[21]), .S(rst), .Z(new_AGEMA_signal_3014) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2975), .B(
        Plaintext_s2[21]), .S(rst), .Z(new_AGEMA_signal_3015) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_0_U1 ( .A(MCOutput[24]), .B(
        Plaintext_s0[24]), .S(rst), .Z(StateRegInput[24]) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3048), .B(
        Plaintext_s1[24]), .S(rst), .Z(new_AGEMA_signal_3062) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3049), .B(
        Plaintext_s2[24]), .S(rst), .Z(new_AGEMA_signal_3063) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_0_U1 ( .A(MCOutput[25]), .B(
        Plaintext_s0[25]), .S(rst), .Z(StateRegInput[25]) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3070), .B(
        Plaintext_s1[25]), .S(rst), .Z(new_AGEMA_signal_3080) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3071), .B(
        Plaintext_s2[25]), .S(rst), .Z(new_AGEMA_signal_3081) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_0_U1 ( .A(MCOutput[28]), .B(
        Plaintext_s0[28]), .S(rst), .Z(StateRegInput[28]) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2886), .B(
        Plaintext_s1[28]), .S(rst), .Z(new_AGEMA_signal_2936) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2887), .B(
        Plaintext_s2[28]), .S(rst), .Z(new_AGEMA_signal_2937) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_0_U1 ( .A(MCOutput[29]), .B(
        Plaintext_s0[29]), .S(rst), .Z(StateRegInput[29]) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2980), .B(
        Plaintext_s1[29]), .S(rst), .Z(new_AGEMA_signal_3022) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2981), .B(
        Plaintext_s2[29]), .S(rst), .Z(new_AGEMA_signal_3023) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_0_U1 ( .A(MCOutput[32]), .B(
        Plaintext_s0[32]), .S(rst), .Z(StateRegInput[32]) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2620), .B(
        Plaintext_s1[32]), .S(rst), .Z(new_AGEMA_signal_2704) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2621), .B(
        Plaintext_s2[32]), .S(rst), .Z(new_AGEMA_signal_2705) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_0_U1 ( .A(MCOutput[33]), .B(
        Plaintext_s0[33]), .S(rst), .Z(StateRegInput[33]) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2744), .B(
        Plaintext_s1[33]), .S(rst), .Z(new_AGEMA_signal_2824) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2745), .B(
        Plaintext_s2[33]), .S(rst), .Z(new_AGEMA_signal_2825) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_0_U1 ( .A(MCOutput[36]), .B(
        Plaintext_s0[36]), .S(rst), .Z(StateRegInput[36]) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2624), .B(
        Plaintext_s1[36]), .S(rst), .Z(new_AGEMA_signal_2708) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2625), .B(
        Plaintext_s2[36]), .S(rst), .Z(new_AGEMA_signal_2709) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_0_U1 ( .A(MCOutput[37]), .B(
        Plaintext_s0[37]), .S(rst), .Z(StateRegInput[37]) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2746), .B(
        Plaintext_s1[37]), .S(rst), .Z(new_AGEMA_signal_2828) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2747), .B(
        Plaintext_s2[37]), .S(rst), .Z(new_AGEMA_signal_2829) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_0_U1 ( .A(MCOutput[40]), .B(
        Plaintext_s0[40]), .S(rst), .Z(StateRegInput[40]) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2628), .B(
        Plaintext_s1[40]), .S(rst), .Z(new_AGEMA_signal_2712) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2629), .B(
        Plaintext_s2[40]), .S(rst), .Z(new_AGEMA_signal_2713) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_0_U1 ( .A(MCOutput[41]), .B(
        Plaintext_s0[41]), .S(rst), .Z(StateRegInput[41]) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2748), .B(
        Plaintext_s1[41]), .S(rst), .Z(new_AGEMA_signal_2832) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2749), .B(
        Plaintext_s2[41]), .S(rst), .Z(new_AGEMA_signal_2833) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_0_U1 ( .A(MCOutput[44]), .B(
        Plaintext_s0[44]), .S(rst), .Z(StateRegInput[44]) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2854), .B(
        Plaintext_s1[44]), .S(rst), .Z(new_AGEMA_signal_2940) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2855), .B(
        Plaintext_s2[44]), .S(rst), .Z(new_AGEMA_signal_2941) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_0_U1 ( .A(MCOutput[45]), .B(
        Plaintext_s0[45]), .S(rst), .Z(StateRegInput[45]) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2960), .B(
        Plaintext_s1[45]), .S(rst), .Z(new_AGEMA_signal_3026) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2961), .B(
        Plaintext_s2[45]), .S(rst), .Z(new_AGEMA_signal_3027) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_0_U1 ( .A(MCOutput[48]), .B(
        Plaintext_s0[48]), .S(rst), .Z(StateRegInput[48]) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2858), .B(
        Plaintext_s1[48]), .S(rst), .Z(new_AGEMA_signal_2944) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2859), .B(
        Plaintext_s2[48]), .S(rst), .Z(new_AGEMA_signal_2945) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_0_U1 ( .A(MCOutput[49]), .B(
        Plaintext_s0[49]), .S(rst), .Z(StateRegInput[49]) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2962), .B(
        Plaintext_s1[49]), .S(rst), .Z(new_AGEMA_signal_3030) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2963), .B(
        Plaintext_s2[49]), .S(rst), .Z(new_AGEMA_signal_3031) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_0_U1 ( .A(MCOutput[52]), .B(
        Plaintext_s0[52]), .S(rst), .Z(StateRegInput[52]) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2862), .B(
        Plaintext_s1[52]), .S(rst), .Z(new_AGEMA_signal_2948) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2863), .B(
        Plaintext_s2[52]), .S(rst), .Z(new_AGEMA_signal_2949) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_0_U1 ( .A(MCOutput[53]), .B(
        Plaintext_s0[53]), .S(rst), .Z(StateRegInput[53]) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2964), .B(
        Plaintext_s1[53]), .S(rst), .Z(new_AGEMA_signal_3034) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2965), .B(
        Plaintext_s2[53]), .S(rst), .Z(new_AGEMA_signal_3035) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_0_U1 ( .A(MCOutput[56]), .B(
        Plaintext_s0[56]), .S(rst), .Z(StateRegInput[56]) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2866), .B(
        Plaintext_s1[56]), .S(rst), .Z(new_AGEMA_signal_2952) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2867), .B(
        Plaintext_s2[56]), .S(rst), .Z(new_AGEMA_signal_2953) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_0_U1 ( .A(MCOutput[57]), .B(
        Plaintext_s0[57]), .S(rst), .Z(StateRegInput[57]) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2966), .B(
        Plaintext_s1[57]), .S(rst), .Z(new_AGEMA_signal_3038) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2967), .B(
        Plaintext_s2[57]), .S(rst), .Z(new_AGEMA_signal_3039) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_0_U1 ( .A(MCOutput[60]), .B(
        Plaintext_s0[60]), .S(rst), .Z(StateRegInput[60]) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3044), .B(
        Plaintext_s1[60]), .S(rst), .Z(new_AGEMA_signal_3066) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3045), .B(
        Plaintext_s2[60]), .S(rst), .Z(new_AGEMA_signal_3067) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_0_U1 ( .A(MCOutput[61]), .B(
        Plaintext_s0[61]), .S(rst), .Z(StateRegInput[61]) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3068), .B(
        Plaintext_s1[61]), .S(rst), .Z(new_AGEMA_signal_3084) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3069), .B(
        Plaintext_s2[61]), .S(rst), .Z(new_AGEMA_signal_3085) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U37 ( .A(new_AGEMA_signal_2028), .B(
        Fresh[98]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U36 ( .A(Fresh[97]), .B(
        SubCellInst_SboxInst_0_Q2), .Z(
        SubCellInst_SboxInst_0_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U35 ( .A(new_AGEMA_signal_2029), .B(
        Fresh[98]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U34 ( .A(Fresh[96]), .B(
        SubCellInst_SboxInst_0_Q2), .Z(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U33 ( .A(Fresh[97]), .B(
        new_AGEMA_signal_2029), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U32 ( .A(new_AGEMA_signal_2028), .B(
        Fresh[96]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U25 ( .A1(Ciphertext_s2[1]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U24 ( .A1(Ciphertext_s2[1]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U23 ( .A1(Ciphertext_s1[1]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U22 ( .A(Fresh[98]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U21 ( .A1(Ciphertext_s1[1]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U20 ( .A1(Ciphertext_s0[1]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U19 ( .A(Fresh[97]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U18 ( .A1(Ciphertext_s0[1]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U17 ( .A(Fresh[96]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U16 ( .A1(new_AGEMA_signal_2029), 
        .A2(Ciphertext_s2[1]), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U15 ( .A1(new_AGEMA_signal_2028), 
        .A2(Ciphertext_s1[1]), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_0_Q2), 
        .A2(Ciphertext_s0[1]), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_n33), .Z(new_AGEMA_signal_2159) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n32), .B(
        SubCellInst_SboxInst_0_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_n30), .Z(new_AGEMA_signal_2158) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n29), .B(
        SubCellInst_SboxInst_0_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_n27), .Z(SubCellInst_SboxInst_0_T1) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n26), .B(
        SubCellInst_SboxInst_0_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_T1), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_L0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2158), 
        .B(new_AGEMA_signal_1934), .Z(new_AGEMA_signal_2286) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2159), 
        .B(new_AGEMA_signal_1935), .Z(new_AGEMA_signal_2287) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U37 ( .A(new_AGEMA_signal_2030), .B(
        Fresh[101]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U36 ( .A(Fresh[100]), .B(
        SubCellInst_SboxInst_0_Q7), .Z(
        SubCellInst_SboxInst_0_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U35 ( .A(new_AGEMA_signal_2031), .B(
        Fresh[101]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U34 ( .A(Fresh[99]), .B(
        SubCellInst_SboxInst_0_Q7), .Z(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U33 ( .A(Fresh[100]), .B(
        new_AGEMA_signal_2031), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U32 ( .A(new_AGEMA_signal_2030), .B(
        Fresh[99]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U25 ( .A1(new_AGEMA_signal_1749), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U24 ( .A1(new_AGEMA_signal_1749), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U23 ( .A1(new_AGEMA_signal_1748), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U22 ( .A(Fresh[101]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U21 ( .A1(new_AGEMA_signal_1748), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_0_Q6), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U19 ( .A(Fresh[100]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_0_Q6), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U17 ( .A(Fresh[99]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U16 ( .A1(new_AGEMA_signal_2031), 
        .A2(new_AGEMA_signal_1749), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U15 ( .A1(new_AGEMA_signal_2030), 
        .A2(new_AGEMA_signal_1748), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_0_Q7), 
        .A2(SubCellInst_SboxInst_0_Q6), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_n33), .Z(new_AGEMA_signal_2161) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n32), .B(
        SubCellInst_SboxInst_0_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_n30), .Z(new_AGEMA_signal_2160) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n29), .B(
        SubCellInst_SboxInst_0_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_n27), .Z(SubCellInst_SboxInst_0_T3) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n26), .B(
        SubCellInst_SboxInst_0_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1748), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1749), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L0), .B(SubCellInst_SboxInst_0_L2), .Z(
        SubCellInst_SboxInst_0_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2286), 
        .B(new_AGEMA_signal_1750), .Z(new_AGEMA_signal_2372) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2287), 
        .B(new_AGEMA_signal_1751), .Z(new_AGEMA_signal_2373) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L0), .B(SubCellInst_SboxInst_0_T3), .Z(
        ShiftRowsOutput[4]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2286), 
        .B(new_AGEMA_signal_2160), .Z(new_AGEMA_signal_2374) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2287), 
        .B(new_AGEMA_signal_2161), .Z(new_AGEMA_signal_2375) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_0_YY_1_), .B(SubCellInst_SboxInst_0_YY_3), .ZN(
        ShiftRowsOutput[5]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2284), .B(new_AGEMA_signal_2372), .Z(new_AGEMA_signal_2488) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2285), .B(new_AGEMA_signal_2373), .Z(new_AGEMA_signal_2489) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U37 ( .A(new_AGEMA_signal_2036), .B(
        Fresh[104]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U36 ( .A(Fresh[103]), .B(
        SubCellInst_SboxInst_1_Q2), .Z(
        SubCellInst_SboxInst_1_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U35 ( .A(new_AGEMA_signal_2037), .B(
        Fresh[104]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U34 ( .A(Fresh[102]), .B(
        SubCellInst_SboxInst_1_Q2), .Z(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U33 ( .A(Fresh[103]), .B(
        new_AGEMA_signal_2037), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U32 ( .A(new_AGEMA_signal_2036), .B(
        Fresh[102]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U25 ( .A1(Ciphertext_s2[5]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U24 ( .A1(Ciphertext_s2[5]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U23 ( .A1(Ciphertext_s1[5]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U22 ( .A(Fresh[104]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U21 ( .A1(Ciphertext_s1[5]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U20 ( .A1(Ciphertext_s0[5]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U19 ( .A(Fresh[103]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U18 ( .A1(Ciphertext_s0[5]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U17 ( .A(Fresh[102]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U16 ( .A1(new_AGEMA_signal_2037), 
        .A2(Ciphertext_s2[5]), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U15 ( .A1(new_AGEMA_signal_2036), 
        .A2(Ciphertext_s1[5]), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_1_Q2), 
        .A2(Ciphertext_s0[5]), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_n33), .Z(new_AGEMA_signal_2167) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n32), .B(
        SubCellInst_SboxInst_1_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_n30), .Z(new_AGEMA_signal_2166) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n29), .B(
        SubCellInst_SboxInst_1_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_n27), .Z(SubCellInst_SboxInst_1_T1) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n26), .B(
        SubCellInst_SboxInst_1_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[5]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[5]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[5]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_T1), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_L0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2166), 
        .B(new_AGEMA_signal_1940), .Z(new_AGEMA_signal_2290) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2167), 
        .B(new_AGEMA_signal_1941), .Z(new_AGEMA_signal_2291) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U37 ( .A(new_AGEMA_signal_2038), .B(
        Fresh[107]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U36 ( .A(Fresh[106]), .B(
        SubCellInst_SboxInst_1_Q7), .Z(
        SubCellInst_SboxInst_1_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U35 ( .A(new_AGEMA_signal_2039), .B(
        Fresh[107]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U34 ( .A(Fresh[105]), .B(
        SubCellInst_SboxInst_1_Q7), .Z(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U33 ( .A(Fresh[106]), .B(
        new_AGEMA_signal_2039), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U32 ( .A(new_AGEMA_signal_2038), .B(
        Fresh[105]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U25 ( .A1(new_AGEMA_signal_1761), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U24 ( .A1(new_AGEMA_signal_1761), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U23 ( .A1(new_AGEMA_signal_1760), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U22 ( .A(Fresh[107]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U21 ( .A1(new_AGEMA_signal_1760), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_1_Q6), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U19 ( .A(Fresh[106]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_1_Q6), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U17 ( .A(Fresh[105]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U16 ( .A1(new_AGEMA_signal_2039), 
        .A2(new_AGEMA_signal_1761), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U15 ( .A1(new_AGEMA_signal_2038), 
        .A2(new_AGEMA_signal_1760), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_1_Q7), 
        .A2(SubCellInst_SboxInst_1_Q6), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_n33), .Z(new_AGEMA_signal_2169) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n32), .B(
        SubCellInst_SboxInst_1_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_n30), .Z(new_AGEMA_signal_2168) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n29), .B(
        SubCellInst_SboxInst_1_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_n27), .Z(SubCellInst_SboxInst_1_T3) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n26), .B(
        SubCellInst_SboxInst_1_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1760), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1761), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L0), .B(SubCellInst_SboxInst_1_L2), .Z(
        SubCellInst_SboxInst_1_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2290), 
        .B(new_AGEMA_signal_1762), .Z(new_AGEMA_signal_2376) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2291), 
        .B(new_AGEMA_signal_1763), .Z(new_AGEMA_signal_2377) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L0), .B(SubCellInst_SboxInst_1_T3), .Z(
        ShiftRowsOutput[8]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2290), 
        .B(new_AGEMA_signal_2168), .Z(new_AGEMA_signal_2378) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2291), 
        .B(new_AGEMA_signal_2169), .Z(new_AGEMA_signal_2379) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_1_YY_1_), .B(SubCellInst_SboxInst_1_YY_3), .ZN(
        ShiftRowsOutput[9]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2288), .B(new_AGEMA_signal_2376), .Z(new_AGEMA_signal_2490) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2289), .B(new_AGEMA_signal_2377), .Z(new_AGEMA_signal_2491) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U37 ( .A(new_AGEMA_signal_2044), .B(
        Fresh[110]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U36 ( .A(Fresh[109]), .B(
        SubCellInst_SboxInst_2_Q2), .Z(
        SubCellInst_SboxInst_2_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U35 ( .A(new_AGEMA_signal_2045), .B(
        Fresh[110]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U34 ( .A(Fresh[108]), .B(
        SubCellInst_SboxInst_2_Q2), .Z(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U33 ( .A(Fresh[109]), .B(
        new_AGEMA_signal_2045), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U32 ( .A(new_AGEMA_signal_2044), .B(
        Fresh[108]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U25 ( .A1(Ciphertext_s2[9]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U24 ( .A1(Ciphertext_s2[9]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U23 ( .A1(Ciphertext_s1[9]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U22 ( .A(Fresh[110]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U21 ( .A1(Ciphertext_s1[9]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U20 ( .A1(Ciphertext_s0[9]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U19 ( .A(Fresh[109]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U18 ( .A1(Ciphertext_s0[9]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U17 ( .A(Fresh[108]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U16 ( .A1(new_AGEMA_signal_2045), 
        .A2(Ciphertext_s2[9]), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U15 ( .A1(new_AGEMA_signal_2044), 
        .A2(Ciphertext_s1[9]), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_2_Q2), 
        .A2(Ciphertext_s0[9]), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_n33), .Z(new_AGEMA_signal_2175) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n32), .B(
        SubCellInst_SboxInst_2_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_n30), .Z(new_AGEMA_signal_2174) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n29), .B(
        SubCellInst_SboxInst_2_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_n27), .Z(SubCellInst_SboxInst_2_T1) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n26), .B(
        SubCellInst_SboxInst_2_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[9]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[9]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[9]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_T1), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_L0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2174), 
        .B(new_AGEMA_signal_1946), .Z(new_AGEMA_signal_2294) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2175), 
        .B(new_AGEMA_signal_1947), .Z(new_AGEMA_signal_2295) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U37 ( .A(new_AGEMA_signal_2046), .B(
        Fresh[113]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U36 ( .A(Fresh[112]), .B(
        SubCellInst_SboxInst_2_Q7), .Z(
        SubCellInst_SboxInst_2_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U35 ( .A(new_AGEMA_signal_2047), .B(
        Fresh[113]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U34 ( .A(Fresh[111]), .B(
        SubCellInst_SboxInst_2_Q7), .Z(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U33 ( .A(Fresh[112]), .B(
        new_AGEMA_signal_2047), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U32 ( .A(new_AGEMA_signal_2046), .B(
        Fresh[111]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U25 ( .A1(new_AGEMA_signal_1773), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U24 ( .A1(new_AGEMA_signal_1773), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U23 ( .A1(new_AGEMA_signal_1772), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U22 ( .A(Fresh[113]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U21 ( .A1(new_AGEMA_signal_1772), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_2_Q6), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U19 ( .A(Fresh[112]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_2_Q6), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U17 ( .A(Fresh[111]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U16 ( .A1(new_AGEMA_signal_2047), 
        .A2(new_AGEMA_signal_1773), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U15 ( .A1(new_AGEMA_signal_2046), 
        .A2(new_AGEMA_signal_1772), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_2_Q7), 
        .A2(SubCellInst_SboxInst_2_Q6), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_n33), .Z(new_AGEMA_signal_2177) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n32), .B(
        SubCellInst_SboxInst_2_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_n30), .Z(new_AGEMA_signal_2176) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n29), .B(
        SubCellInst_SboxInst_2_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_n27), .Z(SubCellInst_SboxInst_2_T3) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n26), .B(
        SubCellInst_SboxInst_2_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1772), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1773), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L0), .B(SubCellInst_SboxInst_2_L2), .Z(
        SubCellInst_SboxInst_2_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2294), 
        .B(new_AGEMA_signal_1774), .Z(new_AGEMA_signal_2380) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2295), 
        .B(new_AGEMA_signal_1775), .Z(new_AGEMA_signal_2381) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L0), .B(SubCellInst_SboxInst_2_T3), .Z(
        ShiftRowsOutput[12]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2294), 
        .B(new_AGEMA_signal_2176), .Z(new_AGEMA_signal_2382) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2295), 
        .B(new_AGEMA_signal_2177), .Z(new_AGEMA_signal_2383) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_2_YY_1_), .B(SubCellInst_SboxInst_2_YY_3), .ZN(
        ShiftRowsOutput[13]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2292), .B(new_AGEMA_signal_2380), .Z(new_AGEMA_signal_2492) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2293), .B(new_AGEMA_signal_2381), .Z(new_AGEMA_signal_2493) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U37 ( .A(new_AGEMA_signal_2052), .B(
        Fresh[116]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U36 ( .A(Fresh[115]), .B(
        SubCellInst_SboxInst_3_Q2), .Z(
        SubCellInst_SboxInst_3_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U35 ( .A(new_AGEMA_signal_2053), .B(
        Fresh[116]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U34 ( .A(Fresh[114]), .B(
        SubCellInst_SboxInst_3_Q2), .Z(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U33 ( .A(Fresh[115]), .B(
        new_AGEMA_signal_2053), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U32 ( .A(new_AGEMA_signal_2052), .B(
        Fresh[114]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U25 ( .A1(Ciphertext_s2[13]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U24 ( .A1(Ciphertext_s2[13]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U23 ( .A1(Ciphertext_s1[13]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U22 ( .A(Fresh[116]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U21 ( .A1(Ciphertext_s1[13]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U20 ( .A1(Ciphertext_s0[13]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U19 ( .A(Fresh[115]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U18 ( .A1(Ciphertext_s0[13]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U17 ( .A(Fresh[114]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U16 ( .A1(new_AGEMA_signal_2053), 
        .A2(Ciphertext_s2[13]), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U15 ( .A1(new_AGEMA_signal_2052), 
        .A2(Ciphertext_s1[13]), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_3_Q2), 
        .A2(Ciphertext_s0[13]), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_n33), .Z(new_AGEMA_signal_2183) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n32), .B(
        SubCellInst_SboxInst_3_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_n30), .Z(new_AGEMA_signal_2182) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n29), .B(
        SubCellInst_SboxInst_3_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_n27), .Z(SubCellInst_SboxInst_3_T1) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n26), .B(
        SubCellInst_SboxInst_3_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[13]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[13]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[13]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_T1), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_L0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2182), 
        .B(new_AGEMA_signal_1952), .Z(new_AGEMA_signal_2298) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2183), 
        .B(new_AGEMA_signal_1953), .Z(new_AGEMA_signal_2299) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U37 ( .A(new_AGEMA_signal_2054), .B(
        Fresh[119]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U36 ( .A(Fresh[118]), .B(
        SubCellInst_SboxInst_3_Q7), .Z(
        SubCellInst_SboxInst_3_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U35 ( .A(new_AGEMA_signal_2055), .B(
        Fresh[119]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U34 ( .A(Fresh[117]), .B(
        SubCellInst_SboxInst_3_Q7), .Z(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U33 ( .A(Fresh[118]), .B(
        new_AGEMA_signal_2055), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U32 ( .A(new_AGEMA_signal_2054), .B(
        Fresh[117]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U25 ( .A1(new_AGEMA_signal_1785), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U24 ( .A1(new_AGEMA_signal_1785), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U23 ( .A1(new_AGEMA_signal_1784), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U22 ( .A(Fresh[119]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U21 ( .A1(new_AGEMA_signal_1784), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_3_Q6), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U19 ( .A(Fresh[118]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_3_Q6), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U17 ( .A(Fresh[117]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U16 ( .A1(new_AGEMA_signal_2055), 
        .A2(new_AGEMA_signal_1785), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U15 ( .A1(new_AGEMA_signal_2054), 
        .A2(new_AGEMA_signal_1784), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_3_Q7), 
        .A2(SubCellInst_SboxInst_3_Q6), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_n33), .Z(new_AGEMA_signal_2185) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n32), .B(
        SubCellInst_SboxInst_3_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_n30), .Z(new_AGEMA_signal_2184) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n29), .B(
        SubCellInst_SboxInst_3_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_n27), .Z(SubCellInst_SboxInst_3_T3) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n26), .B(
        SubCellInst_SboxInst_3_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1784), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1785), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L0), .B(SubCellInst_SboxInst_3_L2), .Z(
        SubCellInst_SboxInst_3_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2298), 
        .B(new_AGEMA_signal_1786), .Z(new_AGEMA_signal_2384) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2299), 
        .B(new_AGEMA_signal_1787), .Z(new_AGEMA_signal_2385) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L0), .B(SubCellInst_SboxInst_3_T3), .Z(
        ShiftRowsOutput[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2298), 
        .B(new_AGEMA_signal_2184), .Z(new_AGEMA_signal_2386) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2299), 
        .B(new_AGEMA_signal_2185), .Z(new_AGEMA_signal_2387) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_3_YY_1_), .B(SubCellInst_SboxInst_3_YY_3), .ZN(
        ShiftRowsOutput[1]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2296), .B(new_AGEMA_signal_2384), .Z(new_AGEMA_signal_2494) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2297), .B(new_AGEMA_signal_2385), .Z(new_AGEMA_signal_2495) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U37 ( .A(new_AGEMA_signal_2060), .B(
        Fresh[122]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U36 ( .A(Fresh[121]), .B(
        SubCellInst_SboxInst_4_Q2), .Z(
        SubCellInst_SboxInst_4_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U35 ( .A(new_AGEMA_signal_2061), .B(
        Fresh[122]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U34 ( .A(Fresh[120]), .B(
        SubCellInst_SboxInst_4_Q2), .Z(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U33 ( .A(Fresh[121]), .B(
        new_AGEMA_signal_2061), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U32 ( .A(new_AGEMA_signal_2060), .B(
        Fresh[120]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U25 ( .A1(Ciphertext_s2[17]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U24 ( .A1(Ciphertext_s2[17]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U23 ( .A1(Ciphertext_s1[17]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U22 ( .A(Fresh[122]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U21 ( .A1(Ciphertext_s1[17]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U20 ( .A1(Ciphertext_s0[17]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U19 ( .A(Fresh[121]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U18 ( .A1(Ciphertext_s0[17]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U17 ( .A(Fresh[120]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U16 ( .A1(new_AGEMA_signal_2061), 
        .A2(Ciphertext_s2[17]), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U15 ( .A1(new_AGEMA_signal_2060), 
        .A2(Ciphertext_s1[17]), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_4_Q2), 
        .A2(Ciphertext_s0[17]), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_n33), .Z(new_AGEMA_signal_2191) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n32), .B(
        SubCellInst_SboxInst_4_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_n30), .Z(new_AGEMA_signal_2190) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n29), .B(
        SubCellInst_SboxInst_4_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_n27), .Z(SubCellInst_SboxInst_4_T1) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n26), .B(
        SubCellInst_SboxInst_4_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[17]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[17]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[17]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_T1), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_L0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2190), 
        .B(new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2302) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2191), 
        .B(new_AGEMA_signal_1959), .Z(new_AGEMA_signal_2303) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U37 ( .A(new_AGEMA_signal_2062), .B(
        Fresh[125]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U36 ( .A(Fresh[124]), .B(
        SubCellInst_SboxInst_4_Q7), .Z(
        SubCellInst_SboxInst_4_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U35 ( .A(new_AGEMA_signal_2063), .B(
        Fresh[125]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U34 ( .A(Fresh[123]), .B(
        SubCellInst_SboxInst_4_Q7), .Z(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U33 ( .A(Fresh[124]), .B(
        new_AGEMA_signal_2063), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U32 ( .A(new_AGEMA_signal_2062), .B(
        Fresh[123]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U25 ( .A1(new_AGEMA_signal_1797), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U24 ( .A1(new_AGEMA_signal_1797), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U23 ( .A1(new_AGEMA_signal_1796), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U22 ( .A(Fresh[125]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U21 ( .A1(new_AGEMA_signal_1796), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_4_Q6), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U19 ( .A(Fresh[124]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_4_Q6), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U17 ( .A(Fresh[123]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U16 ( .A1(new_AGEMA_signal_2063), 
        .A2(new_AGEMA_signal_1797), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U15 ( .A1(new_AGEMA_signal_2062), 
        .A2(new_AGEMA_signal_1796), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_4_Q7), 
        .A2(SubCellInst_SboxInst_4_Q6), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_n33), .Z(new_AGEMA_signal_2193) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n32), .B(
        SubCellInst_SboxInst_4_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_n30), .Z(new_AGEMA_signal_2192) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n29), .B(
        SubCellInst_SboxInst_4_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_n27), .Z(SubCellInst_SboxInst_4_T3) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n26), .B(
        SubCellInst_SboxInst_4_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1796), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1797), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L0), .B(SubCellInst_SboxInst_4_L2), .Z(
        SubCellInst_SboxInst_4_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2302), 
        .B(new_AGEMA_signal_1798), .Z(new_AGEMA_signal_2388) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2303), 
        .B(new_AGEMA_signal_1799), .Z(new_AGEMA_signal_2389) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L0), .B(SubCellInst_SboxInst_4_T3), .Z(
        ShiftRowsOutput[24]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2302), 
        .B(new_AGEMA_signal_2192), .Z(new_AGEMA_signal_2390) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2303), 
        .B(new_AGEMA_signal_2193), .Z(new_AGEMA_signal_2391) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_4_YY_1_), .B(SubCellInst_SboxInst_4_YY_3), .ZN(
        ShiftRowsOutput[25]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2300), .B(new_AGEMA_signal_2388), .Z(new_AGEMA_signal_2496) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2301), .B(new_AGEMA_signal_2389), .Z(new_AGEMA_signal_2497) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U37 ( .A(new_AGEMA_signal_2068), .B(
        Fresh[128]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U36 ( .A(Fresh[127]), .B(
        SubCellInst_SboxInst_5_Q2), .Z(
        SubCellInst_SboxInst_5_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U35 ( .A(new_AGEMA_signal_2069), .B(
        Fresh[128]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U34 ( .A(Fresh[126]), .B(
        SubCellInst_SboxInst_5_Q2), .Z(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U33 ( .A(Fresh[127]), .B(
        new_AGEMA_signal_2069), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U32 ( .A(new_AGEMA_signal_2068), .B(
        Fresh[126]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U25 ( .A1(Ciphertext_s2[21]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U24 ( .A1(Ciphertext_s2[21]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U23 ( .A1(Ciphertext_s1[21]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U22 ( .A(Fresh[128]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U21 ( .A1(Ciphertext_s1[21]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U20 ( .A1(Ciphertext_s0[21]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U19 ( .A(Fresh[127]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U18 ( .A1(Ciphertext_s0[21]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U17 ( .A(Fresh[126]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U16 ( .A1(new_AGEMA_signal_2069), 
        .A2(Ciphertext_s2[21]), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U15 ( .A1(new_AGEMA_signal_2068), 
        .A2(Ciphertext_s1[21]), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_5_Q2), 
        .A2(Ciphertext_s0[21]), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_n33), .Z(new_AGEMA_signal_2199) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n32), .B(
        SubCellInst_SboxInst_5_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_n30), .Z(new_AGEMA_signal_2198) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n29), .B(
        SubCellInst_SboxInst_5_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_n27), .Z(SubCellInst_SboxInst_5_T1) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n26), .B(
        SubCellInst_SboxInst_5_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[21]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[21]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[21]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_T1), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_L0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2198), 
        .B(new_AGEMA_signal_1964), .Z(new_AGEMA_signal_2306) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2199), 
        .B(new_AGEMA_signal_1965), .Z(new_AGEMA_signal_2307) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U37 ( .A(new_AGEMA_signal_2070), .B(
        Fresh[131]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U36 ( .A(Fresh[130]), .B(
        SubCellInst_SboxInst_5_Q7), .Z(
        SubCellInst_SboxInst_5_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U35 ( .A(new_AGEMA_signal_2071), .B(
        Fresh[131]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U34 ( .A(Fresh[129]), .B(
        SubCellInst_SboxInst_5_Q7), .Z(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U33 ( .A(Fresh[130]), .B(
        new_AGEMA_signal_2071), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U32 ( .A(new_AGEMA_signal_2070), .B(
        Fresh[129]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U25 ( .A1(new_AGEMA_signal_1809), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U24 ( .A1(new_AGEMA_signal_1809), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U23 ( .A1(new_AGEMA_signal_1808), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U22 ( .A(Fresh[131]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U21 ( .A1(new_AGEMA_signal_1808), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_5_Q6), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U19 ( .A(Fresh[130]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_5_Q6), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U17 ( .A(Fresh[129]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U16 ( .A1(new_AGEMA_signal_2071), 
        .A2(new_AGEMA_signal_1809), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U15 ( .A1(new_AGEMA_signal_2070), 
        .A2(new_AGEMA_signal_1808), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_5_Q7), 
        .A2(SubCellInst_SboxInst_5_Q6), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_n33), .Z(new_AGEMA_signal_2201) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n32), .B(
        SubCellInst_SboxInst_5_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_n30), .Z(new_AGEMA_signal_2200) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n29), .B(
        SubCellInst_SboxInst_5_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_n27), .Z(SubCellInst_SboxInst_5_T3) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n26), .B(
        SubCellInst_SboxInst_5_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1808), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1809), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L0), .B(SubCellInst_SboxInst_5_L2), .Z(
        SubCellInst_SboxInst_5_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2306), 
        .B(new_AGEMA_signal_1810), .Z(new_AGEMA_signal_2392) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2307), 
        .B(new_AGEMA_signal_1811), .Z(new_AGEMA_signal_2393) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L0), .B(SubCellInst_SboxInst_5_T3), .Z(
        ShiftRowsOutput[28]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2306), 
        .B(new_AGEMA_signal_2200), .Z(new_AGEMA_signal_2394) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2307), 
        .B(new_AGEMA_signal_2201), .Z(new_AGEMA_signal_2395) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_5_YY_1_), .B(SubCellInst_SboxInst_5_YY_3), .ZN(
        ShiftRowsOutput[29]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2304), .B(new_AGEMA_signal_2392), .Z(new_AGEMA_signal_2498) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2305), .B(new_AGEMA_signal_2393), .Z(new_AGEMA_signal_2499) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U37 ( .A(new_AGEMA_signal_2076), .B(
        Fresh[134]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U36 ( .A(Fresh[133]), .B(
        SubCellInst_SboxInst_6_Q2), .Z(
        SubCellInst_SboxInst_6_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U35 ( .A(new_AGEMA_signal_2077), .B(
        Fresh[134]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U34 ( .A(Fresh[132]), .B(
        SubCellInst_SboxInst_6_Q2), .Z(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U33 ( .A(Fresh[133]), .B(
        new_AGEMA_signal_2077), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U32 ( .A(new_AGEMA_signal_2076), .B(
        Fresh[132]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U25 ( .A1(Ciphertext_s2[25]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U24 ( .A1(Ciphertext_s2[25]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U23 ( .A1(Ciphertext_s1[25]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U22 ( .A(Fresh[134]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U21 ( .A1(Ciphertext_s1[25]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U20 ( .A1(Ciphertext_s0[25]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U19 ( .A(Fresh[133]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U18 ( .A1(Ciphertext_s0[25]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U17 ( .A(Fresh[132]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U16 ( .A1(new_AGEMA_signal_2077), 
        .A2(Ciphertext_s2[25]), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U15 ( .A1(new_AGEMA_signal_2076), 
        .A2(Ciphertext_s1[25]), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_6_Q2), 
        .A2(Ciphertext_s0[25]), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_n33), .Z(new_AGEMA_signal_2207) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n32), .B(
        SubCellInst_SboxInst_6_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_n30), .Z(new_AGEMA_signal_2206) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n29), .B(
        SubCellInst_SboxInst_6_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_n27), .Z(SubCellInst_SboxInst_6_T1) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n26), .B(
        SubCellInst_SboxInst_6_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[25]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[25]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[25]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_T1), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_L0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2206), 
        .B(new_AGEMA_signal_1970), .Z(new_AGEMA_signal_2310) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2207), 
        .B(new_AGEMA_signal_1971), .Z(new_AGEMA_signal_2311) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U37 ( .A(new_AGEMA_signal_2078), .B(
        Fresh[137]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U36 ( .A(Fresh[136]), .B(
        SubCellInst_SboxInst_6_Q7), .Z(
        SubCellInst_SboxInst_6_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U35 ( .A(new_AGEMA_signal_2079), .B(
        Fresh[137]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U34 ( .A(Fresh[135]), .B(
        SubCellInst_SboxInst_6_Q7), .Z(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U33 ( .A(Fresh[136]), .B(
        new_AGEMA_signal_2079), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U32 ( .A(new_AGEMA_signal_2078), .B(
        Fresh[135]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U25 ( .A1(new_AGEMA_signal_1821), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U24 ( .A1(new_AGEMA_signal_1821), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U23 ( .A1(new_AGEMA_signal_1820), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U22 ( .A(Fresh[137]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U21 ( .A1(new_AGEMA_signal_1820), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_6_Q6), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U19 ( .A(Fresh[136]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_6_Q6), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U17 ( .A(Fresh[135]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U16 ( .A1(new_AGEMA_signal_2079), 
        .A2(new_AGEMA_signal_1821), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U15 ( .A1(new_AGEMA_signal_2078), 
        .A2(new_AGEMA_signal_1820), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_6_Q7), 
        .A2(SubCellInst_SboxInst_6_Q6), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_n33), .Z(new_AGEMA_signal_2209) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n32), .B(
        SubCellInst_SboxInst_6_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_n30), .Z(new_AGEMA_signal_2208) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n29), .B(
        SubCellInst_SboxInst_6_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_n27), .Z(SubCellInst_SboxInst_6_T3) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n26), .B(
        SubCellInst_SboxInst_6_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1820), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1821), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L0), .B(SubCellInst_SboxInst_6_L2), .Z(
        SubCellInst_SboxInst_6_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2310), 
        .B(new_AGEMA_signal_1822), .Z(new_AGEMA_signal_2396) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2311), 
        .B(new_AGEMA_signal_1823), .Z(new_AGEMA_signal_2397) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L0), .B(SubCellInst_SboxInst_6_T3), .Z(
        ShiftRowsOutput[16]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2310), 
        .B(new_AGEMA_signal_2208), .Z(new_AGEMA_signal_2398) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2311), 
        .B(new_AGEMA_signal_2209), .Z(new_AGEMA_signal_2399) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_6_YY_1_), .B(SubCellInst_SboxInst_6_YY_3), .ZN(
        ShiftRowsOutput[17]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2308), .B(new_AGEMA_signal_2396), .Z(new_AGEMA_signal_2500) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2309), .B(new_AGEMA_signal_2397), .Z(new_AGEMA_signal_2501) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U37 ( .A(new_AGEMA_signal_2084), .B(
        Fresh[140]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U36 ( .A(Fresh[139]), .B(
        SubCellInst_SboxInst_7_Q2), .Z(
        SubCellInst_SboxInst_7_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U35 ( .A(new_AGEMA_signal_2085), .B(
        Fresh[140]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U34 ( .A(Fresh[138]), .B(
        SubCellInst_SboxInst_7_Q2), .Z(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U33 ( .A(Fresh[139]), .B(
        new_AGEMA_signal_2085), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U32 ( .A(new_AGEMA_signal_2084), .B(
        Fresh[138]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U25 ( .A1(Ciphertext_s2[29]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U24 ( .A1(Ciphertext_s2[29]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U23 ( .A1(Ciphertext_s1[29]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U22 ( .A(Fresh[140]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U21 ( .A1(Ciphertext_s1[29]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U20 ( .A1(Ciphertext_s0[29]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U19 ( .A(Fresh[139]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U18 ( .A1(Ciphertext_s0[29]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U17 ( .A(Fresh[138]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U16 ( .A1(new_AGEMA_signal_2085), 
        .A2(Ciphertext_s2[29]), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U15 ( .A1(new_AGEMA_signal_2084), 
        .A2(Ciphertext_s1[29]), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_7_Q2), 
        .A2(Ciphertext_s0[29]), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_n33), .Z(new_AGEMA_signal_2215) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n32), .B(
        SubCellInst_SboxInst_7_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_n30), .Z(new_AGEMA_signal_2214) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n29), .B(
        SubCellInst_SboxInst_7_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_n27), .Z(SubCellInst_SboxInst_7_T1) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n26), .B(
        SubCellInst_SboxInst_7_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[29]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[29]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[29]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_T1), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_L0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2214), 
        .B(new_AGEMA_signal_1976), .Z(new_AGEMA_signal_2314) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2215), 
        .B(new_AGEMA_signal_1977), .Z(new_AGEMA_signal_2315) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U37 ( .A(new_AGEMA_signal_2086), .B(
        Fresh[143]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U36 ( .A(Fresh[142]), .B(
        SubCellInst_SboxInst_7_Q7), .Z(
        SubCellInst_SboxInst_7_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U35 ( .A(new_AGEMA_signal_2087), .B(
        Fresh[143]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U34 ( .A(Fresh[141]), .B(
        SubCellInst_SboxInst_7_Q7), .Z(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U33 ( .A(Fresh[142]), .B(
        new_AGEMA_signal_2087), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U32 ( .A(new_AGEMA_signal_2086), .B(
        Fresh[141]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U25 ( .A1(new_AGEMA_signal_1833), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U24 ( .A1(new_AGEMA_signal_1833), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U23 ( .A1(new_AGEMA_signal_1832), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U22 ( .A(Fresh[143]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U21 ( .A1(new_AGEMA_signal_1832), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_7_Q6), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U19 ( .A(Fresh[142]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_7_Q6), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U17 ( .A(Fresh[141]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U16 ( .A1(new_AGEMA_signal_2087), 
        .A2(new_AGEMA_signal_1833), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U15 ( .A1(new_AGEMA_signal_2086), 
        .A2(new_AGEMA_signal_1832), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_7_Q7), 
        .A2(SubCellInst_SboxInst_7_Q6), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_n33), .Z(new_AGEMA_signal_2217) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n32), .B(
        SubCellInst_SboxInst_7_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_n30), .Z(new_AGEMA_signal_2216) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n29), .B(
        SubCellInst_SboxInst_7_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_n27), .Z(SubCellInst_SboxInst_7_T3) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n26), .B(
        SubCellInst_SboxInst_7_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1832), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1833), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L0), .B(SubCellInst_SboxInst_7_L2), .Z(
        SubCellInst_SboxInst_7_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2314), 
        .B(new_AGEMA_signal_1834), .Z(new_AGEMA_signal_2400) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2315), 
        .B(new_AGEMA_signal_1835), .Z(new_AGEMA_signal_2401) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L0), .B(SubCellInst_SboxInst_7_T3), .Z(
        ShiftRowsOutput[20]) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2314), 
        .B(new_AGEMA_signal_2216), .Z(new_AGEMA_signal_2402) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2315), 
        .B(new_AGEMA_signal_2217), .Z(new_AGEMA_signal_2403) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_7_YY_1_), .B(SubCellInst_SboxInst_7_YY_3), .ZN(
        SubCellOutput_29) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2312), .B(new_AGEMA_signal_2400), .Z(new_AGEMA_signal_2594) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2313), .B(new_AGEMA_signal_2401), .Z(new_AGEMA_signal_2595) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U37 ( .A(new_AGEMA_signal_2092), .B(
        Fresh[146]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U36 ( .A(Fresh[145]), .B(
        SubCellInst_SboxInst_8_Q2), .Z(
        SubCellInst_SboxInst_8_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U35 ( .A(new_AGEMA_signal_2093), .B(
        Fresh[146]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U34 ( .A(Fresh[144]), .B(
        SubCellInst_SboxInst_8_Q2), .Z(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U33 ( .A(Fresh[145]), .B(
        new_AGEMA_signal_2093), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U32 ( .A(new_AGEMA_signal_2092), .B(
        Fresh[144]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U25 ( .A1(Ciphertext_s2[33]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U24 ( .A1(Ciphertext_s2[33]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U23 ( .A1(Ciphertext_s1[33]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U22 ( .A(Fresh[146]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U21 ( .A1(Ciphertext_s1[33]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U20 ( .A1(Ciphertext_s0[33]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U19 ( .A(Fresh[145]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U18 ( .A1(Ciphertext_s0[33]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U17 ( .A(Fresh[144]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U16 ( .A1(new_AGEMA_signal_2093), 
        .A2(Ciphertext_s2[33]), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U15 ( .A1(new_AGEMA_signal_2092), 
        .A2(Ciphertext_s1[33]), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_8_Q2), 
        .A2(Ciphertext_s0[33]), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_n33), .Z(new_AGEMA_signal_2223) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n32), .B(
        SubCellInst_SboxInst_8_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_n30), .Z(new_AGEMA_signal_2222) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n29), .B(
        SubCellInst_SboxInst_8_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_n27), .Z(SubCellInst_SboxInst_8_T1) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n26), .B(
        SubCellInst_SboxInst_8_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[33]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[33]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[33]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_T1), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_L0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2222), 
        .B(new_AGEMA_signal_1982), .Z(new_AGEMA_signal_2318) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2223), 
        .B(new_AGEMA_signal_1983), .Z(new_AGEMA_signal_2319) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U37 ( .A(new_AGEMA_signal_2094), .B(
        Fresh[149]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U36 ( .A(Fresh[148]), .B(
        SubCellInst_SboxInst_8_Q7), .Z(
        SubCellInst_SboxInst_8_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U35 ( .A(new_AGEMA_signal_2095), .B(
        Fresh[149]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U34 ( .A(Fresh[147]), .B(
        SubCellInst_SboxInst_8_Q7), .Z(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U33 ( .A(Fresh[148]), .B(
        new_AGEMA_signal_2095), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U32 ( .A(new_AGEMA_signal_2094), .B(
        Fresh[147]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U25 ( .A1(new_AGEMA_signal_1845), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U24 ( .A1(new_AGEMA_signal_1845), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U23 ( .A1(new_AGEMA_signal_1844), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U22 ( .A(Fresh[149]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U21 ( .A1(new_AGEMA_signal_1844), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_8_Q6), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U19 ( .A(Fresh[148]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_8_Q6), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U17 ( .A(Fresh[147]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U16 ( .A1(new_AGEMA_signal_2095), 
        .A2(new_AGEMA_signal_1845), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U15 ( .A1(new_AGEMA_signal_2094), 
        .A2(new_AGEMA_signal_1844), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_8_Q7), 
        .A2(SubCellInst_SboxInst_8_Q6), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_n33), .Z(new_AGEMA_signal_2225) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n32), .B(
        SubCellInst_SboxInst_8_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_n30), .Z(new_AGEMA_signal_2224) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n29), .B(
        SubCellInst_SboxInst_8_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_n27), .Z(SubCellInst_SboxInst_8_T3) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n26), .B(
        SubCellInst_SboxInst_8_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1844), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1845), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L0), .B(SubCellInst_SboxInst_8_L2), .Z(
        SubCellInst_SboxInst_8_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2318), 
        .B(new_AGEMA_signal_1846), .Z(new_AGEMA_signal_2404) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2319), 
        .B(new_AGEMA_signal_1847), .Z(new_AGEMA_signal_2405) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L0), .B(SubCellInst_SboxInst_8_T3), .Z(
        AddRoundConstantOutput[32]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2318), 
        .B(new_AGEMA_signal_2224), .Z(new_AGEMA_signal_2406) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2319), 
        .B(new_AGEMA_signal_2225), .Z(new_AGEMA_signal_2407) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_8_YY_1_), .B(SubCellInst_SboxInst_8_YY_3), .ZN(
        AddRoundConstantOutput[33]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2316), .B(new_AGEMA_signal_2404), .Z(new_AGEMA_signal_2504) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2317), .B(new_AGEMA_signal_2405), .Z(new_AGEMA_signal_2505) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U37 ( .A(new_AGEMA_signal_2100), .B(
        Fresh[152]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U36 ( .A(Fresh[151]), .B(
        SubCellInst_SboxInst_9_Q2), .Z(
        SubCellInst_SboxInst_9_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U35 ( .A(new_AGEMA_signal_2101), .B(
        Fresh[152]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U34 ( .A(Fresh[150]), .B(
        SubCellInst_SboxInst_9_Q2), .Z(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U33 ( .A(Fresh[151]), .B(
        new_AGEMA_signal_2101), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U32 ( .A(new_AGEMA_signal_2100), .B(
        Fresh[150]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U25 ( .A1(Ciphertext_s2[37]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U24 ( .A1(Ciphertext_s2[37]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U23 ( .A1(Ciphertext_s1[37]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U22 ( .A(Fresh[152]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U21 ( .A1(Ciphertext_s1[37]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U20 ( .A1(Ciphertext_s0[37]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U19 ( .A(Fresh[151]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U18 ( .A1(Ciphertext_s0[37]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U17 ( .A(Fresh[150]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U16 ( .A1(new_AGEMA_signal_2101), 
        .A2(Ciphertext_s2[37]), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U15 ( .A1(new_AGEMA_signal_2100), 
        .A2(Ciphertext_s1[37]), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_9_Q2), 
        .A2(Ciphertext_s0[37]), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_n33), .Z(new_AGEMA_signal_2231) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n32), .B(
        SubCellInst_SboxInst_9_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_n30), .Z(new_AGEMA_signal_2230) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n29), .B(
        SubCellInst_SboxInst_9_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_n27), .Z(SubCellInst_SboxInst_9_T1) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n26), .B(
        SubCellInst_SboxInst_9_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[37]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[37]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[37]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_T1), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_L0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2230), 
        .B(new_AGEMA_signal_1988), .Z(new_AGEMA_signal_2322) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2231), 
        .B(new_AGEMA_signal_1989), .Z(new_AGEMA_signal_2323) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U37 ( .A(new_AGEMA_signal_2102), .B(
        Fresh[155]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U36 ( .A(Fresh[154]), .B(
        SubCellInst_SboxInst_9_Q7), .Z(
        SubCellInst_SboxInst_9_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U35 ( .A(new_AGEMA_signal_2103), .B(
        Fresh[155]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U34 ( .A(Fresh[153]), .B(
        SubCellInst_SboxInst_9_Q7), .Z(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U33 ( .A(Fresh[154]), .B(
        new_AGEMA_signal_2103), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U32 ( .A(new_AGEMA_signal_2102), .B(
        Fresh[153]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U25 ( .A1(new_AGEMA_signal_1857), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U24 ( .A1(new_AGEMA_signal_1857), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U23 ( .A1(new_AGEMA_signal_1856), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U22 ( .A(Fresh[155]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U21 ( .A1(new_AGEMA_signal_1856), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_9_Q6), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U19 ( .A(Fresh[154]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_9_Q6), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U17 ( .A(Fresh[153]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U16 ( .A1(new_AGEMA_signal_2103), 
        .A2(new_AGEMA_signal_1857), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U15 ( .A1(new_AGEMA_signal_2102), 
        .A2(new_AGEMA_signal_1856), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_9_Q7), 
        .A2(SubCellInst_SboxInst_9_Q6), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_n33), .Z(new_AGEMA_signal_2233) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n32), .B(
        SubCellInst_SboxInst_9_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_n30), .Z(new_AGEMA_signal_2232) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n29), .B(
        SubCellInst_SboxInst_9_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_n27), .Z(SubCellInst_SboxInst_9_T3) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n26), .B(
        SubCellInst_SboxInst_9_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1856), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1857), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L0), .B(SubCellInst_SboxInst_9_L2), .Z(
        SubCellInst_SboxInst_9_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2322), 
        .B(new_AGEMA_signal_1858), .Z(new_AGEMA_signal_2408) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2323), 
        .B(new_AGEMA_signal_1859), .Z(new_AGEMA_signal_2409) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L0), .B(SubCellInst_SboxInst_9_T3), .Z(
        AddRoundConstantOutput[36]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2322), 
        .B(new_AGEMA_signal_2232), .Z(new_AGEMA_signal_2410) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2323), 
        .B(new_AGEMA_signal_2233), .Z(new_AGEMA_signal_2411) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_9_YY_1_), .B(SubCellInst_SboxInst_9_YY_3), .ZN(
        AddRoundConstantOutput[37]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2320), .B(new_AGEMA_signal_2408), .Z(new_AGEMA_signal_2506) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2321), .B(new_AGEMA_signal_2409), .Z(new_AGEMA_signal_2507) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U37 ( .A(new_AGEMA_signal_2108), .B(
        Fresh[158]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U36 ( .A(Fresh[157]), .B(
        SubCellInst_SboxInst_10_Q2), .Z(
        SubCellInst_SboxInst_10_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U35 ( .A(new_AGEMA_signal_2109), .B(
        Fresh[158]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U34 ( .A(Fresh[156]), .B(
        SubCellInst_SboxInst_10_Q2), .Z(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U33 ( .A(Fresh[157]), .B(
        new_AGEMA_signal_2109), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U32 ( .A(new_AGEMA_signal_2108), .B(
        Fresh[156]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U25 ( .A1(Ciphertext_s2[41]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U24 ( .A1(Ciphertext_s2[41]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U23 ( .A1(Ciphertext_s1[41]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U22 ( .A(Fresh[158]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U21 ( .A1(Ciphertext_s1[41]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U20 ( .A1(Ciphertext_s0[41]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U19 ( .A(Fresh[157]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U18 ( .A1(Ciphertext_s0[41]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U17 ( .A(Fresh[156]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U16 ( .A1(new_AGEMA_signal_2109), 
        .A2(Ciphertext_s2[41]), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U15 ( .A1(new_AGEMA_signal_2108), 
        .A2(Ciphertext_s1[41]), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_10_Q2), .A2(Ciphertext_s0[41]), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_n33), .Z(new_AGEMA_signal_2239) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n32), .B(
        SubCellInst_SboxInst_10_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_n30), .Z(new_AGEMA_signal_2238) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n29), .B(
        SubCellInst_SboxInst_10_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_n27), .Z(SubCellInst_SboxInst_10_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n26), .B(
        SubCellInst_SboxInst_10_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[41]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[41]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[41]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_T1), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_L0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2238), 
        .B(new_AGEMA_signal_1994), .Z(new_AGEMA_signal_2326) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2239), 
        .B(new_AGEMA_signal_1995), .Z(new_AGEMA_signal_2327) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U37 ( .A(new_AGEMA_signal_2110), .B(
        Fresh[161]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U36 ( .A(Fresh[160]), .B(
        SubCellInst_SboxInst_10_Q7), .Z(
        SubCellInst_SboxInst_10_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U35 ( .A(new_AGEMA_signal_2111), .B(
        Fresh[161]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U34 ( .A(Fresh[159]), .B(
        SubCellInst_SboxInst_10_Q7), .Z(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U33 ( .A(Fresh[160]), .B(
        new_AGEMA_signal_2111), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U32 ( .A(new_AGEMA_signal_2110), .B(
        Fresh[159]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U25 ( .A1(new_AGEMA_signal_1869), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U24 ( .A1(new_AGEMA_signal_1869), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U23 ( .A1(new_AGEMA_signal_1868), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U22 ( .A(Fresh[161]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U21 ( .A1(new_AGEMA_signal_1868), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_10_Q6), .A2(SubCellInst_SboxInst_10_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U19 ( .A(Fresh[160]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_10_Q6), .A2(SubCellInst_SboxInst_10_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U17 ( .A(Fresh[159]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U16 ( .A1(new_AGEMA_signal_2111), 
        .A2(new_AGEMA_signal_1869), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U15 ( .A1(new_AGEMA_signal_2110), 
        .A2(new_AGEMA_signal_1868), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_10_Q7), .A2(SubCellInst_SboxInst_10_Q6), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_n33), .Z(new_AGEMA_signal_2241) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n32), .B(
        SubCellInst_SboxInst_10_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_n30), .Z(new_AGEMA_signal_2240) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n29), .B(
        SubCellInst_SboxInst_10_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_n27), .Z(SubCellInst_SboxInst_10_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n26), .B(
        SubCellInst_SboxInst_10_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1868), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1869), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L0), .B(SubCellInst_SboxInst_10_L2), .Z(
        SubCellInst_SboxInst_10_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2326), 
        .B(new_AGEMA_signal_1870), .Z(new_AGEMA_signal_2412) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2327), 
        .B(new_AGEMA_signal_1871), .Z(new_AGEMA_signal_2413) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L0), .B(SubCellInst_SboxInst_10_T3), .Z(
        AddRoundConstantOutput[40]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2326), .B(new_AGEMA_signal_2240), .Z(new_AGEMA_signal_2414) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2327), .B(new_AGEMA_signal_2241), .Z(new_AGEMA_signal_2415) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_10_YY_1_), .B(SubCellInst_SboxInst_10_YY_3), .ZN(
        AddRoundConstantOutput[41]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2324), .B(new_AGEMA_signal_2412), .Z(
        new_AGEMA_signal_2508) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_2325), .B(new_AGEMA_signal_2413), .Z(
        new_AGEMA_signal_2509) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U37 ( .A(new_AGEMA_signal_2116), .B(
        Fresh[164]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U36 ( .A(Fresh[163]), .B(
        SubCellInst_SboxInst_11_Q2), .Z(
        SubCellInst_SboxInst_11_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U35 ( .A(new_AGEMA_signal_2117), .B(
        Fresh[164]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U34 ( .A(Fresh[162]), .B(
        SubCellInst_SboxInst_11_Q2), .Z(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U33 ( .A(Fresh[163]), .B(
        new_AGEMA_signal_2117), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U32 ( .A(new_AGEMA_signal_2116), .B(
        Fresh[162]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U25 ( .A1(Ciphertext_s2[45]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U24 ( .A1(Ciphertext_s2[45]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U23 ( .A1(Ciphertext_s1[45]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U22 ( .A(Fresh[164]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U21 ( .A1(Ciphertext_s1[45]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U20 ( .A1(Ciphertext_s0[45]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U19 ( .A(Fresh[163]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U18 ( .A1(Ciphertext_s0[45]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U17 ( .A(Fresh[162]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U16 ( .A1(new_AGEMA_signal_2117), 
        .A2(Ciphertext_s2[45]), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U15 ( .A1(new_AGEMA_signal_2116), 
        .A2(Ciphertext_s1[45]), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_11_Q2), .A2(Ciphertext_s0[45]), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_n33), .Z(new_AGEMA_signal_2247) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n32), .B(
        SubCellInst_SboxInst_11_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_n30), .Z(new_AGEMA_signal_2246) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n29), .B(
        SubCellInst_SboxInst_11_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_n27), .Z(SubCellInst_SboxInst_11_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n26), .B(
        SubCellInst_SboxInst_11_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[45]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[45]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[45]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_T1), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_L0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2246), 
        .B(new_AGEMA_signal_2000), .Z(new_AGEMA_signal_2330) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2247), 
        .B(new_AGEMA_signal_2001), .Z(new_AGEMA_signal_2331) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U37 ( .A(new_AGEMA_signal_2118), .B(
        Fresh[167]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U36 ( .A(Fresh[166]), .B(
        SubCellInst_SboxInst_11_Q7), .Z(
        SubCellInst_SboxInst_11_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U35 ( .A(new_AGEMA_signal_2119), .B(
        Fresh[167]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U34 ( .A(Fresh[165]), .B(
        SubCellInst_SboxInst_11_Q7), .Z(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U33 ( .A(Fresh[166]), .B(
        new_AGEMA_signal_2119), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U32 ( .A(new_AGEMA_signal_2118), .B(
        Fresh[165]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U25 ( .A1(new_AGEMA_signal_1881), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U24 ( .A1(new_AGEMA_signal_1881), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U23 ( .A1(new_AGEMA_signal_1880), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U22 ( .A(Fresh[167]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U21 ( .A1(new_AGEMA_signal_1880), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_11_Q6), .A2(SubCellInst_SboxInst_11_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U19 ( .A(Fresh[166]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_11_Q6), .A2(SubCellInst_SboxInst_11_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U17 ( .A(Fresh[165]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U16 ( .A1(new_AGEMA_signal_2119), 
        .A2(new_AGEMA_signal_1881), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U15 ( .A1(new_AGEMA_signal_2118), 
        .A2(new_AGEMA_signal_1880), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_11_Q7), .A2(SubCellInst_SboxInst_11_Q6), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_n33), .Z(new_AGEMA_signal_2249) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n32), .B(
        SubCellInst_SboxInst_11_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_n30), .Z(new_AGEMA_signal_2248) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n29), .B(
        SubCellInst_SboxInst_11_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_n27), .Z(SubCellInst_SboxInst_11_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n26), .B(
        SubCellInst_SboxInst_11_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1880), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1881), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L0), .B(SubCellInst_SboxInst_11_L2), .Z(
        SubCellInst_SboxInst_11_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2330), 
        .B(new_AGEMA_signal_1882), .Z(new_AGEMA_signal_2416) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2331), 
        .B(new_AGEMA_signal_1883), .Z(new_AGEMA_signal_2417) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L0), .B(SubCellInst_SboxInst_11_T3), .Z(
        SubCellOutput_44) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2330), .B(new_AGEMA_signal_2248), .Z(new_AGEMA_signal_2418) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2331), .B(new_AGEMA_signal_2249), .Z(new_AGEMA_signal_2419) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_11_YY_1_), .B(SubCellInst_SboxInst_11_YY_3), .ZN(
        SubCellOutput_45) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2328), .B(new_AGEMA_signal_2416), .Z(
        new_AGEMA_signal_2510) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_2329), .B(new_AGEMA_signal_2417), .Z(
        new_AGEMA_signal_2511) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U37 ( .A(new_AGEMA_signal_2124), .B(
        Fresh[170]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U36 ( .A(Fresh[169]), .B(
        SubCellInst_SboxInst_12_Q2), .Z(
        SubCellInst_SboxInst_12_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U35 ( .A(new_AGEMA_signal_2125), .B(
        Fresh[170]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U34 ( .A(Fresh[168]), .B(
        SubCellInst_SboxInst_12_Q2), .Z(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U33 ( .A(Fresh[169]), .B(
        new_AGEMA_signal_2125), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U32 ( .A(new_AGEMA_signal_2124), .B(
        Fresh[168]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U25 ( .A1(Ciphertext_s2[49]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U24 ( .A1(Ciphertext_s2[49]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U23 ( .A1(Ciphertext_s1[49]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U22 ( .A(Fresh[170]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U21 ( .A1(Ciphertext_s1[49]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U20 ( .A1(Ciphertext_s0[49]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U19 ( .A(Fresh[169]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U18 ( .A1(Ciphertext_s0[49]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U17 ( .A(Fresh[168]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U16 ( .A1(new_AGEMA_signal_2125), 
        .A2(Ciphertext_s2[49]), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U15 ( .A1(new_AGEMA_signal_2124), 
        .A2(Ciphertext_s1[49]), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_12_Q2), .A2(Ciphertext_s0[49]), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_n33), .Z(new_AGEMA_signal_2255) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n32), .B(
        SubCellInst_SboxInst_12_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_n30), .Z(new_AGEMA_signal_2254) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n29), .B(
        SubCellInst_SboxInst_12_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_n27), .Z(SubCellInst_SboxInst_12_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n26), .B(
        SubCellInst_SboxInst_12_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[49]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[49]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[49]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_T1), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_L0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2254), 
        .B(new_AGEMA_signal_2006), .Z(new_AGEMA_signal_2334) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2255), 
        .B(new_AGEMA_signal_2007), .Z(new_AGEMA_signal_2335) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U37 ( .A(new_AGEMA_signal_2126), .B(
        Fresh[173]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U36 ( .A(Fresh[172]), .B(
        SubCellInst_SboxInst_12_Q7), .Z(
        SubCellInst_SboxInst_12_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U35 ( .A(new_AGEMA_signal_2127), .B(
        Fresh[173]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U34 ( .A(Fresh[171]), .B(
        SubCellInst_SboxInst_12_Q7), .Z(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U33 ( .A(Fresh[172]), .B(
        new_AGEMA_signal_2127), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U32 ( .A(new_AGEMA_signal_2126), .B(
        Fresh[171]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U25 ( .A1(new_AGEMA_signal_1893), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U24 ( .A1(new_AGEMA_signal_1893), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U23 ( .A1(new_AGEMA_signal_1892), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U22 ( .A(Fresh[173]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U21 ( .A1(new_AGEMA_signal_1892), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_12_Q6), .A2(SubCellInst_SboxInst_12_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U19 ( .A(Fresh[172]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_12_Q6), .A2(SubCellInst_SboxInst_12_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U17 ( .A(Fresh[171]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U16 ( .A1(new_AGEMA_signal_2127), 
        .A2(new_AGEMA_signal_1893), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U15 ( .A1(new_AGEMA_signal_2126), 
        .A2(new_AGEMA_signal_1892), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_12_Q7), .A2(SubCellInst_SboxInst_12_Q6), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_n33), .Z(new_AGEMA_signal_2257) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n32), .B(
        SubCellInst_SboxInst_12_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_n30), .Z(new_AGEMA_signal_2256) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n29), .B(
        SubCellInst_SboxInst_12_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_n27), .Z(SubCellInst_SboxInst_12_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n26), .B(
        SubCellInst_SboxInst_12_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1892), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1893), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L0), .B(SubCellInst_SboxInst_12_L2), .Z(
        SubCellInst_SboxInst_12_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2334), 
        .B(new_AGEMA_signal_1894), .Z(new_AGEMA_signal_2420) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2335), 
        .B(new_AGEMA_signal_1895), .Z(new_AGEMA_signal_2421) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L0), .B(SubCellInst_SboxInst_12_T3), .Z(
        AddRoundConstantOutput[48]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2334), .B(new_AGEMA_signal_2256), .Z(new_AGEMA_signal_2422) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2335), .B(new_AGEMA_signal_2257), .Z(new_AGEMA_signal_2423) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_12_YY_1_), .B(SubCellInst_SboxInst_12_YY_3), .ZN(
        AddRoundConstantOutput[49]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2332), .B(new_AGEMA_signal_2420), .Z(
        new_AGEMA_signal_2512) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_2333), .B(new_AGEMA_signal_2421), .Z(
        new_AGEMA_signal_2513) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U37 ( .A(new_AGEMA_signal_2132), .B(
        Fresh[176]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U36 ( .A(Fresh[175]), .B(
        SubCellInst_SboxInst_13_Q2), .Z(
        SubCellInst_SboxInst_13_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U35 ( .A(new_AGEMA_signal_2133), .B(
        Fresh[176]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U34 ( .A(Fresh[174]), .B(
        SubCellInst_SboxInst_13_Q2), .Z(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U33 ( .A(Fresh[175]), .B(
        new_AGEMA_signal_2133), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U32 ( .A(new_AGEMA_signal_2132), .B(
        Fresh[174]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U25 ( .A1(Ciphertext_s2[53]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U24 ( .A1(Ciphertext_s2[53]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U23 ( .A1(Ciphertext_s1[53]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U22 ( .A(Fresh[176]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U21 ( .A1(Ciphertext_s1[53]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U20 ( .A1(Ciphertext_s0[53]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U19 ( .A(Fresh[175]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U18 ( .A1(Ciphertext_s0[53]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U17 ( .A(Fresh[174]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U16 ( .A1(new_AGEMA_signal_2133), 
        .A2(Ciphertext_s2[53]), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U15 ( .A1(new_AGEMA_signal_2132), 
        .A2(Ciphertext_s1[53]), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_13_Q2), .A2(Ciphertext_s0[53]), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_n33), .Z(new_AGEMA_signal_2263) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n32), .B(
        SubCellInst_SboxInst_13_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_n30), .Z(new_AGEMA_signal_2262) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n29), .B(
        SubCellInst_SboxInst_13_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_n27), .Z(SubCellInst_SboxInst_13_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n26), .B(
        SubCellInst_SboxInst_13_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[53]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[53]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[53]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_T1), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_L0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2262), 
        .B(new_AGEMA_signal_2012), .Z(new_AGEMA_signal_2338) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2263), 
        .B(new_AGEMA_signal_2013), .Z(new_AGEMA_signal_2339) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U37 ( .A(new_AGEMA_signal_2134), .B(
        Fresh[179]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U36 ( .A(Fresh[178]), .B(
        SubCellInst_SboxInst_13_Q7), .Z(
        SubCellInst_SboxInst_13_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U35 ( .A(new_AGEMA_signal_2135), .B(
        Fresh[179]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U34 ( .A(Fresh[177]), .B(
        SubCellInst_SboxInst_13_Q7), .Z(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U33 ( .A(Fresh[178]), .B(
        new_AGEMA_signal_2135), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U32 ( .A(new_AGEMA_signal_2134), .B(
        Fresh[177]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U25 ( .A1(new_AGEMA_signal_1905), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U24 ( .A1(new_AGEMA_signal_1905), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U23 ( .A1(new_AGEMA_signal_1904), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U22 ( .A(Fresh[179]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U21 ( .A1(new_AGEMA_signal_1904), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_13_Q6), .A2(SubCellInst_SboxInst_13_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U19 ( .A(Fresh[178]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_13_Q6), .A2(SubCellInst_SboxInst_13_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U17 ( .A(Fresh[177]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U16 ( .A1(new_AGEMA_signal_2135), 
        .A2(new_AGEMA_signal_1905), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U15 ( .A1(new_AGEMA_signal_2134), 
        .A2(new_AGEMA_signal_1904), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_13_Q7), .A2(SubCellInst_SboxInst_13_Q6), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_n33), .Z(new_AGEMA_signal_2265) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n32), .B(
        SubCellInst_SboxInst_13_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_n30), .Z(new_AGEMA_signal_2264) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n29), .B(
        SubCellInst_SboxInst_13_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_n27), .Z(SubCellInst_SboxInst_13_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n26), .B(
        SubCellInst_SboxInst_13_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1904), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1905), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L0), .B(SubCellInst_SboxInst_13_L2), .Z(
        SubCellInst_SboxInst_13_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2338), 
        .B(new_AGEMA_signal_1906), .Z(new_AGEMA_signal_2424) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2339), 
        .B(new_AGEMA_signal_1907), .Z(new_AGEMA_signal_2425) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L0), .B(SubCellInst_SboxInst_13_T3), .Z(
        AddRoundConstantOutput[52]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2338), .B(new_AGEMA_signal_2264), .Z(new_AGEMA_signal_2426) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2339), .B(new_AGEMA_signal_2265), .Z(new_AGEMA_signal_2427) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_13_YY_1_), .B(SubCellInst_SboxInst_13_YY_3), .ZN(
        AddRoundConstantOutput[53]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2336), .B(new_AGEMA_signal_2424), .Z(
        new_AGEMA_signal_2514) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_2337), .B(new_AGEMA_signal_2425), .Z(
        new_AGEMA_signal_2515) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U37 ( .A(new_AGEMA_signal_2140), .B(
        Fresh[182]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U36 ( .A(Fresh[181]), .B(
        SubCellInst_SboxInst_14_Q2), .Z(
        SubCellInst_SboxInst_14_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U35 ( .A(new_AGEMA_signal_2141), .B(
        Fresh[182]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U34 ( .A(Fresh[180]), .B(
        SubCellInst_SboxInst_14_Q2), .Z(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U33 ( .A(Fresh[181]), .B(
        new_AGEMA_signal_2141), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U32 ( .A(new_AGEMA_signal_2140), .B(
        Fresh[180]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U25 ( .A1(Ciphertext_s2[57]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U24 ( .A1(Ciphertext_s2[57]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U23 ( .A1(Ciphertext_s1[57]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U22 ( .A(Fresh[182]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U21 ( .A1(Ciphertext_s1[57]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U20 ( .A1(Ciphertext_s0[57]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U19 ( .A(Fresh[181]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U18 ( .A1(Ciphertext_s0[57]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U17 ( .A(Fresh[180]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U16 ( .A1(new_AGEMA_signal_2141), 
        .A2(Ciphertext_s2[57]), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U15 ( .A1(new_AGEMA_signal_2140), 
        .A2(Ciphertext_s1[57]), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_14_Q2), .A2(Ciphertext_s0[57]), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_n33), .Z(new_AGEMA_signal_2271) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n32), .B(
        SubCellInst_SboxInst_14_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_n30), .Z(new_AGEMA_signal_2270) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n29), .B(
        SubCellInst_SboxInst_14_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_n27), .Z(SubCellInst_SboxInst_14_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n26), .B(
        SubCellInst_SboxInst_14_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[57]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[57]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[57]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_T1), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_L0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2270), 
        .B(new_AGEMA_signal_2018), .Z(new_AGEMA_signal_2342) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2271), 
        .B(new_AGEMA_signal_2019), .Z(new_AGEMA_signal_2343) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U37 ( .A(new_AGEMA_signal_2142), .B(
        Fresh[185]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U36 ( .A(Fresh[184]), .B(
        SubCellInst_SboxInst_14_Q7), .Z(
        SubCellInst_SboxInst_14_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U35 ( .A(new_AGEMA_signal_2143), .B(
        Fresh[185]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U34 ( .A(Fresh[183]), .B(
        SubCellInst_SboxInst_14_Q7), .Z(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U33 ( .A(Fresh[184]), .B(
        new_AGEMA_signal_2143), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U32 ( .A(new_AGEMA_signal_2142), .B(
        Fresh[183]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U25 ( .A1(new_AGEMA_signal_1917), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U24 ( .A1(new_AGEMA_signal_1917), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U23 ( .A1(new_AGEMA_signal_1916), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U22 ( .A(Fresh[185]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U21 ( .A1(new_AGEMA_signal_1916), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_14_Q6), .A2(SubCellInst_SboxInst_14_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U19 ( .A(Fresh[184]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_14_Q6), .A2(SubCellInst_SboxInst_14_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U17 ( .A(Fresh[183]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U16 ( .A1(new_AGEMA_signal_2143), 
        .A2(new_AGEMA_signal_1917), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U15 ( .A1(new_AGEMA_signal_2142), 
        .A2(new_AGEMA_signal_1916), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_14_Q7), .A2(SubCellInst_SboxInst_14_Q6), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_n33), .Z(new_AGEMA_signal_2273) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n32), .B(
        SubCellInst_SboxInst_14_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_n30), .Z(new_AGEMA_signal_2272) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n29), .B(
        SubCellInst_SboxInst_14_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_n27), .Z(SubCellInst_SboxInst_14_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n26), .B(
        SubCellInst_SboxInst_14_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1916), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1917), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L0), .B(SubCellInst_SboxInst_14_L2), .Z(
        SubCellInst_SboxInst_14_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2342), 
        .B(new_AGEMA_signal_1918), .Z(new_AGEMA_signal_2428) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2343), 
        .B(new_AGEMA_signal_1919), .Z(new_AGEMA_signal_2429) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L0), .B(SubCellInst_SboxInst_14_T3), .Z(
        AddRoundConstantOutput[56]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2342), .B(new_AGEMA_signal_2272), .Z(new_AGEMA_signal_2430) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2343), .B(new_AGEMA_signal_2273), .Z(new_AGEMA_signal_2431) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_14_YY_1_), .B(SubCellInst_SboxInst_14_YY_3), .ZN(
        AddRoundConstantOutput[57]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2340), .B(new_AGEMA_signal_2428), .Z(
        new_AGEMA_signal_2516) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_2341), .B(new_AGEMA_signal_2429), .Z(
        new_AGEMA_signal_2517) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U37 ( .A(new_AGEMA_signal_2148), .B(
        Fresh[188]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U36 ( .A(Fresh[187]), .B(
        SubCellInst_SboxInst_15_Q2), .Z(
        SubCellInst_SboxInst_15_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U35 ( .A(new_AGEMA_signal_2149), .B(
        Fresh[188]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U34 ( .A(Fresh[186]), .B(
        SubCellInst_SboxInst_15_Q2), .Z(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U33 ( .A(Fresh[187]), .B(
        new_AGEMA_signal_2149), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U32 ( .A(new_AGEMA_signal_2148), .B(
        Fresh[186]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U25 ( .A1(Ciphertext_s2[61]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U24 ( .A1(Ciphertext_s2[61]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U23 ( .A1(Ciphertext_s1[61]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U22 ( .A(Fresh[188]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U21 ( .A1(Ciphertext_s1[61]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U20 ( .A1(Ciphertext_s0[61]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U19 ( .A(Fresh[187]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U18 ( .A1(Ciphertext_s0[61]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U17 ( .A(Fresh[186]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U16 ( .A1(new_AGEMA_signal_2149), 
        .A2(Ciphertext_s2[61]), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U15 ( .A1(new_AGEMA_signal_2148), 
        .A2(Ciphertext_s1[61]), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_15_Q2), .A2(Ciphertext_s0[61]), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_n33), .Z(new_AGEMA_signal_2279) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n32), .B(
        SubCellInst_SboxInst_15_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_n30), .Z(new_AGEMA_signal_2278) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n29), .B(
        SubCellInst_SboxInst_15_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_n27), .Z(SubCellInst_SboxInst_15_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n26), .B(
        SubCellInst_SboxInst_15_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[61]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[61]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[61]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_T1), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_L0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2278), 
        .B(new_AGEMA_signal_2024), .Z(new_AGEMA_signal_2346) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2279), 
        .B(new_AGEMA_signal_2025), .Z(new_AGEMA_signal_2347) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U37 ( .A(new_AGEMA_signal_2150), .B(
        Fresh[191]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U36 ( .A(Fresh[190]), .B(
        SubCellInst_SboxInst_15_Q7), .Z(
        SubCellInst_SboxInst_15_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U35 ( .A(new_AGEMA_signal_2151), .B(
        Fresh[191]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U34 ( .A(Fresh[189]), .B(
        SubCellInst_SboxInst_15_Q7), .Z(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U33 ( .A(Fresh[190]), .B(
        new_AGEMA_signal_2151), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U32 ( .A(new_AGEMA_signal_2150), .B(
        Fresh[189]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U25 ( .A1(new_AGEMA_signal_1929), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U24 ( .A1(new_AGEMA_signal_1929), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U23 ( .A1(new_AGEMA_signal_1928), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U22 ( .A(Fresh[191]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U21 ( .A1(new_AGEMA_signal_1928), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U20 ( .A1(SubCellInst_SboxInst_15_Q6), .A2(SubCellInst_SboxInst_15_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U19 ( .A(Fresh[190]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U18 ( .A1(SubCellInst_SboxInst_15_Q6), .A2(SubCellInst_SboxInst_15_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U17 ( .A(Fresh[189]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U16 ( .A1(new_AGEMA_signal_2151), 
        .A2(new_AGEMA_signal_1929), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U15 ( .A1(new_AGEMA_signal_2150), 
        .A2(new_AGEMA_signal_1928), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_15_Q7), .A2(SubCellInst_SboxInst_15_Q6), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_n33), .Z(new_AGEMA_signal_2281) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n32), .B(
        SubCellInst_SboxInst_15_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_n30), .Z(new_AGEMA_signal_2280) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n29), .B(
        SubCellInst_SboxInst_15_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_n27), .Z(SubCellInst_SboxInst_15_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n26), .B(
        SubCellInst_SboxInst_15_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1928), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_1929), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L0), .B(SubCellInst_SboxInst_15_L2), .Z(
        SubCellInst_SboxInst_15_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2346), 
        .B(new_AGEMA_signal_1930), .Z(new_AGEMA_signal_2432) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2347), 
        .B(new_AGEMA_signal_1931), .Z(new_AGEMA_signal_2433) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L0), .B(SubCellInst_SboxInst_15_T3), .Z(
        SubCellOutput[60]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2346), .B(new_AGEMA_signal_2280), .Z(new_AGEMA_signal_2434) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2347), .B(new_AGEMA_signal_2281), .Z(new_AGEMA_signal_2435) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_15_YY_1_), .B(SubCellInst_SboxInst_15_YY_3), .ZN(
        SubCellOutput[61]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2344), .B(new_AGEMA_signal_2432), .Z(
        new_AGEMA_signal_2518) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_2345), .B(new_AGEMA_signal_2433), .Z(
        new_AGEMA_signal_2519) );
  INV_X1 AddConstXOR_U2_U1 ( .A(SubCellOutput_29), .ZN(ShiftRowsOutput[21]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_0_n1), .B(FSMUpdate[1]), .ZN(
        AddRoundConstantOutput[60]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2520), .B(1'b0), .Z(new_AGEMA_signal_2596) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2521), .B(1'b0), .Z(new_AGEMA_signal_2597) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[60]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_0_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2434), .Z(new_AGEMA_signal_2520) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2435), .Z(new_AGEMA_signal_2521) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_1_n1), .B(FSM_1), .ZN(
        AddRoundConstantOutput[61]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2598), .B(1'b0), .Z(new_AGEMA_signal_2730) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2599), .B(1'b0), .Z(new_AGEMA_signal_2731) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[61]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_1_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2518), .Z(new_AGEMA_signal_2598) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2519), .Z(new_AGEMA_signal_2599) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_0_n1), .B(FSM[4]), .ZN(
        AddRoundConstantOutput[44]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2524), .B(1'b0), .Z(new_AGEMA_signal_2600) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2525), .B(1'b0), .Z(new_AGEMA_signal_2601) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_44), .ZN(AddConstXOR_AddConstXOR_XORInst_1_0_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2418), .Z(new_AGEMA_signal_2524) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2419), .Z(new_AGEMA_signal_2525) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_1_n1), .B(FSM[5]), .ZN(
        AddRoundConstantOutput[45]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2602), .B(1'b0), .Z(new_AGEMA_signal_2732) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2603), .B(1'b0), .Z(new_AGEMA_signal_2733) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_45), .ZN(AddConstXOR_AddConstXOR_XORInst_1_1_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2510), .Z(new_AGEMA_signal_2602) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2511), .Z(new_AGEMA_signal_2603) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_0_n1), .B(
        TweakeyGeneration_key_Feedback[0]), .ZN(ShiftRowsOutput[44]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2528), .B(new_AGEMA_signal_1356), .Z(
        new_AGEMA_signal_2604) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2529), .B(new_AGEMA_signal_1357), .Z(
        new_AGEMA_signal_2605) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[32]), .ZN(AddRoundTweakeyXOR_XORInst_0_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2406), .Z(new_AGEMA_signal_2528) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2407), .Z(new_AGEMA_signal_2529) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_1_n1), .B(
        TweakeyGeneration_key_Feedback[1]), .ZN(ShiftRowsOutput[45]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2606), .B(new_AGEMA_signal_1362), .Z(
        new_AGEMA_signal_2734) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2607), .B(new_AGEMA_signal_1363), .Z(
        new_AGEMA_signal_2735) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[33]), .ZN(AddRoundTweakeyXOR_XORInst_0_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2504), .Z(new_AGEMA_signal_2606) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2505), .Z(new_AGEMA_signal_2607) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_0_n1), .B(
        TweakeyGeneration_key_Feedback[4]), .ZN(ShiftRowsOutput[32]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2532), .B(new_AGEMA_signal_1380), .Z(
        new_AGEMA_signal_2608) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2533), .B(new_AGEMA_signal_1381), .Z(
        new_AGEMA_signal_2609) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[36]), .ZN(AddRoundTweakeyXOR_XORInst_1_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2410), .Z(new_AGEMA_signal_2532) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2411), .Z(new_AGEMA_signal_2533) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_1_n1), .B(
        TweakeyGeneration_key_Feedback[5]), .ZN(ShiftRowsOutput[33]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2610), .B(new_AGEMA_signal_1386), .Z(
        new_AGEMA_signal_2736) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2611), .B(new_AGEMA_signal_1387), .Z(
        new_AGEMA_signal_2737) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[37]), .ZN(AddRoundTweakeyXOR_XORInst_1_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2506), .Z(new_AGEMA_signal_2610) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2507), .Z(new_AGEMA_signal_2611) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_0_n1), .B(
        TweakeyGeneration_key_Feedback[8]), .ZN(ShiftRowsOutput[36]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2536), .B(new_AGEMA_signal_1404), .Z(
        new_AGEMA_signal_2612) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2537), .B(new_AGEMA_signal_1405), .Z(
        new_AGEMA_signal_2613) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[40]), .ZN(AddRoundTweakeyXOR_XORInst_2_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2414), .Z(new_AGEMA_signal_2536) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2415), .Z(new_AGEMA_signal_2537) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_1_n1), .B(
        TweakeyGeneration_key_Feedback[9]), .ZN(ShiftRowsOutput[37]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2614), .B(new_AGEMA_signal_1410), .Z(
        new_AGEMA_signal_2738) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2615), .B(new_AGEMA_signal_1411), .Z(
        new_AGEMA_signal_2739) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[41]), .ZN(AddRoundTweakeyXOR_XORInst_2_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2508), .Z(new_AGEMA_signal_2614) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2509), .Z(new_AGEMA_signal_2615) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_0_n1), .B(
        TweakeyGeneration_key_Feedback[12]), .ZN(ShiftRowsOutput[40]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2740), .B(new_AGEMA_signal_1428), .Z(
        new_AGEMA_signal_2850) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2741), .B(new_AGEMA_signal_1429), .Z(
        new_AGEMA_signal_2851) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[44]), .ZN(AddRoundTweakeyXOR_XORInst_3_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2600), .Z(new_AGEMA_signal_2740) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2601), .Z(new_AGEMA_signal_2741) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_1_n1), .B(
        TweakeyGeneration_key_Feedback[13]), .ZN(ShiftRowsOutput[41]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2852), .B(new_AGEMA_signal_1434), .Z(
        new_AGEMA_signal_2958) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2853), .B(new_AGEMA_signal_1435), .Z(
        new_AGEMA_signal_2959) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[45]), .ZN(AddRoundTweakeyXOR_XORInst_3_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2732), .Z(new_AGEMA_signal_2852) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2733), .Z(new_AGEMA_signal_2853) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_0_n1), .B(
        TweakeyGeneration_key_Feedback[16]), .ZN(MCOutput[32]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2542), .B(new_AGEMA_signal_1452), .Z(
        new_AGEMA_signal_2620) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2543), .B(new_AGEMA_signal_1453), .Z(
        new_AGEMA_signal_2621) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[48]), .ZN(AddRoundTweakeyXOR_XORInst_4_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2422), .Z(new_AGEMA_signal_2542) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2423), .Z(new_AGEMA_signal_2543) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_1_n1), .B(
        TweakeyGeneration_key_Feedback[17]), .ZN(MCOutput[33]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2622), .B(new_AGEMA_signal_1458), .Z(
        new_AGEMA_signal_2744) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2623), .B(new_AGEMA_signal_1459), .Z(
        new_AGEMA_signal_2745) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[49]), .ZN(AddRoundTweakeyXOR_XORInst_4_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2512), .Z(new_AGEMA_signal_2622) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2513), .Z(new_AGEMA_signal_2623) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_0_n1), .B(
        TweakeyGeneration_key_Feedback[20]), .ZN(MCOutput[36]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2546), .B(new_AGEMA_signal_1476), .Z(
        new_AGEMA_signal_2624) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2547), .B(new_AGEMA_signal_1477), .Z(
        new_AGEMA_signal_2625) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[52]), .ZN(AddRoundTweakeyXOR_XORInst_5_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2426), .Z(new_AGEMA_signal_2546) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2427), .Z(new_AGEMA_signal_2547) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_1_n1), .B(
        TweakeyGeneration_key_Feedback[21]), .ZN(MCOutput[37]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2626), .B(new_AGEMA_signal_1482), .Z(
        new_AGEMA_signal_2746) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2627), .B(new_AGEMA_signal_1483), .Z(
        new_AGEMA_signal_2747) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[53]), .ZN(AddRoundTweakeyXOR_XORInst_5_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2514), .Z(new_AGEMA_signal_2626) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2515), .Z(new_AGEMA_signal_2627) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_0_n1), .B(
        TweakeyGeneration_key_Feedback[24]), .ZN(MCOutput[40]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2550), .B(new_AGEMA_signal_1500), .Z(
        new_AGEMA_signal_2628) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2551), .B(new_AGEMA_signal_1501), .Z(
        new_AGEMA_signal_2629) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[56]), .ZN(AddRoundTweakeyXOR_XORInst_6_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2430), .Z(new_AGEMA_signal_2550) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2431), .Z(new_AGEMA_signal_2551) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_1_n1), .B(
        TweakeyGeneration_key_Feedback[25]), .ZN(MCOutput[41]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2630), .B(new_AGEMA_signal_1506), .Z(
        new_AGEMA_signal_2748) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2631), .B(new_AGEMA_signal_1507), .Z(
        new_AGEMA_signal_2749) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[57]), .ZN(AddRoundTweakeyXOR_XORInst_6_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2516), .Z(new_AGEMA_signal_2630) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2517), .Z(new_AGEMA_signal_2631) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_0_n1), .B(
        TweakeyGeneration_key_Feedback[28]), .ZN(MCOutput[44]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2750), .B(new_AGEMA_signal_1524), .Z(
        new_AGEMA_signal_2854) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2751), .B(new_AGEMA_signal_1525), .Z(
        new_AGEMA_signal_2855) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[60]), .ZN(AddRoundTweakeyXOR_XORInst_7_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2596), .Z(new_AGEMA_signal_2750) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2597), .Z(new_AGEMA_signal_2751) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_1_n1), .B(
        TweakeyGeneration_key_Feedback[29]), .ZN(MCOutput[45]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2856), .B(new_AGEMA_signal_1530), .Z(
        new_AGEMA_signal_2960) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2857), .B(new_AGEMA_signal_1531), .Z(
        new_AGEMA_signal_2961) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[61]), .ZN(AddRoundTweakeyXOR_XORInst_7_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2730), .Z(new_AGEMA_signal_2856) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2731), .Z(new_AGEMA_signal_2857) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_0_n2), 
        .B(MCInst_MCR0_XORInst_0_0_n1), .ZN(MCOutput[48]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2754), .B(
        new_AGEMA_signal_2556), .Z(new_AGEMA_signal_2858) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2755), .B(
        new_AGEMA_signal_2557), .Z(new_AGEMA_signal_2859) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[16]), .B(
        ShiftRowsOutput[0]), .ZN(MCInst_MCR0_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2398), .B(
        new_AGEMA_signal_2386), .Z(new_AGEMA_signal_2556) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2399), .B(
        new_AGEMA_signal_2387), .Z(new_AGEMA_signal_2557) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[32]), 
        .Z(MCInst_MCR0_XORInst_0_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2620), .Z(new_AGEMA_signal_2754) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2621), .Z(new_AGEMA_signal_2755) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_1_n2), 
        .B(MCInst_MCR0_XORInst_0_1_n1), .ZN(MCOutput[49]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2860), .B(
        new_AGEMA_signal_2636), .Z(new_AGEMA_signal_2962) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2861), .B(
        new_AGEMA_signal_2637), .Z(new_AGEMA_signal_2963) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[17]), .B(
        ShiftRowsOutput[1]), .ZN(MCInst_MCR0_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2500), .B(
        new_AGEMA_signal_2494), .Z(new_AGEMA_signal_2636) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2501), .B(
        new_AGEMA_signal_2495), .Z(new_AGEMA_signal_2637) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[33]), 
        .Z(MCInst_MCR0_XORInst_0_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2744), .Z(new_AGEMA_signal_2860) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2745), .Z(new_AGEMA_signal_2861) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_0_n2), 
        .B(MCInst_MCR0_XORInst_1_0_n1), .ZN(MCOutput[52]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2758), .B(
        new_AGEMA_signal_2560), .Z(new_AGEMA_signal_2862) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2759), .B(
        new_AGEMA_signal_2561), .Z(new_AGEMA_signal_2863) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[20]), .B(
        ShiftRowsOutput[4]), .ZN(MCInst_MCR0_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2402), .B(
        new_AGEMA_signal_2374), .Z(new_AGEMA_signal_2560) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2403), .B(
        new_AGEMA_signal_2375), .Z(new_AGEMA_signal_2561) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[36]), 
        .Z(MCInst_MCR0_XORInst_1_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2624), .Z(new_AGEMA_signal_2758) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2625), .Z(new_AGEMA_signal_2759) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_1_n2), 
        .B(MCInst_MCR0_XORInst_1_1_n1), .ZN(MCOutput[53]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2864), .B(
        new_AGEMA_signal_2760), .Z(new_AGEMA_signal_2964) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2865), .B(
        new_AGEMA_signal_2761), .Z(new_AGEMA_signal_2965) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[21]), .B(
        ShiftRowsOutput[5]), .ZN(MCInst_MCR0_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2594), .B(
        new_AGEMA_signal_2488), .Z(new_AGEMA_signal_2760) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2595), .B(
        new_AGEMA_signal_2489), .Z(new_AGEMA_signal_2761) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[37]), 
        .Z(MCInst_MCR0_XORInst_1_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2746), .Z(new_AGEMA_signal_2864) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2747), .Z(new_AGEMA_signal_2865) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_0_n2), 
        .B(MCInst_MCR0_XORInst_2_0_n1), .ZN(MCOutput[56]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2764), .B(
        new_AGEMA_signal_2564), .Z(new_AGEMA_signal_2866) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2765), .B(
        new_AGEMA_signal_2565), .Z(new_AGEMA_signal_2867) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[24]), .B(
        ShiftRowsOutput[8]), .ZN(MCInst_MCR0_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2390), .B(
        new_AGEMA_signal_2378), .Z(new_AGEMA_signal_2564) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2391), .B(
        new_AGEMA_signal_2379), .Z(new_AGEMA_signal_2565) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[40]), 
        .Z(MCInst_MCR0_XORInst_2_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2628), .Z(new_AGEMA_signal_2764) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2629), .Z(new_AGEMA_signal_2765) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_1_n2), 
        .B(MCInst_MCR0_XORInst_2_1_n1), .ZN(MCOutput[57]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2868), .B(
        new_AGEMA_signal_2646), .Z(new_AGEMA_signal_2966) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2869), .B(
        new_AGEMA_signal_2647), .Z(new_AGEMA_signal_2967) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[25]), .B(
        ShiftRowsOutput[9]), .ZN(MCInst_MCR0_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2496), .B(
        new_AGEMA_signal_2490), .Z(new_AGEMA_signal_2646) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2497), .B(
        new_AGEMA_signal_2491), .Z(new_AGEMA_signal_2647) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[41]), 
        .Z(MCInst_MCR0_XORInst_2_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2748), .Z(new_AGEMA_signal_2868) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2749), .Z(new_AGEMA_signal_2869) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_0_n2), 
        .B(MCInst_MCR0_XORInst_3_0_n1), .ZN(MCOutput[60]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2968), .B(
        new_AGEMA_signal_2568), .Z(new_AGEMA_signal_3044) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2969), .B(
        new_AGEMA_signal_2569), .Z(new_AGEMA_signal_3045) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[28]), .B(
        ShiftRowsOutput[12]), .ZN(MCInst_MCR0_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2394), .B(
        new_AGEMA_signal_2382), .Z(new_AGEMA_signal_2568) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2395), .B(
        new_AGEMA_signal_2383), .Z(new_AGEMA_signal_2569) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[44]), 
        .Z(MCInst_MCR0_XORInst_3_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2854), .Z(new_AGEMA_signal_2968) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2855), .Z(new_AGEMA_signal_2969) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_1_n2), 
        .B(MCInst_MCR0_XORInst_3_1_n1), .ZN(MCOutput[61]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3046), .B(
        new_AGEMA_signal_2652), .Z(new_AGEMA_signal_3068) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3047), .B(
        new_AGEMA_signal_2653), .Z(new_AGEMA_signal_3069) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[29]), .B(
        ShiftRowsOutput[13]), .ZN(MCInst_MCR0_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2498), .B(
        new_AGEMA_signal_2492), .Z(new_AGEMA_signal_2652) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2499), .B(
        new_AGEMA_signal_2493), .Z(new_AGEMA_signal_2653) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[45]), 
        .Z(MCInst_MCR0_XORInst_3_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2960), .Z(new_AGEMA_signal_3046) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2961), .Z(new_AGEMA_signal_3047) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_0_n1), 
        .B(ShiftRowsOutput[16]), .ZN(MCOutput[16]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2770), .B(
        new_AGEMA_signal_2398), .Z(new_AGEMA_signal_2874) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2771), .B(
        new_AGEMA_signal_2399), .Z(new_AGEMA_signal_2875) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[32]), .ZN(MCInst_MCR2_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2608), .Z(new_AGEMA_signal_2770) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2609), .Z(new_AGEMA_signal_2771) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_1_n1), 
        .B(ShiftRowsOutput[17]), .ZN(MCOutput[17]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2876), .B(
        new_AGEMA_signal_2500), .Z(new_AGEMA_signal_2972) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2877), .B(
        new_AGEMA_signal_2501), .Z(new_AGEMA_signal_2973) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[33]), .ZN(MCInst_MCR2_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2736), .Z(new_AGEMA_signal_2876) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2737), .Z(new_AGEMA_signal_2877) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_0_n1), 
        .B(ShiftRowsOutput[20]), .ZN(MCOutput[20]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2774), .B(
        new_AGEMA_signal_2402), .Z(new_AGEMA_signal_2878) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2775), .B(
        new_AGEMA_signal_2403), .Z(new_AGEMA_signal_2879) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[36]), .ZN(MCInst_MCR2_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2612), .Z(new_AGEMA_signal_2774) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2613), .Z(new_AGEMA_signal_2775) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_1_n1), 
        .B(ShiftRowsOutput[21]), .ZN(MCOutput[21]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2880), .B(
        new_AGEMA_signal_2594), .Z(new_AGEMA_signal_2974) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2881), .B(
        new_AGEMA_signal_2595), .Z(new_AGEMA_signal_2975) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[37]), .ZN(MCInst_MCR2_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2738), .Z(new_AGEMA_signal_2880) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2739), .Z(new_AGEMA_signal_2881) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_0_n1), 
        .B(ShiftRowsOutput[24]), .ZN(MCOutput[24]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2976), .B(
        new_AGEMA_signal_2390), .Z(new_AGEMA_signal_3048) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2977), .B(
        new_AGEMA_signal_2391), .Z(new_AGEMA_signal_3049) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[40]), .ZN(MCInst_MCR2_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2850), .Z(new_AGEMA_signal_2976) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2851), .Z(new_AGEMA_signal_2977) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_1_n1), 
        .B(ShiftRowsOutput[25]), .ZN(MCOutput[25]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3050), .B(
        new_AGEMA_signal_2496), .Z(new_AGEMA_signal_3070) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3051), .B(
        new_AGEMA_signal_2497), .Z(new_AGEMA_signal_3071) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[41]), .ZN(MCInst_MCR2_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2958), .Z(new_AGEMA_signal_3050) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2959), .Z(new_AGEMA_signal_3051) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_0_n1), 
        .B(ShiftRowsOutput[28]), .ZN(MCOutput[28]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2780), .B(
        new_AGEMA_signal_2394), .Z(new_AGEMA_signal_2886) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2781), .B(
        new_AGEMA_signal_2395), .Z(new_AGEMA_signal_2887) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[44]), .ZN(MCInst_MCR2_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2604), .Z(new_AGEMA_signal_2780) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2605), .Z(new_AGEMA_signal_2781) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_1_n1), 
        .B(ShiftRowsOutput[29]), .ZN(MCOutput[29]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2888), .B(
        new_AGEMA_signal_2498), .Z(new_AGEMA_signal_2980) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2889), .B(
        new_AGEMA_signal_2499), .Z(new_AGEMA_signal_2981) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[45]), .ZN(MCInst_MCR2_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2734), .Z(new_AGEMA_signal_2888) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2735), .Z(new_AGEMA_signal_2889) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_0_n1), 
        .B(ShiftRowsOutput[16]), .ZN(MCOutput[0]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2784), .B(
        new_AGEMA_signal_2398), .Z(new_AGEMA_signal_2890) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2785), .B(
        new_AGEMA_signal_2399), .Z(new_AGEMA_signal_2891) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[32]), 
        .ZN(MCInst_MCR3_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2620), .Z(new_AGEMA_signal_2784) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2621), .Z(new_AGEMA_signal_2785) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_1_n1), 
        .B(ShiftRowsOutput[17]), .ZN(MCOutput[1]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2892), .B(
        new_AGEMA_signal_2500), .Z(new_AGEMA_signal_2982) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2893), .B(
        new_AGEMA_signal_2501), .Z(new_AGEMA_signal_2983) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[33]), 
        .ZN(MCInst_MCR3_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2744), .Z(new_AGEMA_signal_2892) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2745), .Z(new_AGEMA_signal_2893) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_0_n1), 
        .B(ShiftRowsOutput[20]), .ZN(MCOutput[4]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2788), .B(
        new_AGEMA_signal_2402), .Z(new_AGEMA_signal_2894) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2789), .B(
        new_AGEMA_signal_2403), .Z(new_AGEMA_signal_2895) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[36]), 
        .ZN(MCInst_MCR3_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2624), .Z(new_AGEMA_signal_2788) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2625), .Z(new_AGEMA_signal_2789) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_1_n1), 
        .B(ShiftRowsOutput[21]), .ZN(MCOutput[5]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2896), .B(
        new_AGEMA_signal_2594), .Z(new_AGEMA_signal_2984) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2897), .B(
        new_AGEMA_signal_2595), .Z(new_AGEMA_signal_2985) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[37]), 
        .ZN(MCInst_MCR3_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2746), .Z(new_AGEMA_signal_2896) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2747), .Z(new_AGEMA_signal_2897) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_0_n1), 
        .B(ShiftRowsOutput[24]), .ZN(MCOutput[8]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2792), .B(
        new_AGEMA_signal_2390), .Z(new_AGEMA_signal_2898) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2793), .B(
        new_AGEMA_signal_2391), .Z(new_AGEMA_signal_2899) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[40]), 
        .ZN(MCInst_MCR3_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2628), .Z(new_AGEMA_signal_2792) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2629), .Z(new_AGEMA_signal_2793) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_1_n1), 
        .B(ShiftRowsOutput[25]), .ZN(MCOutput[9]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2900), .B(
        new_AGEMA_signal_2496), .Z(new_AGEMA_signal_2986) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2901), .B(
        new_AGEMA_signal_2497), .Z(new_AGEMA_signal_2987) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[41]), 
        .ZN(MCInst_MCR3_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2748), .Z(new_AGEMA_signal_2900) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2749), .Z(new_AGEMA_signal_2901) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_0_n1), 
        .B(ShiftRowsOutput[28]), .ZN(MCOutput[12]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2988), .B(
        new_AGEMA_signal_2394), .Z(new_AGEMA_signal_3052) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2989), .B(
        new_AGEMA_signal_2395), .Z(new_AGEMA_signal_3053) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[44]), 
        .ZN(MCInst_MCR3_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2854), .Z(new_AGEMA_signal_2988) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2855), .Z(new_AGEMA_signal_2989) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_1_n1), 
        .B(ShiftRowsOutput[29]), .ZN(MCOutput[13]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3054), .B(
        new_AGEMA_signal_2498), .Z(new_AGEMA_signal_3072) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3055), .B(
        new_AGEMA_signal_2499), .Z(new_AGEMA_signal_3073) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[45]), 
        .ZN(MCInst_MCR3_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2960), .Z(new_AGEMA_signal_3054) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2961), .Z(new_AGEMA_signal_3055) );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[63]), .CK(clk_gated), .Q(Ciphertext_s0[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3042), .CK(clk_gated), .Q(Ciphertext_s1[63]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3043), .CK(clk_gated), .Q(Ciphertext_s2[63]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[62]), .CK(clk_gated), .Q(Ciphertext_s0[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2956), .CK(clk_gated), .Q(Ciphertext_s1[62]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2957), .CK(clk_gated), .Q(Ciphertext_s2[62]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[61]), .CK(clk_gated), .Q(Ciphertext_s0[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3084), .CK(clk_gated), .Q(Ciphertext_s1[61]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3085), .CK(clk_gated), .Q(Ciphertext_s2[61]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[60]), .CK(clk_gated), .Q(Ciphertext_s0[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3066), .CK(clk_gated), .Q(Ciphertext_s1[60]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3067), .CK(clk_gated), .Q(Ciphertext_s2[60]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[59]), .CK(clk_gated), .Q(Ciphertext_s0[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2848), .CK(clk_gated), .Q(Ciphertext_s1[59]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2849), .CK(clk_gated), .Q(Ciphertext_s2[59]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[58]), .CK(clk_gated), .Q(Ciphertext_s0[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2728), .CK(clk_gated), .Q(Ciphertext_s1[58]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2729), .CK(clk_gated), .Q(Ciphertext_s2[58]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[57]), .CK(clk_gated), .Q(Ciphertext_s0[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3038), .CK(clk_gated), .Q(Ciphertext_s1[57]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3039), .CK(clk_gated), .Q(Ciphertext_s2[57]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[56]), .CK(clk_gated), .Q(Ciphertext_s0[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2952), .CK(clk_gated), .Q(Ciphertext_s1[56]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2953), .CK(clk_gated), .Q(Ciphertext_s2[56]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[55]), .CK(clk_gated), .Q(Ciphertext_s0[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2844), .CK(clk_gated), .Q(Ciphertext_s1[55]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2845), .CK(clk_gated), .Q(Ciphertext_s2[55]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[54]), .CK(clk_gated), .Q(Ciphertext_s0[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2724), .CK(clk_gated), .Q(Ciphertext_s1[54]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2725), .CK(clk_gated), .Q(Ciphertext_s2[54]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[53]), .CK(clk_gated), .Q(Ciphertext_s0[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3034), .CK(clk_gated), .Q(Ciphertext_s1[53]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3035), .CK(clk_gated), .Q(Ciphertext_s2[53]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[52]), .CK(clk_gated), .Q(Ciphertext_s0[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2948), .CK(clk_gated), .Q(Ciphertext_s1[52]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2949), .CK(clk_gated), .Q(Ciphertext_s2[52]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[51]), .CK(clk_gated), .Q(Ciphertext_s0[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2840), .CK(clk_gated), .Q(Ciphertext_s1[51]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2841), .CK(clk_gated), .Q(Ciphertext_s2[51]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[50]), .CK(clk_gated), .Q(Ciphertext_s0[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2720), .CK(clk_gated), .Q(Ciphertext_s1[50]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2721), .CK(clk_gated), .Q(Ciphertext_s2[50]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[49]), .CK(clk_gated), .Q(Ciphertext_s0[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3030), .CK(clk_gated), .Q(Ciphertext_s1[49]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3031), .CK(clk_gated), .Q(Ciphertext_s2[49]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[48]), .CK(clk_gated), .Q(Ciphertext_s0[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2944), .CK(clk_gated), .Q(Ciphertext_s1[48]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2945), .CK(clk_gated), .Q(Ciphertext_s2[48]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[47]), .CK(clk_gated), .Q(Ciphertext_s0[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2836), .CK(clk_gated), .Q(Ciphertext_s1[47]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2837), .CK(clk_gated), .Q(Ciphertext_s2[47]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[46]), .CK(clk_gated), .Q(Ciphertext_s0[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2716), .CK(clk_gated), .Q(Ciphertext_s1[46]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2717), .CK(clk_gated), .Q(Ciphertext_s2[46]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[45]), .CK(clk_gated), .Q(Ciphertext_s0[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3026), .CK(clk_gated), .Q(Ciphertext_s1[45]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3027), .CK(clk_gated), .Q(Ciphertext_s2[45]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[44]), .CK(clk_gated), .Q(Ciphertext_s0[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2940), .CK(clk_gated), .Q(Ciphertext_s1[44]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2941), .CK(clk_gated), .Q(Ciphertext_s2[44]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[43]), .CK(clk_gated), .Q(Ciphertext_s0[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2592), .CK(clk_gated), .Q(Ciphertext_s1[43]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2593), .CK(clk_gated), .Q(Ciphertext_s2[43]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[42]), .CK(clk_gated), .Q(Ciphertext_s0[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2486), .CK(clk_gated), .Q(Ciphertext_s1[42]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2487), .CK(clk_gated), .Q(Ciphertext_s2[42]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[41]), .CK(clk_gated), .Q(Ciphertext_s0[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2832), .CK(clk_gated), .Q(Ciphertext_s1[41]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2833), .CK(clk_gated), .Q(Ciphertext_s2[41]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[40]), .CK(clk_gated), .Q(Ciphertext_s0[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2712), .CK(clk_gated), .Q(Ciphertext_s1[40]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2713), .CK(clk_gated), .Q(Ciphertext_s2[40]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[39]), .CK(clk_gated), .Q(Ciphertext_s0[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2588), .CK(clk_gated), .Q(Ciphertext_s1[39]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2589), .CK(clk_gated), .Q(Ciphertext_s2[39]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[38]), .CK(clk_gated), .Q(Ciphertext_s0[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2482), .CK(clk_gated), .Q(Ciphertext_s1[38]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2483), .CK(clk_gated), .Q(Ciphertext_s2[38]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[37]), .CK(clk_gated), .Q(Ciphertext_s0[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2828), .CK(clk_gated), .Q(Ciphertext_s1[37]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2829), .CK(clk_gated), .Q(Ciphertext_s2[37]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[36]), .CK(clk_gated), .Q(Ciphertext_s0[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2708), .CK(clk_gated), .Q(Ciphertext_s1[36]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2709), .CK(clk_gated), .Q(Ciphertext_s2[36]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[35]), .CK(clk_gated), .Q(Ciphertext_s0[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2584), .CK(clk_gated), .Q(Ciphertext_s1[35]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2585), .CK(clk_gated), .Q(Ciphertext_s2[35]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[34]), .CK(clk_gated), .Q(Ciphertext_s0[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2478), .CK(clk_gated), .Q(Ciphertext_s1[34]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2479), .CK(clk_gated), .Q(Ciphertext_s2[34]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[33]), .CK(clk_gated), .Q(Ciphertext_s0[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2824), .CK(clk_gated), .Q(Ciphertext_s1[33]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2825), .CK(clk_gated), .Q(Ciphertext_s2[33]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[32]), .CK(clk_gated), .Q(Ciphertext_s0[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2704), .CK(clk_gated), .Q(Ciphertext_s1[32]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2705), .CK(clk_gated), .Q(Ciphertext_s2[32]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[31]), .CK(clk_gated), .Q(Ciphertext_s0[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2820), .CK(clk_gated), .Q(Ciphertext_s1[31]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2821), .CK(clk_gated), .Q(Ciphertext_s2[31]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[30]), .CK(clk_gated), .Q(Ciphertext_s0[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2700), .CK(clk_gated), .Q(Ciphertext_s1[30]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2701), .CK(clk_gated), .Q(Ciphertext_s2[30]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[29]), .CK(clk_gated), .Q(Ciphertext_s0[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3022), .CK(clk_gated), .Q(Ciphertext_s1[29]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3023), .CK(clk_gated), .Q(Ciphertext_s2[29]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[28]), .CK(clk_gated), .Q(Ciphertext_s0[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2936), .CK(clk_gated), .Q(Ciphertext_s1[28]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2937), .CK(clk_gated), .Q(Ciphertext_s2[28]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[27]), .CK(clk_gated), .Q(Ciphertext_s0[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3018), .CK(clk_gated), .Q(Ciphertext_s1[27]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3019), .CK(clk_gated), .Q(Ciphertext_s2[27]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[26]), .CK(clk_gated), .Q(Ciphertext_s0[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2932), .CK(clk_gated), .Q(Ciphertext_s1[26]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2933), .CK(clk_gated), .Q(Ciphertext_s2[26]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[25]), .CK(clk_gated), .Q(Ciphertext_s0[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3080), .CK(clk_gated), .Q(Ciphertext_s1[25]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3081), .CK(clk_gated), .Q(Ciphertext_s2[25]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[24]), .CK(clk_gated), .Q(Ciphertext_s0[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3062), .CK(clk_gated), .Q(Ciphertext_s1[24]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3063), .CK(clk_gated), .Q(Ciphertext_s2[24]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[23]), .CK(clk_gated), .Q(Ciphertext_s0[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2816), .CK(clk_gated), .Q(Ciphertext_s1[23]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2817), .CK(clk_gated), .Q(Ciphertext_s2[23]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[22]), .CK(clk_gated), .Q(Ciphertext_s0[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2696), .CK(clk_gated), .Q(Ciphertext_s1[22]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2697), .CK(clk_gated), .Q(Ciphertext_s2[22]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[21]), .CK(clk_gated), .Q(Ciphertext_s0[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3014), .CK(clk_gated), .Q(Ciphertext_s1[21]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3015), .CK(clk_gated), .Q(Ciphertext_s2[21]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[20]), .CK(clk_gated), .Q(Ciphertext_s0[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2928), .CK(clk_gated), .Q(Ciphertext_s1[20]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2929), .CK(clk_gated), .Q(Ciphertext_s2[20]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[19]), .CK(clk_gated), .Q(Ciphertext_s0[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2812), .CK(clk_gated), .Q(Ciphertext_s1[19]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2813), .CK(clk_gated), .Q(Ciphertext_s2[19]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[18]), .CK(clk_gated), .Q(Ciphertext_s0[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2692), .CK(clk_gated), .Q(Ciphertext_s1[18]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2693), .CK(clk_gated), .Q(Ciphertext_s2[18]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[17]), .CK(clk_gated), .Q(Ciphertext_s0[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3010), .CK(clk_gated), .Q(Ciphertext_s1[17]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3011), .CK(clk_gated), .Q(Ciphertext_s2[17]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[16]), .CK(clk_gated), .Q(Ciphertext_s0[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2924), .CK(clk_gated), .Q(Ciphertext_s1[16]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2925), .CK(clk_gated), .Q(Ciphertext_s2[16]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[15]), .CK(clk_gated), .Q(Ciphertext_s0[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3006), .CK(clk_gated), .Q(Ciphertext_s1[15]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3007), .CK(clk_gated), .Q(Ciphertext_s2[15]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[14]), .CK(clk_gated), .Q(Ciphertext_s0[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2920), .CK(clk_gated), .Q(Ciphertext_s1[14]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2921), .CK(clk_gated), .Q(Ciphertext_s2[14]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[13]), .CK(clk_gated), .Q(Ciphertext_s0[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3076), .CK(clk_gated), .Q(Ciphertext_s1[13]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3077), .CK(clk_gated), .Q(Ciphertext_s2[13]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[12]), .CK(clk_gated), .Q(Ciphertext_s0[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3058), .CK(clk_gated), .Q(Ciphertext_s1[12]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3059), .CK(clk_gated), .Q(Ciphertext_s2[12]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[11]), .CK(clk_gated), .Q(Ciphertext_s0[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2808), .CK(clk_gated), .Q(Ciphertext_s1[11]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2809), .CK(clk_gated), .Q(Ciphertext_s2[11]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[10]), .CK(clk_gated), .Q(Ciphertext_s0[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2688), .CK(clk_gated), .Q(Ciphertext_s1[10]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2689), .CK(clk_gated), .Q(Ciphertext_s2[10]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[9]), .CK(clk_gated), .Q(Ciphertext_s0[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3002), .CK(clk_gated), .Q(Ciphertext_s1[9]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3003), .CK(clk_gated), .Q(Ciphertext_s2[9]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[8]), .CK(clk_gated), .Q(Ciphertext_s0[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2916), .CK(clk_gated), .Q(Ciphertext_s1[8]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2917), .CK(clk_gated), .Q(Ciphertext_s2[8]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[7]), .CK(clk_gated), .Q(Ciphertext_s0[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2804), .CK(clk_gated), .Q(Ciphertext_s1[7]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2805), .CK(clk_gated), .Q(Ciphertext_s2[7]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[6]), .CK(clk_gated), .Q(Ciphertext_s0[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2684), .CK(clk_gated), .Q(Ciphertext_s1[6]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2685), .CK(clk_gated), .Q(Ciphertext_s2[6]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[5]), .CK(clk_gated), .Q(Ciphertext_s0[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2998), .CK(clk_gated), .Q(Ciphertext_s1[5]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2999), .CK(clk_gated), .Q(Ciphertext_s2[5]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[4]), .CK(clk_gated), .Q(Ciphertext_s0[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2912), .CK(clk_gated), .Q(Ciphertext_s1[4]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2913), .CK(clk_gated), .Q(Ciphertext_s2[4]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[3]), .CK(clk_gated), .Q(Ciphertext_s0[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2800), .CK(clk_gated), .Q(Ciphertext_s1[3]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2801), .CK(clk_gated), .Q(Ciphertext_s2[3]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[2]), .CK(clk_gated), .Q(Ciphertext_s0[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2680), .CK(clk_gated), .Q(Ciphertext_s1[2]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2681), .CK(clk_gated), .Q(Ciphertext_s2[2]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[1]), .CK(clk_gated), .Q(Ciphertext_s0[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2994), .CK(clk_gated), .Q(Ciphertext_s1[1]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2995), .CK(clk_gated), .Q(Ciphertext_s2[1]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[0]), .CK(clk_gated), .Q(Ciphertext_s0[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2908), .CK(clk_gated), .Q(Ciphertext_s1[0]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2909), .CK(clk_gated), .Q(Ciphertext_s2[0]), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[63]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[31]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1738), .CK(clk_gated), .Q(new_AGEMA_signal_1542), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1739), .CK(clk_gated), .Q(new_AGEMA_signal_1543), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[62]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[30]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1732), .CK(clk_gated), .Q(new_AGEMA_signal_1536), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1733), .CK(clk_gated), .Q(new_AGEMA_signal_1537), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[61]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[29]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1726), .CK(clk_gated), .Q(new_AGEMA_signal_1530), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1727), .CK(clk_gated), .Q(new_AGEMA_signal_1531), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[60]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[28]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1720), .CK(clk_gated), .Q(new_AGEMA_signal_1524), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1721), .CK(clk_gated), .Q(new_AGEMA_signal_1525), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[59]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[27]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1714), .CK(clk_gated), .Q(new_AGEMA_signal_1518), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1715), .CK(clk_gated), .Q(new_AGEMA_signal_1519), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[58]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[26]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1708), .CK(clk_gated), .Q(new_AGEMA_signal_1512), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1709), .CK(clk_gated), .Q(new_AGEMA_signal_1513), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[57]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[25]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1702), .CK(clk_gated), .Q(new_AGEMA_signal_1506), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1703), .CK(clk_gated), .Q(new_AGEMA_signal_1507), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[56]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[24]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1696), .CK(clk_gated), .Q(new_AGEMA_signal_1500), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1697), .CK(clk_gated), .Q(new_AGEMA_signal_1501), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[55]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[23]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1690), .CK(clk_gated), .Q(new_AGEMA_signal_1494), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1691), .CK(clk_gated), .Q(new_AGEMA_signal_1495), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[54]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[22]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1684), .CK(clk_gated), .Q(new_AGEMA_signal_1488), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1685), .CK(clk_gated), .Q(new_AGEMA_signal_1489), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[53]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[21]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1678), .CK(clk_gated), .Q(new_AGEMA_signal_1482), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1679), .CK(clk_gated), .Q(new_AGEMA_signal_1483), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[52]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[20]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1672), .CK(clk_gated), .Q(new_AGEMA_signal_1476), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1673), .CK(clk_gated), .Q(new_AGEMA_signal_1477), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[51]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[19]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1666), .CK(clk_gated), .Q(new_AGEMA_signal_1470), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1667), .CK(clk_gated), .Q(new_AGEMA_signal_1471), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[50]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[18]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1660), .CK(clk_gated), .Q(new_AGEMA_signal_1464), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1661), .CK(clk_gated), .Q(new_AGEMA_signal_1465), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[49]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[17]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1654), .CK(clk_gated), .Q(new_AGEMA_signal_1458), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1655), .CK(clk_gated), .Q(new_AGEMA_signal_1459), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[48]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[16]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1648), .CK(clk_gated), .Q(new_AGEMA_signal_1452), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1649), .CK(clk_gated), .Q(new_AGEMA_signal_1453), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[47]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[15]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1642), .CK(clk_gated), .Q(new_AGEMA_signal_1446), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1643), .CK(clk_gated), .Q(new_AGEMA_signal_1447), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[46]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[14]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1636), .CK(clk_gated), .Q(new_AGEMA_signal_1440), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1637), .CK(clk_gated), .Q(new_AGEMA_signal_1441), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[45]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[13]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1630), .CK(clk_gated), .Q(new_AGEMA_signal_1434), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1631), .CK(clk_gated), .Q(new_AGEMA_signal_1435), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[44]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[12]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1624), .CK(clk_gated), .Q(new_AGEMA_signal_1428), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1625), .CK(clk_gated), .Q(new_AGEMA_signal_1429), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[43]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[11]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1618), .CK(clk_gated), .Q(new_AGEMA_signal_1422), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1619), .CK(clk_gated), .Q(new_AGEMA_signal_1423), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[42]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[10]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1612), .CK(clk_gated), .Q(new_AGEMA_signal_1416), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1613), .CK(clk_gated), .Q(new_AGEMA_signal_1417), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[41]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[9]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1606), .CK(clk_gated), .Q(new_AGEMA_signal_1410), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1607), .CK(clk_gated), .Q(new_AGEMA_signal_1411), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[40]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[8]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1600), .CK(clk_gated), .Q(new_AGEMA_signal_1404), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1601), .CK(clk_gated), .Q(new_AGEMA_signal_1405), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[39]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[7]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1594), .CK(clk_gated), .Q(new_AGEMA_signal_1398), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1595), .CK(clk_gated), .Q(new_AGEMA_signal_1399), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[38]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[6]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1588), .CK(clk_gated), .Q(new_AGEMA_signal_1392), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1589), .CK(clk_gated), .Q(new_AGEMA_signal_1393), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[37]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[5]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1582), .CK(clk_gated), .Q(new_AGEMA_signal_1386), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1583), .CK(clk_gated), .Q(new_AGEMA_signal_1387), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[36]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[4]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1576), .CK(clk_gated), .Q(new_AGEMA_signal_1380), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1577), .CK(clk_gated), .Q(new_AGEMA_signal_1381), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[35]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[3]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1570), .CK(clk_gated), .Q(new_AGEMA_signal_1374), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1571), .CK(clk_gated), .Q(new_AGEMA_signal_1375), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[34]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[2]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1564), .CK(clk_gated), .Q(new_AGEMA_signal_1368), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1565), .CK(clk_gated), .Q(new_AGEMA_signal_1369), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[33]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[1]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1558), .CK(clk_gated), .Q(new_AGEMA_signal_1362), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1559), .CK(clk_gated), .Q(new_AGEMA_signal_1363), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[32]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[0]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1552), .CK(clk_gated), .Q(new_AGEMA_signal_1356), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1553), .CK(clk_gated), .Q(new_AGEMA_signal_1357), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[31]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[55]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1546), .CK(clk_gated), .Q(new_AGEMA_signal_1686), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1547), .CK(clk_gated), .Q(new_AGEMA_signal_1687), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[30]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[54]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1540), .CK(clk_gated), .Q(new_AGEMA_signal_1680), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1541), .CK(clk_gated), .Q(new_AGEMA_signal_1681), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[29]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[53]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1534), .CK(clk_gated), .Q(new_AGEMA_signal_1674), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1535), .CK(clk_gated), .Q(new_AGEMA_signal_1675), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[28]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[52]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1528), .CK(clk_gated), .Q(new_AGEMA_signal_1668), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1529), .CK(clk_gated), .Q(new_AGEMA_signal_1669), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[27]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[63]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1522), .CK(clk_gated), .Q(new_AGEMA_signal_1734), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1523), .CK(clk_gated), .Q(new_AGEMA_signal_1735), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[26]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[62]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1516), .CK(clk_gated), .Q(new_AGEMA_signal_1728), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1517), .CK(clk_gated), .Q(new_AGEMA_signal_1729), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[25]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[61]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1510), .CK(clk_gated), .Q(new_AGEMA_signal_1722), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1511), .CK(clk_gated), .Q(new_AGEMA_signal_1723), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[24]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[60]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1504), .CK(clk_gated), .Q(new_AGEMA_signal_1716), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1505), .CK(clk_gated), .Q(new_AGEMA_signal_1717), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[23]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[47]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1498), .CK(clk_gated), .Q(new_AGEMA_signal_1638), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1499), .CK(clk_gated), .Q(new_AGEMA_signal_1639), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[22]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[46]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1492), .CK(clk_gated), .Q(new_AGEMA_signal_1632), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1493), .CK(clk_gated), .Q(new_AGEMA_signal_1633), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[21]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[45]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1486), .CK(clk_gated), .Q(new_AGEMA_signal_1626), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1487), .CK(clk_gated), .Q(new_AGEMA_signal_1627), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[20]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[44]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1480), .CK(clk_gated), .Q(new_AGEMA_signal_1620), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1481), .CK(clk_gated), .Q(new_AGEMA_signal_1621), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[19]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[35]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1474), .CK(clk_gated), .Q(new_AGEMA_signal_1566), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1475), .CK(clk_gated), .Q(new_AGEMA_signal_1567), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[18]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[34]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1468), .CK(clk_gated), .Q(new_AGEMA_signal_1560), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1469), .CK(clk_gated), .Q(new_AGEMA_signal_1561), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[17]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[33]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1462), .CK(clk_gated), .Q(new_AGEMA_signal_1554), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1463), .CK(clk_gated), .Q(new_AGEMA_signal_1555), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[16]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[32]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1456), .CK(clk_gated), .Q(new_AGEMA_signal_1548), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1457), .CK(clk_gated), .Q(new_AGEMA_signal_1549), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[15]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[39]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1450), .CK(clk_gated), .Q(new_AGEMA_signal_1590), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1451), .CK(clk_gated), .Q(new_AGEMA_signal_1591), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[14]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[38]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1444), .CK(clk_gated), .Q(new_AGEMA_signal_1584), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1445), .CK(clk_gated), .Q(new_AGEMA_signal_1585), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[13]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[37]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1438), .CK(clk_gated), .Q(new_AGEMA_signal_1578), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1439), .CK(clk_gated), .Q(new_AGEMA_signal_1579), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[12]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[36]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1432), .CK(clk_gated), .Q(new_AGEMA_signal_1572), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1433), .CK(clk_gated), .Q(new_AGEMA_signal_1573), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[11]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[51]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1426), .CK(clk_gated), .Q(new_AGEMA_signal_1662), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1427), .CK(clk_gated), .Q(new_AGEMA_signal_1663), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[10]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[50]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1420), .CK(clk_gated), .Q(new_AGEMA_signal_1656), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1421), .CK(clk_gated), .Q(new_AGEMA_signal_1657), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[9]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[49]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1414), .CK(clk_gated), .Q(new_AGEMA_signal_1650), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1415), .CK(clk_gated), .Q(new_AGEMA_signal_1651), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[8]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[48]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1408), .CK(clk_gated), .Q(new_AGEMA_signal_1644), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1409), .CK(clk_gated), .Q(new_AGEMA_signal_1645), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[7]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[43]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1402), .CK(clk_gated), .Q(new_AGEMA_signal_1614), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1403), .CK(clk_gated), .Q(new_AGEMA_signal_1615), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[6]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[42]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1396), .CK(clk_gated), .Q(new_AGEMA_signal_1608), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1397), .CK(clk_gated), .Q(new_AGEMA_signal_1609), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[5]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[41]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1390), .CK(clk_gated), .Q(new_AGEMA_signal_1602), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1391), .CK(clk_gated), .Q(new_AGEMA_signal_1603), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[4]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[40]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1384), .CK(clk_gated), .Q(new_AGEMA_signal_1596), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1385), .CK(clk_gated), .Q(new_AGEMA_signal_1597), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[3]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[59]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1378), .CK(clk_gated), .Q(new_AGEMA_signal_1710), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1379), .CK(clk_gated), .Q(new_AGEMA_signal_1711), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[2]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[58]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1372), .CK(clk_gated), .Q(new_AGEMA_signal_1704), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1373), .CK(clk_gated), .Q(new_AGEMA_signal_1705), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[1]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[57]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1366), .CK(clk_gated), .Q(new_AGEMA_signal_1698), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1367), .CK(clk_gated), .Q(new_AGEMA_signal_1699), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[0]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[56]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1360), .CK(clk_gated), .Q(new_AGEMA_signal_1692), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_1361), .CK(clk_gated), .Q(new_AGEMA_signal_1693), 
        .QN() );
endmodule

