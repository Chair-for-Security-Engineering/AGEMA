/* modified netlist. Source: module LED in file ../CaseStudies/11_LED_round_based_encryption/netlists/LED.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module LED_LMDPL_Pipeline_d1 (IN_plaintext_s0, IN_key_s0, IN_reset, CLK, Po_rst, Fresh, IN_plaintext_s1, IN_key_s1, OUT_ciphertext_s0, OUT_done, OUT_ciphertext_s1);
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input IN_reset ;
    input CLK ;
    input Po_rst ;
    input [63:0] IN_plaintext_s1 ;
    input [127:0] IN_key_s1 ;
    input [63:0] Fresh ;
    output [63:0] OUT_ciphertext_s0 ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s1 ;
    wire n15 ;
    wire n14 ;
    wire n16 ;
    wire n17 ;
    wire n18 ;
    wire n19 ;
    wire n20 ;
    wire LED_128_Instance_n34 ;
    wire LED_128_Instance_n33 ;
    wire LED_128_Instance_n32 ;
    wire LED_128_Instance_n23 ;
    wire LED_128_Instance_n21 ;
    wire LED_128_Instance_n20 ;
    wire LED_128_Instance_n19 ;
    wire LED_128_Instance_n18 ;
    wire LED_128_Instance_n17 ;
    wire LED_128_Instance_n16 ;
    wire LED_128_Instance_n15 ;
    wire LED_128_Instance_n14 ;
    wire LED_128_Instance_n13 ;
    wire LED_128_Instance_n12 ;
    wire LED_128_Instance_n11 ;
    wire LED_128_Instance_n10 ;
    wire LED_128_Instance_n2 ;
    wire LED_128_Instance_n1 ;
    wire LED_128_Instance_n27 ;
    wire LED_128_Instance_N9 ;
    wire LED_128_Instance_n28 ;
    wire LED_128_Instance_N8 ;
    wire LED_128_Instance_n30 ;
    wire LED_128_Instance_N7 ;
    wire LED_128_Instance_n5 ;
    wire LED_128_Instance_N6 ;
    wire LED_128_Instance_n29 ;
    wire LED_128_Instance_N5 ;
    wire LED_128_Instance_n6 ;
    wire LED_128_Instance_N4 ;
    wire LED_128_Instance_n24 ;
    wire LED_128_Instance_N13 ;
    wire LED_128_Instance_n25 ;
    wire LED_128_Instance_N12 ;
    wire LED_128_Instance_n8 ;
    wire LED_128_Instance_n26 ;
    wire LED_128_Instance_N11 ;
    wire LED_128_Instance_n4 ;
    wire LED_128_Instance_N10 ;
    wire LED_128_Instance_n31 ;
    wire LED_128_Instance_addroundkey_out_0_ ;
    wire LED_128_Instance_addroundkey_out_1_ ;
    wire LED_128_Instance_addroundkey_out_2_ ;
    wire LED_128_Instance_addroundkey_out_3_ ;
    wire LED_128_Instance_addroundkey_out_4_ ;
    wire LED_128_Instance_addroundkey_out_5_ ;
    wire LED_128_Instance_addroundkey_out_6_ ;
    wire LED_128_Instance_addroundkey_out_16_ ;
    wire LED_128_Instance_addroundkey_out_17_ ;
    wire LED_128_Instance_addroundkey_out_18_ ;
    wire LED_128_Instance_addroundkey_out_19_ ;
    wire LED_128_Instance_addroundkey_out_20_ ;
    wire LED_128_Instance_addroundkey_out_21_ ;
    wire LED_128_Instance_addroundkey_out_22_ ;
    wire LED_128_Instance_addroundkey_out_32_ ;
    wire LED_128_Instance_addroundkey_out_33_ ;
    wire LED_128_Instance_addroundkey_out_34_ ;
    wire LED_128_Instance_addroundkey_out_35_ ;
    wire LED_128_Instance_addroundkey_out_36_ ;
    wire LED_128_Instance_addroundkey_out_37_ ;
    wire LED_128_Instance_addroundkey_out_38_ ;
    wire LED_128_Instance_addroundkey_out_48_ ;
    wire LED_128_Instance_addroundkey_out_49_ ;
    wire LED_128_Instance_addroundkey_out_50_ ;
    wire LED_128_Instance_addroundkey_out_51_ ;
    wire LED_128_Instance_addroundkey_out_52_ ;
    wire LED_128_Instance_addroundkey_out_53_ ;
    wire LED_128_Instance_addroundkey_out_54_ ;
    wire LED_128_Instance_n22 ;
    wire LED_128_Instance_MUX_state0_n11 ;
    wire LED_128_Instance_MUX_state0_n10 ;
    wire LED_128_Instance_MUX_state0_n9 ;
    wire LED_128_Instance_MUX_state0_n8 ;
    wire LED_128_Instance_MUX_current_roundkey_n10 ;
    wire LED_128_Instance_MUX_current_roundkey_n9 ;
    wire LED_128_Instance_MUX_current_roundkey_n8 ;
    wire LED_128_Instance_MUX_current_roundkey_n7 ;
    wire LED_128_Instance_MUX_addroundkey_out_n9 ;
    wire LED_128_Instance_MUX_addroundkey_out_n8 ;
    wire LED_128_Instance_MUX_addroundkey_out_n7 ;
    wire LED_128_Instance_SBox_Instance_0_n3 ;
    wire LED_128_Instance_SBox_Instance_0_n2 ;
    wire LED_128_Instance_SBox_Instance_0_n1 ;
    wire LED_128_Instance_SBox_Instance_0_L8 ;
    wire LED_128_Instance_SBox_Instance_0_L7 ;
    wire LED_128_Instance_SBox_Instance_0_T3 ;
    wire LED_128_Instance_SBox_Instance_0_T1 ;
    wire LED_128_Instance_SBox_Instance_0_Q7 ;
    wire LED_128_Instance_SBox_Instance_0_Q6 ;
    wire LED_128_Instance_SBox_Instance_0_L5 ;
    wire LED_128_Instance_SBox_Instance_0_T2 ;
    wire LED_128_Instance_SBox_Instance_0_L4 ;
    wire LED_128_Instance_SBox_Instance_0_Q3 ;
    wire LED_128_Instance_SBox_Instance_0_L3 ;
    wire LED_128_Instance_SBox_Instance_0_Q2 ;
    wire LED_128_Instance_SBox_Instance_0_T0 ;
    wire LED_128_Instance_SBox_Instance_0_L2 ;
    wire LED_128_Instance_SBox_Instance_0_L1 ;
    wire LED_128_Instance_SBox_Instance_0_L0 ;
    wire LED_128_Instance_SBox_Instance_1_n3 ;
    wire LED_128_Instance_SBox_Instance_1_n2 ;
    wire LED_128_Instance_SBox_Instance_1_n1 ;
    wire LED_128_Instance_SBox_Instance_1_L8 ;
    wire LED_128_Instance_SBox_Instance_1_L7 ;
    wire LED_128_Instance_SBox_Instance_1_T3 ;
    wire LED_128_Instance_SBox_Instance_1_T1 ;
    wire LED_128_Instance_SBox_Instance_1_Q7 ;
    wire LED_128_Instance_SBox_Instance_1_Q6 ;
    wire LED_128_Instance_SBox_Instance_1_L5 ;
    wire LED_128_Instance_SBox_Instance_1_T2 ;
    wire LED_128_Instance_SBox_Instance_1_L4 ;
    wire LED_128_Instance_SBox_Instance_1_Q3 ;
    wire LED_128_Instance_SBox_Instance_1_L3 ;
    wire LED_128_Instance_SBox_Instance_1_Q2 ;
    wire LED_128_Instance_SBox_Instance_1_T0 ;
    wire LED_128_Instance_SBox_Instance_1_L2 ;
    wire LED_128_Instance_SBox_Instance_1_L1 ;
    wire LED_128_Instance_SBox_Instance_1_L0 ;
    wire LED_128_Instance_SBox_Instance_2_n3 ;
    wire LED_128_Instance_SBox_Instance_2_n2 ;
    wire LED_128_Instance_SBox_Instance_2_n1 ;
    wire LED_128_Instance_SBox_Instance_2_L8 ;
    wire LED_128_Instance_SBox_Instance_2_L7 ;
    wire LED_128_Instance_SBox_Instance_2_T3 ;
    wire LED_128_Instance_SBox_Instance_2_T1 ;
    wire LED_128_Instance_SBox_Instance_2_Q7 ;
    wire LED_128_Instance_SBox_Instance_2_Q6 ;
    wire LED_128_Instance_SBox_Instance_2_L5 ;
    wire LED_128_Instance_SBox_Instance_2_T2 ;
    wire LED_128_Instance_SBox_Instance_2_L4 ;
    wire LED_128_Instance_SBox_Instance_2_Q3 ;
    wire LED_128_Instance_SBox_Instance_2_L3 ;
    wire LED_128_Instance_SBox_Instance_2_Q2 ;
    wire LED_128_Instance_SBox_Instance_2_T0 ;
    wire LED_128_Instance_SBox_Instance_2_L2 ;
    wire LED_128_Instance_SBox_Instance_2_L1 ;
    wire LED_128_Instance_SBox_Instance_2_L0 ;
    wire LED_128_Instance_SBox_Instance_3_n3 ;
    wire LED_128_Instance_SBox_Instance_3_n2 ;
    wire LED_128_Instance_SBox_Instance_3_n1 ;
    wire LED_128_Instance_SBox_Instance_3_L8 ;
    wire LED_128_Instance_SBox_Instance_3_L7 ;
    wire LED_128_Instance_SBox_Instance_3_T3 ;
    wire LED_128_Instance_SBox_Instance_3_T1 ;
    wire LED_128_Instance_SBox_Instance_3_Q7 ;
    wire LED_128_Instance_SBox_Instance_3_Q6 ;
    wire LED_128_Instance_SBox_Instance_3_L5 ;
    wire LED_128_Instance_SBox_Instance_3_T2 ;
    wire LED_128_Instance_SBox_Instance_3_L4 ;
    wire LED_128_Instance_SBox_Instance_3_Q3 ;
    wire LED_128_Instance_SBox_Instance_3_L3 ;
    wire LED_128_Instance_SBox_Instance_3_Q2 ;
    wire LED_128_Instance_SBox_Instance_3_T0 ;
    wire LED_128_Instance_SBox_Instance_3_L2 ;
    wire LED_128_Instance_SBox_Instance_3_L1 ;
    wire LED_128_Instance_SBox_Instance_3_L0 ;
    wire LED_128_Instance_SBox_Instance_4_n3 ;
    wire LED_128_Instance_SBox_Instance_4_n2 ;
    wire LED_128_Instance_SBox_Instance_4_n1 ;
    wire LED_128_Instance_SBox_Instance_4_L8 ;
    wire LED_128_Instance_SBox_Instance_4_L7 ;
    wire LED_128_Instance_SBox_Instance_4_T3 ;
    wire LED_128_Instance_SBox_Instance_4_T1 ;
    wire LED_128_Instance_SBox_Instance_4_Q7 ;
    wire LED_128_Instance_SBox_Instance_4_Q6 ;
    wire LED_128_Instance_SBox_Instance_4_L5 ;
    wire LED_128_Instance_SBox_Instance_4_T2 ;
    wire LED_128_Instance_SBox_Instance_4_L4 ;
    wire LED_128_Instance_SBox_Instance_4_Q3 ;
    wire LED_128_Instance_SBox_Instance_4_L3 ;
    wire LED_128_Instance_SBox_Instance_4_Q2 ;
    wire LED_128_Instance_SBox_Instance_4_T0 ;
    wire LED_128_Instance_SBox_Instance_4_L2 ;
    wire LED_128_Instance_SBox_Instance_4_L1 ;
    wire LED_128_Instance_SBox_Instance_4_L0 ;
    wire LED_128_Instance_SBox_Instance_5_n3 ;
    wire LED_128_Instance_SBox_Instance_5_n2 ;
    wire LED_128_Instance_SBox_Instance_5_n1 ;
    wire LED_128_Instance_SBox_Instance_5_L8 ;
    wire LED_128_Instance_SBox_Instance_5_L7 ;
    wire LED_128_Instance_SBox_Instance_5_T3 ;
    wire LED_128_Instance_SBox_Instance_5_T1 ;
    wire LED_128_Instance_SBox_Instance_5_Q7 ;
    wire LED_128_Instance_SBox_Instance_5_Q6 ;
    wire LED_128_Instance_SBox_Instance_5_L5 ;
    wire LED_128_Instance_SBox_Instance_5_T2 ;
    wire LED_128_Instance_SBox_Instance_5_L4 ;
    wire LED_128_Instance_SBox_Instance_5_Q3 ;
    wire LED_128_Instance_SBox_Instance_5_L3 ;
    wire LED_128_Instance_SBox_Instance_5_Q2 ;
    wire LED_128_Instance_SBox_Instance_5_T0 ;
    wire LED_128_Instance_SBox_Instance_5_L2 ;
    wire LED_128_Instance_SBox_Instance_5_L1 ;
    wire LED_128_Instance_SBox_Instance_5_L0 ;
    wire LED_128_Instance_SBox_Instance_6_n3 ;
    wire LED_128_Instance_SBox_Instance_6_n2 ;
    wire LED_128_Instance_SBox_Instance_6_n1 ;
    wire LED_128_Instance_SBox_Instance_6_L8 ;
    wire LED_128_Instance_SBox_Instance_6_L7 ;
    wire LED_128_Instance_SBox_Instance_6_T3 ;
    wire LED_128_Instance_SBox_Instance_6_T1 ;
    wire LED_128_Instance_SBox_Instance_6_Q7 ;
    wire LED_128_Instance_SBox_Instance_6_Q6 ;
    wire LED_128_Instance_SBox_Instance_6_L5 ;
    wire LED_128_Instance_SBox_Instance_6_T2 ;
    wire LED_128_Instance_SBox_Instance_6_L4 ;
    wire LED_128_Instance_SBox_Instance_6_Q3 ;
    wire LED_128_Instance_SBox_Instance_6_L3 ;
    wire LED_128_Instance_SBox_Instance_6_Q2 ;
    wire LED_128_Instance_SBox_Instance_6_T0 ;
    wire LED_128_Instance_SBox_Instance_6_L2 ;
    wire LED_128_Instance_SBox_Instance_6_L1 ;
    wire LED_128_Instance_SBox_Instance_6_L0 ;
    wire LED_128_Instance_SBox_Instance_7_n3 ;
    wire LED_128_Instance_SBox_Instance_7_n2 ;
    wire LED_128_Instance_SBox_Instance_7_n1 ;
    wire LED_128_Instance_SBox_Instance_7_L8 ;
    wire LED_128_Instance_SBox_Instance_7_L7 ;
    wire LED_128_Instance_SBox_Instance_7_T3 ;
    wire LED_128_Instance_SBox_Instance_7_T1 ;
    wire LED_128_Instance_SBox_Instance_7_Q7 ;
    wire LED_128_Instance_SBox_Instance_7_Q6 ;
    wire LED_128_Instance_SBox_Instance_7_L5 ;
    wire LED_128_Instance_SBox_Instance_7_T2 ;
    wire LED_128_Instance_SBox_Instance_7_L4 ;
    wire LED_128_Instance_SBox_Instance_7_Q3 ;
    wire LED_128_Instance_SBox_Instance_7_L3 ;
    wire LED_128_Instance_SBox_Instance_7_Q2 ;
    wire LED_128_Instance_SBox_Instance_7_T0 ;
    wire LED_128_Instance_SBox_Instance_7_L2 ;
    wire LED_128_Instance_SBox_Instance_7_L1 ;
    wire LED_128_Instance_SBox_Instance_7_L0 ;
    wire LED_128_Instance_SBox_Instance_8_n3 ;
    wire LED_128_Instance_SBox_Instance_8_n2 ;
    wire LED_128_Instance_SBox_Instance_8_n1 ;
    wire LED_128_Instance_SBox_Instance_8_L8 ;
    wire LED_128_Instance_SBox_Instance_8_L7 ;
    wire LED_128_Instance_SBox_Instance_8_T3 ;
    wire LED_128_Instance_SBox_Instance_8_T1 ;
    wire LED_128_Instance_SBox_Instance_8_Q7 ;
    wire LED_128_Instance_SBox_Instance_8_Q6 ;
    wire LED_128_Instance_SBox_Instance_8_L5 ;
    wire LED_128_Instance_SBox_Instance_8_T2 ;
    wire LED_128_Instance_SBox_Instance_8_L4 ;
    wire LED_128_Instance_SBox_Instance_8_Q3 ;
    wire LED_128_Instance_SBox_Instance_8_L3 ;
    wire LED_128_Instance_SBox_Instance_8_Q2 ;
    wire LED_128_Instance_SBox_Instance_8_T0 ;
    wire LED_128_Instance_SBox_Instance_8_L2 ;
    wire LED_128_Instance_SBox_Instance_8_L1 ;
    wire LED_128_Instance_SBox_Instance_8_L0 ;
    wire LED_128_Instance_SBox_Instance_9_n3 ;
    wire LED_128_Instance_SBox_Instance_9_n2 ;
    wire LED_128_Instance_SBox_Instance_9_n1 ;
    wire LED_128_Instance_SBox_Instance_9_L8 ;
    wire LED_128_Instance_SBox_Instance_9_L7 ;
    wire LED_128_Instance_SBox_Instance_9_T3 ;
    wire LED_128_Instance_SBox_Instance_9_T1 ;
    wire LED_128_Instance_SBox_Instance_9_Q7 ;
    wire LED_128_Instance_SBox_Instance_9_Q6 ;
    wire LED_128_Instance_SBox_Instance_9_L5 ;
    wire LED_128_Instance_SBox_Instance_9_T2 ;
    wire LED_128_Instance_SBox_Instance_9_L4 ;
    wire LED_128_Instance_SBox_Instance_9_Q3 ;
    wire LED_128_Instance_SBox_Instance_9_L3 ;
    wire LED_128_Instance_SBox_Instance_9_Q2 ;
    wire LED_128_Instance_SBox_Instance_9_T0 ;
    wire LED_128_Instance_SBox_Instance_9_L2 ;
    wire LED_128_Instance_SBox_Instance_9_L1 ;
    wire LED_128_Instance_SBox_Instance_9_L0 ;
    wire LED_128_Instance_SBox_Instance_10_n3 ;
    wire LED_128_Instance_SBox_Instance_10_n2 ;
    wire LED_128_Instance_SBox_Instance_10_n1 ;
    wire LED_128_Instance_SBox_Instance_10_L8 ;
    wire LED_128_Instance_SBox_Instance_10_L7 ;
    wire LED_128_Instance_SBox_Instance_10_T3 ;
    wire LED_128_Instance_SBox_Instance_10_T1 ;
    wire LED_128_Instance_SBox_Instance_10_Q7 ;
    wire LED_128_Instance_SBox_Instance_10_Q6 ;
    wire LED_128_Instance_SBox_Instance_10_L5 ;
    wire LED_128_Instance_SBox_Instance_10_T2 ;
    wire LED_128_Instance_SBox_Instance_10_L4 ;
    wire LED_128_Instance_SBox_Instance_10_Q3 ;
    wire LED_128_Instance_SBox_Instance_10_L3 ;
    wire LED_128_Instance_SBox_Instance_10_Q2 ;
    wire LED_128_Instance_SBox_Instance_10_T0 ;
    wire LED_128_Instance_SBox_Instance_10_L2 ;
    wire LED_128_Instance_SBox_Instance_10_L1 ;
    wire LED_128_Instance_SBox_Instance_10_L0 ;
    wire LED_128_Instance_SBox_Instance_11_n3 ;
    wire LED_128_Instance_SBox_Instance_11_n2 ;
    wire LED_128_Instance_SBox_Instance_11_n1 ;
    wire LED_128_Instance_SBox_Instance_11_L8 ;
    wire LED_128_Instance_SBox_Instance_11_L7 ;
    wire LED_128_Instance_SBox_Instance_11_T3 ;
    wire LED_128_Instance_SBox_Instance_11_T1 ;
    wire LED_128_Instance_SBox_Instance_11_Q7 ;
    wire LED_128_Instance_SBox_Instance_11_Q6 ;
    wire LED_128_Instance_SBox_Instance_11_L5 ;
    wire LED_128_Instance_SBox_Instance_11_T2 ;
    wire LED_128_Instance_SBox_Instance_11_L4 ;
    wire LED_128_Instance_SBox_Instance_11_Q3 ;
    wire LED_128_Instance_SBox_Instance_11_L3 ;
    wire LED_128_Instance_SBox_Instance_11_Q2 ;
    wire LED_128_Instance_SBox_Instance_11_T0 ;
    wire LED_128_Instance_SBox_Instance_11_L2 ;
    wire LED_128_Instance_SBox_Instance_11_L1 ;
    wire LED_128_Instance_SBox_Instance_11_L0 ;
    wire LED_128_Instance_SBox_Instance_12_n3 ;
    wire LED_128_Instance_SBox_Instance_12_n2 ;
    wire LED_128_Instance_SBox_Instance_12_n1 ;
    wire LED_128_Instance_SBox_Instance_12_L8 ;
    wire LED_128_Instance_SBox_Instance_12_L7 ;
    wire LED_128_Instance_SBox_Instance_12_T3 ;
    wire LED_128_Instance_SBox_Instance_12_T1 ;
    wire LED_128_Instance_SBox_Instance_12_Q7 ;
    wire LED_128_Instance_SBox_Instance_12_Q6 ;
    wire LED_128_Instance_SBox_Instance_12_L5 ;
    wire LED_128_Instance_SBox_Instance_12_T2 ;
    wire LED_128_Instance_SBox_Instance_12_L4 ;
    wire LED_128_Instance_SBox_Instance_12_Q3 ;
    wire LED_128_Instance_SBox_Instance_12_L3 ;
    wire LED_128_Instance_SBox_Instance_12_Q2 ;
    wire LED_128_Instance_SBox_Instance_12_T0 ;
    wire LED_128_Instance_SBox_Instance_12_L2 ;
    wire LED_128_Instance_SBox_Instance_12_L1 ;
    wire LED_128_Instance_SBox_Instance_12_L0 ;
    wire LED_128_Instance_SBox_Instance_13_n3 ;
    wire LED_128_Instance_SBox_Instance_13_n2 ;
    wire LED_128_Instance_SBox_Instance_13_n1 ;
    wire LED_128_Instance_SBox_Instance_13_L8 ;
    wire LED_128_Instance_SBox_Instance_13_L7 ;
    wire LED_128_Instance_SBox_Instance_13_T3 ;
    wire LED_128_Instance_SBox_Instance_13_T1 ;
    wire LED_128_Instance_SBox_Instance_13_Q7 ;
    wire LED_128_Instance_SBox_Instance_13_Q6 ;
    wire LED_128_Instance_SBox_Instance_13_L5 ;
    wire LED_128_Instance_SBox_Instance_13_T2 ;
    wire LED_128_Instance_SBox_Instance_13_L4 ;
    wire LED_128_Instance_SBox_Instance_13_Q3 ;
    wire LED_128_Instance_SBox_Instance_13_L3 ;
    wire LED_128_Instance_SBox_Instance_13_Q2 ;
    wire LED_128_Instance_SBox_Instance_13_T0 ;
    wire LED_128_Instance_SBox_Instance_13_L2 ;
    wire LED_128_Instance_SBox_Instance_13_L1 ;
    wire LED_128_Instance_SBox_Instance_13_L0 ;
    wire LED_128_Instance_SBox_Instance_14_n3 ;
    wire LED_128_Instance_SBox_Instance_14_n2 ;
    wire LED_128_Instance_SBox_Instance_14_n1 ;
    wire LED_128_Instance_SBox_Instance_14_L8 ;
    wire LED_128_Instance_SBox_Instance_14_L7 ;
    wire LED_128_Instance_SBox_Instance_14_T3 ;
    wire LED_128_Instance_SBox_Instance_14_T1 ;
    wire LED_128_Instance_SBox_Instance_14_Q7 ;
    wire LED_128_Instance_SBox_Instance_14_Q6 ;
    wire LED_128_Instance_SBox_Instance_14_L5 ;
    wire LED_128_Instance_SBox_Instance_14_T2 ;
    wire LED_128_Instance_SBox_Instance_14_L4 ;
    wire LED_128_Instance_SBox_Instance_14_Q3 ;
    wire LED_128_Instance_SBox_Instance_14_L3 ;
    wire LED_128_Instance_SBox_Instance_14_Q2 ;
    wire LED_128_Instance_SBox_Instance_14_T0 ;
    wire LED_128_Instance_SBox_Instance_14_L2 ;
    wire LED_128_Instance_SBox_Instance_14_L1 ;
    wire LED_128_Instance_SBox_Instance_14_L0 ;
    wire LED_128_Instance_SBox_Instance_15_n3 ;
    wire LED_128_Instance_SBox_Instance_15_n2 ;
    wire LED_128_Instance_SBox_Instance_15_n1 ;
    wire LED_128_Instance_SBox_Instance_15_L8 ;
    wire LED_128_Instance_SBox_Instance_15_L7 ;
    wire LED_128_Instance_SBox_Instance_15_T3 ;
    wire LED_128_Instance_SBox_Instance_15_T1 ;
    wire LED_128_Instance_SBox_Instance_15_Q7 ;
    wire LED_128_Instance_SBox_Instance_15_Q6 ;
    wire LED_128_Instance_SBox_Instance_15_L5 ;
    wire LED_128_Instance_SBox_Instance_15_T2 ;
    wire LED_128_Instance_SBox_Instance_15_L4 ;
    wire LED_128_Instance_SBox_Instance_15_Q3 ;
    wire LED_128_Instance_SBox_Instance_15_L3 ;
    wire LED_128_Instance_SBox_Instance_15_Q2 ;
    wire LED_128_Instance_SBox_Instance_15_T0 ;
    wire LED_128_Instance_SBox_Instance_15_L2 ;
    wire LED_128_Instance_SBox_Instance_15_L1 ;
    wire LED_128_Instance_SBox_Instance_15_L0 ;
    wire LED_128_Instance_MCS_Instance_0_n38 ;
    wire LED_128_Instance_MCS_Instance_0_n37 ;
    wire LED_128_Instance_MCS_Instance_0_n36 ;
    wire LED_128_Instance_MCS_Instance_0_n35 ;
    wire LED_128_Instance_MCS_Instance_0_n34 ;
    wire LED_128_Instance_MCS_Instance_0_n33 ;
    wire LED_128_Instance_MCS_Instance_0_n32 ;
    wire LED_128_Instance_MCS_Instance_0_n31 ;
    wire LED_128_Instance_MCS_Instance_0_n30 ;
    wire LED_128_Instance_MCS_Instance_0_n29 ;
    wire LED_128_Instance_MCS_Instance_0_n28 ;
    wire LED_128_Instance_MCS_Instance_0_n27 ;
    wire LED_128_Instance_MCS_Instance_0_n26 ;
    wire LED_128_Instance_MCS_Instance_0_n25 ;
    wire LED_128_Instance_MCS_Instance_0_n24 ;
    wire LED_128_Instance_MCS_Instance_0_n23 ;
    wire LED_128_Instance_MCS_Instance_0_n22 ;
    wire LED_128_Instance_MCS_Instance_0_n21 ;
    wire LED_128_Instance_MCS_Instance_0_n20 ;
    wire LED_128_Instance_MCS_Instance_0_n19 ;
    wire LED_128_Instance_MCS_Instance_0_n18 ;
    wire LED_128_Instance_MCS_Instance_0_n17 ;
    wire LED_128_Instance_MCS_Instance_0_n16 ;
    wire LED_128_Instance_MCS_Instance_0_n15 ;
    wire LED_128_Instance_MCS_Instance_0_n14 ;
    wire LED_128_Instance_MCS_Instance_0_n13 ;
    wire LED_128_Instance_MCS_Instance_0_n12 ;
    wire LED_128_Instance_MCS_Instance_0_n11 ;
    wire LED_128_Instance_MCS_Instance_0_n10 ;
    wire LED_128_Instance_MCS_Instance_0_n9 ;
    wire LED_128_Instance_MCS_Instance_0_n8 ;
    wire LED_128_Instance_MCS_Instance_0_n7 ;
    wire LED_128_Instance_MCS_Instance_0_n6 ;
    wire LED_128_Instance_MCS_Instance_0_n5 ;
    wire LED_128_Instance_MCS_Instance_0_n4 ;
    wire LED_128_Instance_MCS_Instance_0_n3 ;
    wire LED_128_Instance_MCS_Instance_0_n2 ;
    wire LED_128_Instance_MCS_Instance_0_n1 ;
    wire LED_128_Instance_MCS_Instance_1_n38 ;
    wire LED_128_Instance_MCS_Instance_1_n37 ;
    wire LED_128_Instance_MCS_Instance_1_n36 ;
    wire LED_128_Instance_MCS_Instance_1_n35 ;
    wire LED_128_Instance_MCS_Instance_1_n34 ;
    wire LED_128_Instance_MCS_Instance_1_n33 ;
    wire LED_128_Instance_MCS_Instance_1_n32 ;
    wire LED_128_Instance_MCS_Instance_1_n31 ;
    wire LED_128_Instance_MCS_Instance_1_n30 ;
    wire LED_128_Instance_MCS_Instance_1_n29 ;
    wire LED_128_Instance_MCS_Instance_1_n28 ;
    wire LED_128_Instance_MCS_Instance_1_n27 ;
    wire LED_128_Instance_MCS_Instance_1_n26 ;
    wire LED_128_Instance_MCS_Instance_1_n25 ;
    wire LED_128_Instance_MCS_Instance_1_n24 ;
    wire LED_128_Instance_MCS_Instance_1_n23 ;
    wire LED_128_Instance_MCS_Instance_1_n22 ;
    wire LED_128_Instance_MCS_Instance_1_n21 ;
    wire LED_128_Instance_MCS_Instance_1_n20 ;
    wire LED_128_Instance_MCS_Instance_1_n19 ;
    wire LED_128_Instance_MCS_Instance_1_n18 ;
    wire LED_128_Instance_MCS_Instance_1_n17 ;
    wire LED_128_Instance_MCS_Instance_1_n16 ;
    wire LED_128_Instance_MCS_Instance_1_n15 ;
    wire LED_128_Instance_MCS_Instance_1_n14 ;
    wire LED_128_Instance_MCS_Instance_1_n13 ;
    wire LED_128_Instance_MCS_Instance_1_n12 ;
    wire LED_128_Instance_MCS_Instance_1_n11 ;
    wire LED_128_Instance_MCS_Instance_1_n10 ;
    wire LED_128_Instance_MCS_Instance_1_n9 ;
    wire LED_128_Instance_MCS_Instance_1_n8 ;
    wire LED_128_Instance_MCS_Instance_1_n7 ;
    wire LED_128_Instance_MCS_Instance_1_n6 ;
    wire LED_128_Instance_MCS_Instance_1_n5 ;
    wire LED_128_Instance_MCS_Instance_1_n4 ;
    wire LED_128_Instance_MCS_Instance_1_n3 ;
    wire LED_128_Instance_MCS_Instance_1_n2 ;
    wire LED_128_Instance_MCS_Instance_1_n1 ;
    wire LED_128_Instance_MCS_Instance_2_n38 ;
    wire LED_128_Instance_MCS_Instance_2_n37 ;
    wire LED_128_Instance_MCS_Instance_2_n36 ;
    wire LED_128_Instance_MCS_Instance_2_n35 ;
    wire LED_128_Instance_MCS_Instance_2_n34 ;
    wire LED_128_Instance_MCS_Instance_2_n33 ;
    wire LED_128_Instance_MCS_Instance_2_n32 ;
    wire LED_128_Instance_MCS_Instance_2_n31 ;
    wire LED_128_Instance_MCS_Instance_2_n30 ;
    wire LED_128_Instance_MCS_Instance_2_n29 ;
    wire LED_128_Instance_MCS_Instance_2_n28 ;
    wire LED_128_Instance_MCS_Instance_2_n27 ;
    wire LED_128_Instance_MCS_Instance_2_n26 ;
    wire LED_128_Instance_MCS_Instance_2_n25 ;
    wire LED_128_Instance_MCS_Instance_2_n24 ;
    wire LED_128_Instance_MCS_Instance_2_n23 ;
    wire LED_128_Instance_MCS_Instance_2_n22 ;
    wire LED_128_Instance_MCS_Instance_2_n21 ;
    wire LED_128_Instance_MCS_Instance_2_n20 ;
    wire LED_128_Instance_MCS_Instance_2_n19 ;
    wire LED_128_Instance_MCS_Instance_2_n18 ;
    wire LED_128_Instance_MCS_Instance_2_n17 ;
    wire LED_128_Instance_MCS_Instance_2_n16 ;
    wire LED_128_Instance_MCS_Instance_2_n15 ;
    wire LED_128_Instance_MCS_Instance_2_n14 ;
    wire LED_128_Instance_MCS_Instance_2_n13 ;
    wire LED_128_Instance_MCS_Instance_2_n12 ;
    wire LED_128_Instance_MCS_Instance_2_n11 ;
    wire LED_128_Instance_MCS_Instance_2_n10 ;
    wire LED_128_Instance_MCS_Instance_2_n9 ;
    wire LED_128_Instance_MCS_Instance_2_n8 ;
    wire LED_128_Instance_MCS_Instance_2_n7 ;
    wire LED_128_Instance_MCS_Instance_2_n6 ;
    wire LED_128_Instance_MCS_Instance_2_n5 ;
    wire LED_128_Instance_MCS_Instance_2_n4 ;
    wire LED_128_Instance_MCS_Instance_2_n3 ;
    wire LED_128_Instance_MCS_Instance_2_n2 ;
    wire LED_128_Instance_MCS_Instance_2_n1 ;
    wire LED_128_Instance_MCS_Instance_3_n38 ;
    wire LED_128_Instance_MCS_Instance_3_n37 ;
    wire LED_128_Instance_MCS_Instance_3_n36 ;
    wire LED_128_Instance_MCS_Instance_3_n35 ;
    wire LED_128_Instance_MCS_Instance_3_n34 ;
    wire LED_128_Instance_MCS_Instance_3_n33 ;
    wire LED_128_Instance_MCS_Instance_3_n32 ;
    wire LED_128_Instance_MCS_Instance_3_n31 ;
    wire LED_128_Instance_MCS_Instance_3_n30 ;
    wire LED_128_Instance_MCS_Instance_3_n29 ;
    wire LED_128_Instance_MCS_Instance_3_n28 ;
    wire LED_128_Instance_MCS_Instance_3_n27 ;
    wire LED_128_Instance_MCS_Instance_3_n26 ;
    wire LED_128_Instance_MCS_Instance_3_n25 ;
    wire LED_128_Instance_MCS_Instance_3_n24 ;
    wire LED_128_Instance_MCS_Instance_3_n23 ;
    wire LED_128_Instance_MCS_Instance_3_n22 ;
    wire LED_128_Instance_MCS_Instance_3_n21 ;
    wire LED_128_Instance_MCS_Instance_3_n20 ;
    wire LED_128_Instance_MCS_Instance_3_n19 ;
    wire LED_128_Instance_MCS_Instance_3_n18 ;
    wire LED_128_Instance_MCS_Instance_3_n17 ;
    wire LED_128_Instance_MCS_Instance_3_n16 ;
    wire LED_128_Instance_MCS_Instance_3_n15 ;
    wire LED_128_Instance_MCS_Instance_3_n14 ;
    wire LED_128_Instance_MCS_Instance_3_n13 ;
    wire LED_128_Instance_MCS_Instance_3_n12 ;
    wire LED_128_Instance_MCS_Instance_3_n11 ;
    wire LED_128_Instance_MCS_Instance_3_n10 ;
    wire LED_128_Instance_MCS_Instance_3_n9 ;
    wire LED_128_Instance_MCS_Instance_3_n8 ;
    wire LED_128_Instance_MCS_Instance_3_n7 ;
    wire LED_128_Instance_MCS_Instance_3_n6 ;
    wire LED_128_Instance_MCS_Instance_3_n5 ;
    wire LED_128_Instance_MCS_Instance_3_n4 ;
    wire LED_128_Instance_MCS_Instance_3_n3 ;
    wire LED_128_Instance_MCS_Instance_3_n2 ;
    wire LED_128_Instance_MCS_Instance_3_n1 ;
    wire LED_128_Instance_ks_reg_0__Q ;
    wire [5:0] roundconstant ;
    wire [63:0] LED_128_Instance_subcells_out ;
    wire [63:0] LED_128_Instance_addconst_out ;
    wire [63:0] LED_128_Instance_addroundkey_tmp ;
    wire [63:0] LED_128_Instance_current_roundkey ;
    wire [63:0] LED_128_Instance_state1 ;
    wire [63:0] LED_128_Instance_state0 ;
    wire [63:0] LED_128_Instance_mixcolumns_out ;
    wire LMDPL_pre1 ;
    wire LMDPL_pre2 ;
    wire mid_rst ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;

    /* cells in depth 0 */
    NOR2_X1 U16 ( .A1 (roundconstant[4]), .A2 (roundconstant[1]), .ZN (n14) ) ;
    NAND2_X1 U17 ( .A1 (roundconstant[0]), .A2 (n14), .ZN (n16) ) ;
    NOR2_X1 U18 ( .A1 (roundconstant[5]), .A2 (n16), .ZN (n17) ) ;
    NAND2_X1 U19 ( .A1 (roundconstant[3]), .A2 (n17), .ZN (n18) ) ;
    NOR2_X1 U20 ( .A1 (roundconstant[2]), .A2 (n18), .ZN (n19) ) ;
    NOR2_X1 U21 ( .A1 (OUT_done), .A2 (n19), .ZN (n20) ) ;
    NOR2_X1 U22 ( .A1 (IN_reset), .A2 (n20), .ZN (n15) ) ;
    NAND2_X1 LED_128_Instance_U30 ( .A1 (LED_128_Instance_n33), .A2 (LED_128_Instance_n32), .ZN (LED_128_Instance_n34) ) ;
    XNOR2_X1 LED_128_Instance_U29 ( .A (LED_128_Instance_n25), .B (LED_128_Instance_n23), .ZN (LED_128_Instance_n32) ) ;
    XOR2_X1 LED_128_Instance_U28 ( .A (LED_128_Instance_n4), .B (LED_128_Instance_n26), .Z (LED_128_Instance_n23) ) ;
    NAND2_X1 LED_128_Instance_U27 ( .A1 (LED_128_Instance_n21), .A2 (LED_128_Instance_n20), .ZN (LED_128_Instance_n33) ) ;
    NAND2_X1 LED_128_Instance_U26 ( .A1 (LED_128_Instance_n19), .A2 (LED_128_Instance_n18), .ZN (LED_128_Instance_n20) ) ;
    NOR2_X1 LED_128_Instance_U25 ( .A1 (LED_128_Instance_n24), .A2 (LED_128_Instance_n1), .ZN (LED_128_Instance_n18) ) ;
    NOR2_X1 LED_128_Instance_U24 ( .A1 (LED_128_Instance_n8), .A2 (LED_128_Instance_n4), .ZN (LED_128_Instance_n19) ) ;
    NAND2_X1 LED_128_Instance_U23 ( .A1 (LED_128_Instance_n1), .A2 (LED_128_Instance_n17), .ZN (LED_128_Instance_n21) ) ;
    AND2_X1 LED_128_Instance_U22 ( .A1 (LED_128_Instance_n8), .A2 (LED_128_Instance_n4), .ZN (LED_128_Instance_n17) ) ;
    NAND2_X1 LED_128_Instance_U21 ( .A1 (LED_128_Instance_n29), .A2 (LED_128_Instance_n14), .ZN (LED_128_Instance_n15) ) ;
    NOR2_X1 LED_128_Instance_U20 ( .A1 (LED_128_Instance_n6), .A2 (LED_128_Instance_n13), .ZN (LED_128_Instance_n14) ) ;
    NAND2_X1 LED_128_Instance_U19 ( .A1 (LED_128_Instance_n5), .A2 (roundconstant[3]), .ZN (LED_128_Instance_n13) ) ;
    NAND2_X1 LED_128_Instance_U18 ( .A1 (LED_128_Instance_n28), .A2 (LED_128_Instance_n27), .ZN (LED_128_Instance_n16) ) ;
    NOR2_X1 LED_128_Instance_U17 ( .A1 (LED_128_Instance_n28), .A2 (IN_reset), .ZN (LED_128_Instance_N9) ) ;
    NOR2_X1 LED_128_Instance_U16 ( .A1 (IN_reset), .A2 (LED_128_Instance_n30), .ZN (LED_128_Instance_N8) ) ;
    NOR2_X1 LED_128_Instance_U15 ( .A1 (IN_reset), .A2 (LED_128_Instance_n5), .ZN (LED_128_Instance_N7) ) ;
    NOR2_X1 LED_128_Instance_U14 ( .A1 (IN_reset), .A2 (LED_128_Instance_n29), .ZN (LED_128_Instance_N6) ) ;
    NOR2_X1 LED_128_Instance_U13 ( .A1 (IN_reset), .A2 (LED_128_Instance_n6), .ZN (LED_128_Instance_N5) ) ;
    NOR2_X1 LED_128_Instance_U12 ( .A1 (LED_128_Instance_n1), .A2 (IN_reset), .ZN (LED_128_Instance_N13) ) ;
    NOR2_X1 LED_128_Instance_U11 ( .A1 (LED_128_Instance_n8), .A2 (IN_reset), .ZN (LED_128_Instance_N12) ) ;
    NOR2_X1 LED_128_Instance_U10 ( .A1 (LED_128_Instance_n4), .A2 (IN_reset), .ZN (LED_128_Instance_N11) ) ;
    NOR2_X1 LED_128_Instance_U9 ( .A1 (LED_128_Instance_n2), .A2 (IN_reset), .ZN (LED_128_Instance_N10) ) ;
    OR2_X1 LED_128_Instance_U8 ( .A1 (LED_128_Instance_n2), .A2 (LED_128_Instance_n21), .ZN (LED_128_Instance_n11) ) ;
    NAND2_X1 LED_128_Instance_U7 ( .A1 (LED_128_Instance_n34), .A2 (LED_128_Instance_n11), .ZN (LED_128_Instance_n31) ) ;
    NOR2_X1 LED_128_Instance_U6 ( .A1 (LED_128_Instance_n16), .A2 (LED_128_Instance_n15), .ZN (LED_128_Instance_n22) ) ;
    INV_X1 LED_128_Instance_U5 ( .A (LED_128_Instance_n11), .ZN (LED_128_Instance_n12) ) ;
    OR2_X1 LED_128_Instance_U4 ( .A1 (IN_reset), .A2 (LED_128_Instance_n10), .ZN (LED_128_Instance_N4) ) ;
    XNOR2_X1 LED_128_Instance_U3 ( .A (LED_128_Instance_n28), .B (LED_128_Instance_n27), .ZN (LED_128_Instance_n10) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U4 ( .A (LED_128_Instance_n22), .ZN (LED_128_Instance_MUX_state0_n11) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U3 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n8) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U2 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n10) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U1 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n9) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, LED_128_Instance_mixcolumns_out[0]}), .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, LED_128_Instance_addroundkey_out_0_}), .c ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, LED_128_Instance_state0[0]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, LED_128_Instance_mixcolumns_out[1]}), .a ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, LED_128_Instance_addroundkey_out_1_}), .c ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, LED_128_Instance_state0[1]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[2]}), .a ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, LED_128_Instance_addroundkey_out_2_}), .c ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, LED_128_Instance_state0[2]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, LED_128_Instance_mixcolumns_out[3]}), .a ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, LED_128_Instance_addroundkey_out_3_}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, LED_128_Instance_state0[3]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, LED_128_Instance_mixcolumns_out[4]}), .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, LED_128_Instance_addroundkey_out_4_}), .c ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, LED_128_Instance_state0[4]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, LED_128_Instance_mixcolumns_out[5]}), .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, LED_128_Instance_addroundkey_out_5_}), .c ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, LED_128_Instance_state0[5]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, LED_128_Instance_mixcolumns_out[6]}), .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, LED_128_Instance_addroundkey_out_6_}), .c ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, LED_128_Instance_state0[6]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, LED_128_Instance_mixcolumns_out[7]}), .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, LED_128_Instance_addconst_out[7]}), .c ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, LED_128_Instance_state0[7]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_8_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, LED_128_Instance_mixcolumns_out[8]}), .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, LED_128_Instance_addconst_out[8]}), .c ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, LED_128_Instance_state0[8]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_9_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, LED_128_Instance_mixcolumns_out[9]}), .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, LED_128_Instance_addconst_out[9]}), .c ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, LED_128_Instance_state0[9]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_10_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, LED_128_Instance_mixcolumns_out[10]}), .a ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, LED_128_Instance_addconst_out[10]}), .c ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, LED_128_Instance_state0[10]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_11_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, LED_128_Instance_mixcolumns_out[11]}), .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[11]}), .c ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, LED_128_Instance_state0[11]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_12_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, LED_128_Instance_mixcolumns_out[12]}), .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, LED_128_Instance_addconst_out[12]}), .c ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, LED_128_Instance_state0[12]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_13_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, LED_128_Instance_mixcolumns_out[13]}), .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[13]}), .c ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, LED_128_Instance_state0[13]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_14_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, LED_128_Instance_mixcolumns_out[14]}), .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, LED_128_Instance_addconst_out[14]}), .c ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, LED_128_Instance_state0[14]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_15_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, LED_128_Instance_mixcolumns_out[15]}), .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, LED_128_Instance_addconst_out[15]}), .c ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, LED_128_Instance_state0[15]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_16_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, LED_128_Instance_mixcolumns_out[16]}), .a ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, LED_128_Instance_addroundkey_out_16_}), .c ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, LED_128_Instance_state0[16]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_17_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, LED_128_Instance_mixcolumns_out[17]}), .a ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, LED_128_Instance_addroundkey_out_17_}), .c ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, LED_128_Instance_state0[17]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_18_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, LED_128_Instance_mixcolumns_out[18]}), .a ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, LED_128_Instance_addroundkey_out_18_}), .c ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, LED_128_Instance_state0[18]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_19_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, LED_128_Instance_mixcolumns_out[19]}), .a ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, LED_128_Instance_addroundkey_out_19_}), .c ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, LED_128_Instance_state0[19]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_20_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, LED_128_Instance_mixcolumns_out[20]}), .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, LED_128_Instance_addroundkey_out_20_}), .c ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, LED_128_Instance_state0[20]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_21_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, LED_128_Instance_mixcolumns_out[21]}), .a ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, LED_128_Instance_addroundkey_out_21_}), .c ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, LED_128_Instance_state0[21]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_22_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, LED_128_Instance_mixcolumns_out[22]}), .a ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, LED_128_Instance_addroundkey_out_22_}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, LED_128_Instance_state0[22]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_23_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, LED_128_Instance_mixcolumns_out[23]}), .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, LED_128_Instance_addconst_out[23]}), .c ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, LED_128_Instance_state0[23]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_24_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, LED_128_Instance_mixcolumns_out[24]}), .a ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, LED_128_Instance_addconst_out[24]}), .c ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, LED_128_Instance_state0[24]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_25_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, LED_128_Instance_mixcolumns_out[25]}), .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[25]}), .c ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, LED_128_Instance_state0[25]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_26_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, LED_128_Instance_mixcolumns_out[26]}), .a ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, LED_128_Instance_addconst_out[26]}), .c ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, LED_128_Instance_state0[26]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_27_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, LED_128_Instance_mixcolumns_out[27]}), .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, LED_128_Instance_addconst_out[27]}), .c ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, LED_128_Instance_state0[27]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_28_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, LED_128_Instance_mixcolumns_out[28]}), .a ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, LED_128_Instance_addconst_out[28]}), .c ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, LED_128_Instance_state0[28]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_29_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, LED_128_Instance_mixcolumns_out[29]}), .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[29]}), .c ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, LED_128_Instance_state0[29]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_30_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, LED_128_Instance_mixcolumns_out[30]}), .a ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, LED_128_Instance_addconst_out[30]}), .c ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, LED_128_Instance_state0[30]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_31_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, LED_128_Instance_mixcolumns_out[31]}), .a ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[31]}), .c ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, LED_128_Instance_state0[31]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_32_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, LED_128_Instance_mixcolumns_out[32]}), .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, LED_128_Instance_addroundkey_out_32_}), .c ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, LED_128_Instance_state0[32]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_33_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, LED_128_Instance_mixcolumns_out[33]}), .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, LED_128_Instance_addroundkey_out_33_}), .c ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, LED_128_Instance_state0[33]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_34_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, LED_128_Instance_mixcolumns_out[34]}), .a ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, LED_128_Instance_addroundkey_out_34_}), .c ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, LED_128_Instance_state0[34]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_35_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, LED_128_Instance_mixcolumns_out[35]}), .a ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, LED_128_Instance_addroundkey_out_35_}), .c ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, LED_128_Instance_state0[35]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_36_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, LED_128_Instance_mixcolumns_out[36]}), .a ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, LED_128_Instance_addroundkey_out_36_}), .c ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, LED_128_Instance_state0[36]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_37_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, LED_128_Instance_mixcolumns_out[37]}), .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, LED_128_Instance_addroundkey_out_37_}), .c ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, LED_128_Instance_state0[37]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_38_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, LED_128_Instance_mixcolumns_out[38]}), .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, LED_128_Instance_addroundkey_out_38_}), .c ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, LED_128_Instance_state0[38]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_39_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, LED_128_Instance_mixcolumns_out[39]}), .a ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, LED_128_Instance_addconst_out[39]}), .c ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, LED_128_Instance_state0[39]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_40_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, LED_128_Instance_mixcolumns_out[40]}), .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, LED_128_Instance_addconst_out[40]}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, LED_128_Instance_state0[40]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_41_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, LED_128_Instance_mixcolumns_out[41]}), .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, LED_128_Instance_addconst_out[41]}), .c ({new_AGEMA_signal_3427, new_AGEMA_signal_3426, LED_128_Instance_state0[41]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_42_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, LED_128_Instance_mixcolumns_out[42]}), .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, LED_128_Instance_addconst_out[42]}), .c ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, LED_128_Instance_state0[42]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_43_U1 ( .s ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, LED_128_Instance_n22}), .b ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, LED_128_Instance_mixcolumns_out[43]}), .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, LED_128_Instance_addconst_out[43]}), .c ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, LED_128_Instance_state0[43]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_44_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, LED_128_Instance_mixcolumns_out[44]}), .a ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, LED_128_Instance_addconst_out[44]}), .c ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, LED_128_Instance_state0[44]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_45_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, LED_128_Instance_mixcolumns_out[45]}), .a ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, LED_128_Instance_addconst_out[45]}), .c ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, LED_128_Instance_state0[45]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_46_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, LED_128_Instance_mixcolumns_out[46]}), .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, LED_128_Instance_addconst_out[46]}), .c ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, LED_128_Instance_state0[46]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_47_U1 ( .s ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, LED_128_Instance_n22}), .b ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, LED_128_Instance_mixcolumns_out[47]}), .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, LED_128_Instance_addconst_out[47]}), .c ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, LED_128_Instance_state0[47]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_48_U1 ( .s ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, LED_128_Instance_n22}), .b ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, LED_128_Instance_mixcolumns_out[48]}), .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, LED_128_Instance_addroundkey_out_48_}), .c ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, LED_128_Instance_state0[48]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_49_U1 ( .s ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, LED_128_Instance_n22}), .b ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, LED_128_Instance_mixcolumns_out[49]}), .a ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, LED_128_Instance_addroundkey_out_49_}), .c ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, LED_128_Instance_state0[49]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_50_U1 ( .s ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, LED_128_Instance_n22}), .b ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, LED_128_Instance_mixcolumns_out[50]}), .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, LED_128_Instance_addroundkey_out_50_}), .c ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, LED_128_Instance_state0[50]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_51_U1 ( .s ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, LED_128_Instance_n22}), .b ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, LED_128_Instance_mixcolumns_out[51]}), .a ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, LED_128_Instance_addroundkey_out_51_}), .c ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, LED_128_Instance_state0[51]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_52_U1 ( .s ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, LED_128_Instance_n22}), .b ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, LED_128_Instance_mixcolumns_out[52]}), .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, LED_128_Instance_addroundkey_out_52_}), .c ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, LED_128_Instance_state0[52]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_53_U1 ( .s ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, LED_128_Instance_n22}), .b ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, LED_128_Instance_mixcolumns_out[53]}), .a ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, LED_128_Instance_addroundkey_out_53_}), .c ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, LED_128_Instance_state0[53]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_54_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, LED_128_Instance_mixcolumns_out[54]}), .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, LED_128_Instance_addroundkey_out_54_}), .c ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, LED_128_Instance_state0[54]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_55_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, LED_128_Instance_mixcolumns_out[55]}), .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, LED_128_Instance_addconst_out[55]}), .c ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, LED_128_Instance_state0[55]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_56_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, LED_128_Instance_mixcolumns_out[56]}), .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, LED_128_Instance_addconst_out[56]}), .c ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, LED_128_Instance_state0[56]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_57_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, LED_128_Instance_mixcolumns_out[57]}), .a ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, LED_128_Instance_addconst_out[57]}), .c ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, LED_128_Instance_state0[57]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_58_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, LED_128_Instance_mixcolumns_out[58]}), .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, LED_128_Instance_addconst_out[58]}), .c ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, LED_128_Instance_state0[58]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_59_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, LED_128_Instance_mixcolumns_out[59]}), .a ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, LED_128_Instance_addconst_out[59]}), .c ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, LED_128_Instance_state0[59]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_60_U1 ( .s ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, LED_128_Instance_MUX_state0_n9}), .b ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, LED_128_Instance_mixcolumns_out[60]}), .a ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, LED_128_Instance_addconst_out[60]}), .c ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, LED_128_Instance_state0[60]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_61_U1 ( .s ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, LED_128_Instance_MUX_state0_n10}), .b ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, LED_128_Instance_mixcolumns_out[61]}), .a ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, LED_128_Instance_addconst_out[61]}), .c ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, LED_128_Instance_state0[61]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_62_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, LED_128_Instance_mixcolumns_out[62]}), .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, LED_128_Instance_addconst_out[62]}), .c ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, LED_128_Instance_state0[62]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state0_mux_inst_63_U1 ( .s ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, LED_128_Instance_MUX_state0_n8}), .b ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, LED_128_Instance_mixcolumns_out[63]}), .a ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, LED_128_Instance_addconst_out[63]}), .c ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, LED_128_Instance_state0[63]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, LED_128_Instance_state0[0]}), .a ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, IN_plaintext_s0[0]}), .c ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, LED_128_Instance_state1[0]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, LED_128_Instance_state0[1]}), .a ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, IN_plaintext_s0[1]}), .c ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, LED_128_Instance_state1[1]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, LED_128_Instance_state0[2]}), .a ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, IN_plaintext_s0[2]}), .c ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, LED_128_Instance_state1[2]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, LED_128_Instance_state0[3]}), .a ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, IN_plaintext_s0[3]}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, LED_128_Instance_state1[3]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, LED_128_Instance_state0[4]}), .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, IN_plaintext_s0[4]}), .c ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, LED_128_Instance_state1[4]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, LED_128_Instance_state0[5]}), .a ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, IN_plaintext_s0[5]}), .c ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, LED_128_Instance_state1[5]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, LED_128_Instance_state0[6]}), .a ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, IN_plaintext_s0[6]}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, LED_128_Instance_state1[6]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, LED_128_Instance_state0[7]}), .a ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, IN_plaintext_s0[7]}), .c ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, LED_128_Instance_state1[7]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_8_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, LED_128_Instance_state0[8]}), .a ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, IN_plaintext_s0[8]}), .c ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, LED_128_Instance_state1[8]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_9_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, LED_128_Instance_state0[9]}), .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, IN_plaintext_s0[9]}), .c ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, LED_128_Instance_state1[9]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_10_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, LED_128_Instance_state0[10]}), .a ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, IN_plaintext_s0[10]}), .c ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, LED_128_Instance_state1[10]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_11_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, LED_128_Instance_state0[11]}), .a ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, IN_plaintext_s0[11]}), .c ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, LED_128_Instance_state1[11]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_12_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, LED_128_Instance_state0[12]}), .a ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, IN_plaintext_s0[12]}), .c ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, LED_128_Instance_state1[12]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_13_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, LED_128_Instance_state0[13]}), .a ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, IN_plaintext_s0[13]}), .c ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, LED_128_Instance_state1[13]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_14_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, LED_128_Instance_state0[14]}), .a ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, IN_plaintext_s0[14]}), .c ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, LED_128_Instance_state1[14]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_15_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, LED_128_Instance_state0[15]}), .a ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, IN_plaintext_s0[15]}), .c ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, LED_128_Instance_state1[15]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_16_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, LED_128_Instance_state0[16]}), .a ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, IN_plaintext_s0[16]}), .c ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, LED_128_Instance_state1[16]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_17_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, LED_128_Instance_state0[17]}), .a ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, IN_plaintext_s0[17]}), .c ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, LED_128_Instance_state1[17]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_18_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, LED_128_Instance_state0[18]}), .a ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, IN_plaintext_s0[18]}), .c ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, LED_128_Instance_state1[18]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_19_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, LED_128_Instance_state0[19]}), .a ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, IN_plaintext_s0[19]}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, LED_128_Instance_state1[19]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_20_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, LED_128_Instance_state0[20]}), .a ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, IN_plaintext_s0[20]}), .c ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, LED_128_Instance_state1[20]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_21_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, LED_128_Instance_state0[21]}), .a ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, IN_plaintext_s0[21]}), .c ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, LED_128_Instance_state1[21]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_22_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, LED_128_Instance_state0[22]}), .a ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, IN_plaintext_s0[22]}), .c ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, LED_128_Instance_state1[22]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_23_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, LED_128_Instance_state0[23]}), .a ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, IN_plaintext_s0[23]}), .c ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, LED_128_Instance_state1[23]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_24_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, LED_128_Instance_state0[24]}), .a ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, IN_plaintext_s0[24]}), .c ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, LED_128_Instance_state1[24]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_25_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, LED_128_Instance_state0[25]}), .a ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, IN_plaintext_s0[25]}), .c ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, LED_128_Instance_state1[25]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_26_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, LED_128_Instance_state0[26]}), .a ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, IN_plaintext_s0[26]}), .c ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, LED_128_Instance_state1[26]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_27_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, LED_128_Instance_state0[27]}), .a ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, IN_plaintext_s0[27]}), .c ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, LED_128_Instance_state1[27]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_28_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, LED_128_Instance_state0[28]}), .a ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, IN_plaintext_s0[28]}), .c ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, LED_128_Instance_state1[28]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_29_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, LED_128_Instance_state0[29]}), .a ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, IN_plaintext_s0[29]}), .c ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, LED_128_Instance_state1[29]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_30_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, LED_128_Instance_state0[30]}), .a ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, IN_plaintext_s0[30]}), .c ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, LED_128_Instance_state1[30]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_31_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, LED_128_Instance_state0[31]}), .a ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, IN_plaintext_s0[31]}), .c ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, LED_128_Instance_state1[31]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_32_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, LED_128_Instance_state0[32]}), .a ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, IN_plaintext_s0[32]}), .c ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, LED_128_Instance_state1[32]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_33_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, LED_128_Instance_state0[33]}), .a ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, IN_plaintext_s0[33]}), .c ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, LED_128_Instance_state1[33]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_34_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, LED_128_Instance_state0[34]}), .a ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, IN_plaintext_s0[34]}), .c ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, LED_128_Instance_state1[34]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_35_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, LED_128_Instance_state0[35]}), .a ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, IN_plaintext_s0[35]}), .c ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, LED_128_Instance_state1[35]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_36_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, LED_128_Instance_state0[36]}), .a ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, IN_plaintext_s0[36]}), .c ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, LED_128_Instance_state1[36]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_37_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, LED_128_Instance_state0[37]}), .a ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, IN_plaintext_s0[37]}), .c ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, LED_128_Instance_state1[37]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_38_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, LED_128_Instance_state0[38]}), .a ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, IN_plaintext_s0[38]}), .c ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, LED_128_Instance_state1[38]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_39_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, LED_128_Instance_state0[39]}), .a ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, IN_plaintext_s0[39]}), .c ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, LED_128_Instance_state1[39]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_40_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, LED_128_Instance_state0[40]}), .a ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, IN_plaintext_s0[40]}), .c ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, LED_128_Instance_state1[40]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_41_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3427, new_AGEMA_signal_3426, LED_128_Instance_state0[41]}), .a ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, IN_plaintext_s0[41]}), .c ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, LED_128_Instance_state1[41]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_42_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, LED_128_Instance_state0[42]}), .a ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, IN_plaintext_s0[42]}), .c ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, LED_128_Instance_state1[42]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_43_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, LED_128_Instance_state0[43]}), .a ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, IN_plaintext_s0[43]}), .c ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, LED_128_Instance_state1[43]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_44_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, LED_128_Instance_state0[44]}), .a ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, IN_plaintext_s0[44]}), .c ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, LED_128_Instance_state1[44]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_45_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, LED_128_Instance_state0[45]}), .a ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, IN_plaintext_s0[45]}), .c ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, LED_128_Instance_state1[45]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_46_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, LED_128_Instance_state0[46]}), .a ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, IN_plaintext_s0[46]}), .c ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, LED_128_Instance_state1[46]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_47_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, LED_128_Instance_state0[47]}), .a ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, IN_plaintext_s0[47]}), .c ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, LED_128_Instance_state1[47]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_48_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, LED_128_Instance_state0[48]}), .a ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, IN_plaintext_s0[48]}), .c ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, LED_128_Instance_state1[48]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_49_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, LED_128_Instance_state0[49]}), .a ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, IN_plaintext_s0[49]}), .c ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, LED_128_Instance_state1[49]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_50_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, LED_128_Instance_state0[50]}), .a ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, IN_plaintext_s0[50]}), .c ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, LED_128_Instance_state1[50]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_51_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, LED_128_Instance_state0[51]}), .a ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, IN_plaintext_s0[51]}), .c ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, LED_128_Instance_state1[51]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_52_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, LED_128_Instance_state0[52]}), .a ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, IN_plaintext_s0[52]}), .c ({new_AGEMA_signal_3715, new_AGEMA_signal_3714, LED_128_Instance_state1[52]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_53_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, LED_128_Instance_state0[53]}), .a ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, IN_plaintext_s0[53]}), .c ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, LED_128_Instance_state1[53]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_54_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, LED_128_Instance_state0[54]}), .a ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, IN_plaintext_s0[54]}), .c ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, LED_128_Instance_state1[54]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_55_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, LED_128_Instance_state0[55]}), .a ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, IN_plaintext_s0[55]}), .c ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, LED_128_Instance_state1[55]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_56_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, LED_128_Instance_state0[56]}), .a ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, IN_plaintext_s0[56]}), .c ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, LED_128_Instance_state1[56]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_57_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, LED_128_Instance_state0[57]}), .a ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, IN_plaintext_s0[57]}), .c ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, LED_128_Instance_state1[57]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_58_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, LED_128_Instance_state0[58]}), .a ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, IN_plaintext_s0[58]}), .c ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, LED_128_Instance_state1[58]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_59_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, LED_128_Instance_state0[59]}), .a ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, IN_plaintext_s0[59]}), .c ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, LED_128_Instance_state1[59]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_60_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, LED_128_Instance_state0[60]}), .a ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, IN_plaintext_s0[60]}), .c ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, LED_128_Instance_state1[60]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_61_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, LED_128_Instance_state0[61]}), .a ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, IN_plaintext_s0[61]}), .c ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, LED_128_Instance_state1[61]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_62_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, LED_128_Instance_state0[62]}), .a ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, IN_plaintext_s0[62]}), .c ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, LED_128_Instance_state1[62]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_state1_mux_inst_63_U1 ( .s ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, IN_reset}), .b ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, LED_128_Instance_state0[63]}), .a ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, IN_plaintext_s0[63]}), .c ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, LED_128_Instance_state1[63]}) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U4 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n9) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U3 ( .A (LED_128_Instance_n12), .ZN (LED_128_Instance_MUX_current_roundkey_n10) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U2 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n7) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U1 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n8) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, IN_key_s0[64]}), .a ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, IN_key_s0[0]}), .c ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, LED_128_Instance_current_roundkey[0]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, IN_key_s0[65]}), .a ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, IN_key_s0[1]}), .c ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, LED_128_Instance_current_roundkey[1]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, IN_key_s0[66]}), .a ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, IN_key_s0[2]}), .c ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, LED_128_Instance_current_roundkey[2]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, IN_key_s0[67]}), .a ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, IN_key_s0[3]}), .c ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, LED_128_Instance_current_roundkey[3]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, IN_key_s0[68]}), .a ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, IN_key_s0[4]}), .c ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, LED_128_Instance_current_roundkey[4]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, IN_key_s0[69]}), .a ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, IN_key_s0[5]}), .c ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, LED_128_Instance_current_roundkey[5]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, IN_key_s0[70]}), .a ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, IN_key_s0[6]}), .c ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, LED_128_Instance_current_roundkey[6]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, IN_key_s0[71]}), .a ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, IN_key_s0[7]}), .c ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, LED_128_Instance_current_roundkey[7]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, IN_key_s0[72]}), .a ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, IN_key_s0[8]}), .c ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, LED_128_Instance_current_roundkey[8]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, IN_key_s0[73]}), .a ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, IN_key_s0[9]}), .c ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, LED_128_Instance_current_roundkey[9]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, IN_key_s0[74]}), .a ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, IN_key_s0[10]}), .c ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, LED_128_Instance_current_roundkey[10]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, IN_key_s0[75]}), .a ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, IN_key_s0[11]}), .c ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, LED_128_Instance_current_roundkey[11]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, IN_key_s0[76]}), .a ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, IN_key_s0[12]}), .c ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, LED_128_Instance_current_roundkey[12]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, IN_key_s0[77]}), .a ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, IN_key_s0[13]}), .c ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, LED_128_Instance_current_roundkey[13]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, IN_key_s0[78]}), .a ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, IN_key_s0[14]}), .c ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, LED_128_Instance_current_roundkey[14]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, IN_key_s0[79]}), .a ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, IN_key_s0[15]}), .c ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, LED_128_Instance_current_roundkey[15]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, IN_key_s0[80]}), .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, IN_key_s0[16]}), .c ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, LED_128_Instance_current_roundkey[16]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, IN_key_s0[81]}), .a ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, IN_key_s0[17]}), .c ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, LED_128_Instance_current_roundkey[17]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, IN_key_s0[82]}), .a ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, IN_key_s0[18]}), .c ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, LED_128_Instance_current_roundkey[18]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, IN_key_s0[83]}), .a ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, IN_key_s0[19]}), .c ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, LED_128_Instance_current_roundkey[19]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1 ( .s ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, LED_128_Instance_MUX_current_roundkey_n9}), .b ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, IN_key_s0[84]}), .a ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, IN_key_s0[20]}), .c ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, LED_128_Instance_current_roundkey[20]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, IN_key_s0[85]}), .a ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, IN_key_s0[21]}), .c ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, LED_128_Instance_current_roundkey[21]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, IN_key_s0[86]}), .a ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, IN_key_s0[22]}), .c ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, LED_128_Instance_current_roundkey[22]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, IN_key_s0[87]}), .a ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, IN_key_s0[23]}), .c ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, LED_128_Instance_current_roundkey[23]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, IN_key_s0[88]}), .a ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, IN_key_s0[24]}), .c ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, LED_128_Instance_current_roundkey[24]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, IN_key_s0[89]}), .a ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, IN_key_s0[25]}), .c ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, LED_128_Instance_current_roundkey[25]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1371, new_AGEMA_signal_1370, IN_key_s0[90]}), .a ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, IN_key_s0[26]}), .c ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, LED_128_Instance_current_roundkey[26]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, IN_key_s0[91]}), .a ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, IN_key_s0[27]}), .c ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, LED_128_Instance_current_roundkey[27]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, IN_key_s0[92]}), .a ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, IN_key_s0[28]}), .c ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, LED_128_Instance_current_roundkey[28]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, IN_key_s0[93]}), .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, IN_key_s0[29]}), .c ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, LED_128_Instance_current_roundkey[29]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, IN_key_s0[94]}), .a ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, IN_key_s0[30]}), .c ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, LED_128_Instance_current_roundkey[30]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, IN_key_s0[95]}), .a ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, IN_key_s0[31]}), .c ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, LED_128_Instance_current_roundkey[31]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1383, new_AGEMA_signal_1382, IN_key_s0[96]}), .a ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, IN_key_s0[32]}), .c ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, LED_128_Instance_current_roundkey[32]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, IN_key_s0[97]}), .a ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, IN_key_s0[33]}), .c ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, LED_128_Instance_current_roundkey[33]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, IN_key_s0[98]}), .a ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, IN_key_s0[34]}), .c ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, LED_128_Instance_current_roundkey[34]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, IN_key_s0[99]}), .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, IN_key_s0[35]}), .c ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, LED_128_Instance_current_roundkey[35]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, IN_key_s0[100]}), .a ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, IN_key_s0[36]}), .c ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, LED_128_Instance_current_roundkey[36]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, IN_key_s0[101]}), .a ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, IN_key_s0[37]}), .c ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, LED_128_Instance_current_roundkey[37]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, IN_key_s0[102]}), .a ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, IN_key_s0[38]}), .c ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, LED_128_Instance_current_roundkey[38]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1 ( .s ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, LED_128_Instance_n12}), .b ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, IN_key_s0[103]}), .a ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, IN_key_s0[39]}), .c ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, LED_128_Instance_current_roundkey[39]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, IN_key_s0[104]}), .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, IN_key_s0[40]}), .c ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, LED_128_Instance_current_roundkey[40]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, IN_key_s0[105]}), .a ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, IN_key_s0[41]}), .c ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, LED_128_Instance_current_roundkey[41]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, IN_key_s0[106]}), .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, IN_key_s0[42]}), .c ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, LED_128_Instance_current_roundkey[42]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, IN_key_s0[107]}), .a ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, IN_key_s0[43]}), .c ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, LED_128_Instance_current_roundkey[43]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, IN_key_s0[108]}), .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, IN_key_s0[44]}), .c ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, LED_128_Instance_current_roundkey[44]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, IN_key_s0[109]}), .a ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, IN_key_s0[45]}), .c ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, LED_128_Instance_current_roundkey[45]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, IN_key_s0[110]}), .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, IN_key_s0[46]}), .c ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, LED_128_Instance_current_roundkey[46]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, IN_key_s0[111]}), .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, IN_key_s0[47]}), .c ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, LED_128_Instance_current_roundkey[47]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, IN_key_s0[112]}), .a ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, IN_key_s0[48]}), .c ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, LED_128_Instance_current_roundkey[48]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, IN_key_s0[113]}), .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, IN_key_s0[49]}), .c ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, LED_128_Instance_current_roundkey[49]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, IN_key_s0[114]}), .a ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, IN_key_s0[50]}), .c ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, LED_128_Instance_current_roundkey[50]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1 ( .s ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, LED_128_Instance_MUX_current_roundkey_n8}), .b ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, IN_key_s0[115]}), .a ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, IN_key_s0[51]}), .c ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, LED_128_Instance_current_roundkey[51]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, IN_key_s0[116]}), .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, IN_key_s0[52]}), .c ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, LED_128_Instance_current_roundkey[52]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, IN_key_s0[117]}), .a ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, IN_key_s0[53]}), .c ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, LED_128_Instance_current_roundkey[53]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, IN_key_s0[118]}), .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, IN_key_s0[54]}), .c ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, LED_128_Instance_current_roundkey[54]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, IN_key_s0[119]}), .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, IN_key_s0[55]}), .c ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, LED_128_Instance_current_roundkey[55]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, IN_key_s0[120]}), .a ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, IN_key_s0[56]}), .c ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, LED_128_Instance_current_roundkey[56]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, IN_key_s0[121]}), .a ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, IN_key_s0[57]}), .c ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, LED_128_Instance_current_roundkey[57]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, IN_key_s0[122]}), .a ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, IN_key_s0[58]}), .c ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, LED_128_Instance_current_roundkey[58]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, IN_key_s0[123]}), .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, IN_key_s0[59]}), .c ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, LED_128_Instance_current_roundkey[59]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, IN_key_s0[124]}), .a ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, IN_key_s0[60]}), .c ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, LED_128_Instance_current_roundkey[60]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, IN_key_s0[125]}), .a ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, IN_key_s0[61]}), .c ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, LED_128_Instance_current_roundkey[61]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, IN_key_s0[126]}), .a ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, IN_key_s0[62]}), .c ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, LED_128_Instance_current_roundkey[62]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1 ( .s ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, LED_128_Instance_MUX_current_roundkey_n7}), .b ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, IN_key_s0[127]}), .a ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, IN_key_s0[63]}), .c ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, LED_128_Instance_current_roundkey[63]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U64 ( .a ({new_AGEMA_signal_1793, OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .b ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, LED_128_Instance_current_roundkey[9]}), .c ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, LED_128_Instance_addroundkey_tmp[9]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U63 ( .a ({new_AGEMA_signal_1797, OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, LED_128_Instance_current_roundkey[8]}), .c ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, LED_128_Instance_addroundkey_tmp[8]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U62 ( .a ({new_AGEMA_signal_1801, OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, LED_128_Instance_current_roundkey[7]}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, LED_128_Instance_addroundkey_tmp[7]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U61 ( .a ({new_AGEMA_signal_1805, OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .b ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, LED_128_Instance_current_roundkey[6]}), .c ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, LED_128_Instance_addroundkey_tmp[6]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U60 ( .a ({new_AGEMA_signal_1809, OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .b ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, LED_128_Instance_current_roundkey[63]}), .c ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, LED_128_Instance_addroundkey_tmp[63]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U59 ( .a ({new_AGEMA_signal_1813, OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .b ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, LED_128_Instance_current_roundkey[62]}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, LED_128_Instance_addroundkey_tmp[62]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U58 ( .a ({new_AGEMA_signal_1817, OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .b ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, LED_128_Instance_current_roundkey[61]}), .c ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, LED_128_Instance_addroundkey_tmp[61]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U57 ( .a ({new_AGEMA_signal_1821, OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .b ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, LED_128_Instance_current_roundkey[60]}), .c ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, LED_128_Instance_addroundkey_tmp[60]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U56 ( .a ({new_AGEMA_signal_1825, OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .b ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, LED_128_Instance_current_roundkey[5]}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, LED_128_Instance_addroundkey_tmp[5]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U55 ( .a ({new_AGEMA_signal_1829, OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .b ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, LED_128_Instance_current_roundkey[59]}), .c ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, LED_128_Instance_addroundkey_tmp[59]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U54 ( .a ({new_AGEMA_signal_1833, OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .b ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, LED_128_Instance_current_roundkey[58]}), .c ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, LED_128_Instance_addroundkey_tmp[58]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U53 ( .a ({new_AGEMA_signal_1837, OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .b ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, LED_128_Instance_current_roundkey[57]}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, LED_128_Instance_addroundkey_tmp[57]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U52 ( .a ({new_AGEMA_signal_1841, OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .b ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, LED_128_Instance_current_roundkey[56]}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, LED_128_Instance_addroundkey_tmp[56]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U51 ( .a ({new_AGEMA_signal_1845, OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .b ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, LED_128_Instance_current_roundkey[55]}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, LED_128_Instance_addroundkey_tmp[55]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U50 ( .a ({new_AGEMA_signal_1849, OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .b ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, LED_128_Instance_current_roundkey[54]}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, LED_128_Instance_addroundkey_tmp[54]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U49 ( .a ({new_AGEMA_signal_1853, OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .b ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, LED_128_Instance_current_roundkey[53]}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, LED_128_Instance_addroundkey_tmp[53]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U48 ( .a ({new_AGEMA_signal_1857, OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .b ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, LED_128_Instance_current_roundkey[52]}), .c ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, LED_128_Instance_addroundkey_tmp[52]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U47 ( .a ({new_AGEMA_signal_1861, OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .b ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, LED_128_Instance_current_roundkey[51]}), .c ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, LED_128_Instance_addroundkey_tmp[51]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U46 ( .a ({new_AGEMA_signal_1865, OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .b ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, LED_128_Instance_current_roundkey[50]}), .c ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, LED_128_Instance_addroundkey_tmp[50]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U45 ( .a ({new_AGEMA_signal_1869, OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, LED_128_Instance_current_roundkey[4]}), .c ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, LED_128_Instance_addroundkey_tmp[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U44 ( .a ({new_AGEMA_signal_1873, OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .b ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, LED_128_Instance_current_roundkey[49]}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, LED_128_Instance_addroundkey_tmp[49]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U43 ( .a ({new_AGEMA_signal_1877, OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .b ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, LED_128_Instance_current_roundkey[48]}), .c ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, LED_128_Instance_addroundkey_tmp[48]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U42 ( .a ({new_AGEMA_signal_1881, OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .b ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, LED_128_Instance_current_roundkey[47]}), .c ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, LED_128_Instance_addroundkey_tmp[47]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U41 ( .a ({new_AGEMA_signal_1885, OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .b ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, LED_128_Instance_current_roundkey[46]}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, LED_128_Instance_addroundkey_tmp[46]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U40 ( .a ({new_AGEMA_signal_1889, OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .b ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, LED_128_Instance_current_roundkey[45]}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, LED_128_Instance_addroundkey_tmp[45]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U39 ( .a ({new_AGEMA_signal_1893, OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .b ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, LED_128_Instance_current_roundkey[44]}), .c ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, LED_128_Instance_addroundkey_tmp[44]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U38 ( .a ({new_AGEMA_signal_1897, OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .b ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, LED_128_Instance_current_roundkey[43]}), .c ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, LED_128_Instance_addroundkey_tmp[43]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U37 ( .a ({new_AGEMA_signal_1901, OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .b ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, LED_128_Instance_current_roundkey[42]}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, LED_128_Instance_addroundkey_tmp[42]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U36 ( .a ({new_AGEMA_signal_1905, OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .b ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, LED_128_Instance_current_roundkey[41]}), .c ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, LED_128_Instance_addroundkey_tmp[41]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U35 ( .a ({new_AGEMA_signal_1909, OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .b ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, LED_128_Instance_current_roundkey[40]}), .c ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, LED_128_Instance_addroundkey_tmp[40]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U34 ( .a ({new_AGEMA_signal_1413, OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .b ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, LED_128_Instance_current_roundkey[3]}), .c ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, LED_128_Instance_addroundkey_tmp[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U33 ( .a ({new_AGEMA_signal_1417, OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, LED_128_Instance_current_roundkey[39]}), .c ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, LED_128_Instance_addroundkey_tmp[39]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U32 ( .a ({new_AGEMA_signal_1913, OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .b ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, LED_128_Instance_current_roundkey[38]}), .c ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, LED_128_Instance_addroundkey_tmp[38]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U31 ( .a ({new_AGEMA_signal_1917, OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .b ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, LED_128_Instance_current_roundkey[37]}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, LED_128_Instance_addroundkey_tmp[37]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U30 ( .a ({new_AGEMA_signal_1421, OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .b ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, LED_128_Instance_current_roundkey[36]}), .c ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, LED_128_Instance_addroundkey_tmp[36]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U29 ( .a ({new_AGEMA_signal_1425, OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, LED_128_Instance_current_roundkey[35]}), .c ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, LED_128_Instance_addroundkey_tmp[35]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U28 ( .a ({new_AGEMA_signal_1429, OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, LED_128_Instance_current_roundkey[34]}), .c ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, LED_128_Instance_addroundkey_tmp[34]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U27 ( .a ({new_AGEMA_signal_1921, OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .b ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, LED_128_Instance_current_roundkey[33]}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, LED_128_Instance_addroundkey_tmp[33]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U26 ( .a ({new_AGEMA_signal_1433, OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .b ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, LED_128_Instance_current_roundkey[32]}), .c ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, LED_128_Instance_addroundkey_tmp[32]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U25 ( .a ({new_AGEMA_signal_1925, OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .b ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, LED_128_Instance_current_roundkey[31]}), .c ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, LED_128_Instance_addroundkey_tmp[31]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U24 ( .a ({new_AGEMA_signal_1929, OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, LED_128_Instance_current_roundkey[30]}), .c ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, LED_128_Instance_addroundkey_tmp[30]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U23 ( .a ({new_AGEMA_signal_1933, OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .b ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, LED_128_Instance_current_roundkey[2]}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, LED_128_Instance_addroundkey_tmp[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U22 ( .a ({new_AGEMA_signal_1937, OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .b ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, LED_128_Instance_current_roundkey[29]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, LED_128_Instance_addroundkey_tmp[29]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U21 ( .a ({new_AGEMA_signal_1437, OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .b ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, LED_128_Instance_current_roundkey[28]}), .c ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, LED_128_Instance_addroundkey_tmp[28]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U20 ( .a ({new_AGEMA_signal_1941, OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .b ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, LED_128_Instance_current_roundkey[27]}), .c ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, LED_128_Instance_addroundkey_tmp[27]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U19 ( .a ({new_AGEMA_signal_1441, OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, LED_128_Instance_current_roundkey[26]}), .c ({new_AGEMA_signal_1443, new_AGEMA_signal_1442, LED_128_Instance_addroundkey_tmp[26]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U18 ( .a ({new_AGEMA_signal_1945, OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .b ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, LED_128_Instance_current_roundkey[25]}), .c ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, LED_128_Instance_addroundkey_tmp[25]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U17 ( .a ({new_AGEMA_signal_1445, OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, LED_128_Instance_current_roundkey[24]}), .c ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, LED_128_Instance_addroundkey_tmp[24]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U16 ( .a ({new_AGEMA_signal_1949, OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .b ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, LED_128_Instance_current_roundkey[23]}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, LED_128_Instance_addroundkey_tmp[23]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U15 ( .a ({new_AGEMA_signal_1449, OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .b ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, LED_128_Instance_current_roundkey[22]}), .c ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, LED_128_Instance_addroundkey_tmp[22]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U14 ( .a ({new_AGEMA_signal_1953, OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .b ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, LED_128_Instance_current_roundkey[21]}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, LED_128_Instance_addroundkey_tmp[21]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U13 ( .a ({new_AGEMA_signal_1957, OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .b ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, LED_128_Instance_current_roundkey[20]}), .c ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, LED_128_Instance_addroundkey_tmp[20]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U12 ( .a ({new_AGEMA_signal_1961, OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .b ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, LED_128_Instance_current_roundkey[1]}), .c ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, LED_128_Instance_addroundkey_tmp[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U11 ( .a ({new_AGEMA_signal_1453, OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, LED_128_Instance_current_roundkey[19]}), .c ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, LED_128_Instance_addroundkey_tmp[19]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U10 ( .a ({new_AGEMA_signal_1965, OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .b ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, LED_128_Instance_current_roundkey[18]}), .c ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, LED_128_Instance_addroundkey_tmp[18]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U9 ( .a ({new_AGEMA_signal_1969, OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .b ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, LED_128_Instance_current_roundkey[17]}), .c ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, LED_128_Instance_addroundkey_tmp[17]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U8 ( .a ({new_AGEMA_signal_1457, OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, LED_128_Instance_current_roundkey[16]}), .c ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, LED_128_Instance_addroundkey_tmp[16]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U7 ( .a ({new_AGEMA_signal_1973, OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .b ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, LED_128_Instance_current_roundkey[15]}), .c ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, LED_128_Instance_addroundkey_tmp[15]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U6 ( .a ({new_AGEMA_signal_1977, OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .b ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, LED_128_Instance_current_roundkey[14]}), .c ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, LED_128_Instance_addroundkey_tmp[14]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U5 ( .a ({new_AGEMA_signal_1981, OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .b ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, LED_128_Instance_current_roundkey[13]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, LED_128_Instance_addroundkey_tmp[13]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U4 ( .a ({new_AGEMA_signal_1985, OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .b ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, LED_128_Instance_current_roundkey[12]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, LED_128_Instance_addroundkey_tmp[12]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U3 ( .a ({new_AGEMA_signal_1989, OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .b ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, LED_128_Instance_current_roundkey[11]}), .c ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, LED_128_Instance_addroundkey_tmp[11]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U2 ( .a ({new_AGEMA_signal_1993, OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .b ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, LED_128_Instance_current_roundkey[10]}), .c ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, LED_128_Instance_addroundkey_tmp[10]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_addRoundKey_instance_U1 ( .a ({new_AGEMA_signal_1461, OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .b ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, LED_128_Instance_current_roundkey[0]}), .c ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, LED_128_Instance_addroundkey_tmp[0]}) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U3 ( .A (LED_128_Instance_MUX_addroundkey_out_n9), .ZN (LED_128_Instance_MUX_addroundkey_out_n7) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U2 ( .A (LED_128_Instance_n31), .ZN (LED_128_Instance_MUX_addroundkey_out_n9) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U1 ( .A (LED_128_Instance_MUX_addroundkey_out_n9), .ZN (LED_128_Instance_MUX_addroundkey_out_n8) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1461, OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .a ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, LED_128_Instance_addroundkey_tmp[0]}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, LED_128_Instance_addroundkey_out_0_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1961, OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .a ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, LED_128_Instance_addroundkey_tmp[1]}), .c ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, LED_128_Instance_addroundkey_out_1_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1933, OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .a ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, LED_128_Instance_addroundkey_tmp[2]}), .c ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, LED_128_Instance_addroundkey_out_2_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1413, OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .a ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, LED_128_Instance_addroundkey_tmp[3]}), .c ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, LED_128_Instance_addroundkey_out_3_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1869, OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .a ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, LED_128_Instance_addroundkey_tmp[4]}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, LED_128_Instance_addroundkey_out_4_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1825, OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .a ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, LED_128_Instance_addroundkey_tmp[5]}), .c ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, LED_128_Instance_addroundkey_out_5_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1805, OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .a ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, LED_128_Instance_addroundkey_tmp[6]}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, LED_128_Instance_addroundkey_out_6_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1801, OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .a ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, LED_128_Instance_addroundkey_tmp[7]}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, LED_128_Instance_addconst_out[7]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1797, OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .a ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, LED_128_Instance_addroundkey_tmp[8]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, LED_128_Instance_addconst_out[8]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1793, OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .a ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, LED_128_Instance_addroundkey_tmp[9]}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, LED_128_Instance_addconst_out[9]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1993, OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, LED_128_Instance_addroundkey_tmp[10]}), .c ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, LED_128_Instance_addconst_out[10]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1989, OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .a ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, LED_128_Instance_addroundkey_tmp[11]}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[11]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1985, OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .a ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, LED_128_Instance_addroundkey_tmp[12]}), .c ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, LED_128_Instance_addconst_out[12]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1981, OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .a ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, LED_128_Instance_addroundkey_tmp[13]}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[13]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1977, OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, LED_128_Instance_addroundkey_tmp[14]}), .c ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, LED_128_Instance_addconst_out[14]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1973, OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .a ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, LED_128_Instance_addroundkey_tmp[15]}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, LED_128_Instance_addconst_out[15]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1457, OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .a ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, LED_128_Instance_addroundkey_tmp[16]}), .c ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, LED_128_Instance_addroundkey_out_16_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1969, OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .a ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, LED_128_Instance_addroundkey_tmp[17]}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, LED_128_Instance_addroundkey_out_17_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1965, OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .a ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, LED_128_Instance_addroundkey_tmp[18]}), .c ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, LED_128_Instance_addroundkey_out_18_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1453, OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .a ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, LED_128_Instance_addroundkey_tmp[19]}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, LED_128_Instance_addroundkey_out_19_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1 ( .s ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, LED_128_Instance_MUX_addroundkey_out_n8}), .b ({new_AGEMA_signal_1957, OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, LED_128_Instance_addroundkey_tmp[20]}), .c ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, LED_128_Instance_addroundkey_out_20_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1953, OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .a ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, LED_128_Instance_addroundkey_tmp[21]}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, LED_128_Instance_addroundkey_out_21_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1449, OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .a ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, LED_128_Instance_addroundkey_tmp[22]}), .c ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, LED_128_Instance_addroundkey_out_22_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1949, OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .a ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, LED_128_Instance_addroundkey_tmp[23]}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, LED_128_Instance_addconst_out[23]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1445, OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .a ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, LED_128_Instance_addroundkey_tmp[24]}), .c ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, LED_128_Instance_addconst_out[24]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1945, OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, LED_128_Instance_addroundkey_tmp[25]}), .c ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[25]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1441, OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .a ({new_AGEMA_signal_1443, new_AGEMA_signal_1442, LED_128_Instance_addroundkey_tmp[26]}), .c ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, LED_128_Instance_addconst_out[26]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1941, OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .a ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, LED_128_Instance_addroundkey_tmp[27]}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, LED_128_Instance_addconst_out[27]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1437, OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .a ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, LED_128_Instance_addroundkey_tmp[28]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, LED_128_Instance_addconst_out[28]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1937, OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .a ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, LED_128_Instance_addroundkey_tmp[29]}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[29]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1929, OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .a ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, LED_128_Instance_addroundkey_tmp[30]}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, LED_128_Instance_addconst_out[30]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1925, OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .a ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, LED_128_Instance_addroundkey_tmp[31]}), .c ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[31]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1433, OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .a ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, LED_128_Instance_addroundkey_tmp[32]}), .c ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, LED_128_Instance_addroundkey_out_32_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1921, OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .a ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, LED_128_Instance_addroundkey_tmp[33]}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, LED_128_Instance_addroundkey_out_33_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1429, OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .a ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, LED_128_Instance_addroundkey_tmp[34]}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, LED_128_Instance_addroundkey_out_34_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1425, OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .a ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, LED_128_Instance_addroundkey_tmp[35]}), .c ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, LED_128_Instance_addroundkey_out_35_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1421, OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .a ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, LED_128_Instance_addroundkey_tmp[36]}), .c ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, LED_128_Instance_addroundkey_out_36_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1917, OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .a ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, LED_128_Instance_addroundkey_tmp[37]}), .c ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, LED_128_Instance_addroundkey_out_37_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1913, OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .a ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, LED_128_Instance_addroundkey_tmp[38]}), .c ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, LED_128_Instance_addroundkey_out_38_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1417, OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .a ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, LED_128_Instance_addroundkey_tmp[39]}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, LED_128_Instance_addconst_out[39]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1909, OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .a ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, LED_128_Instance_addroundkey_tmp[40]}), .c ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, LED_128_Instance_addconst_out[40]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1905, OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .a ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, LED_128_Instance_addroundkey_tmp[41]}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, LED_128_Instance_addconst_out[41]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1901, OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .a ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, LED_128_Instance_addroundkey_tmp[42]}), .c ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, LED_128_Instance_addconst_out[42]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1897, OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, LED_128_Instance_addroundkey_tmp[43]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, LED_128_Instance_addconst_out[43]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1893, OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .a ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, LED_128_Instance_addroundkey_tmp[44]}), .c ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, LED_128_Instance_addconst_out[44]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1889, OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .a ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, LED_128_Instance_addroundkey_tmp[45]}), .c ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, LED_128_Instance_addconst_out[45]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1885, OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .a ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, LED_128_Instance_addroundkey_tmp[46]}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, LED_128_Instance_addconst_out[46]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1881, OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, LED_128_Instance_addroundkey_tmp[47]}), .c ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, LED_128_Instance_addconst_out[47]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1877, OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .a ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, LED_128_Instance_addroundkey_tmp[48]}), .c ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, LED_128_Instance_addroundkey_out_48_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1873, OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .a ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, LED_128_Instance_addroundkey_tmp[49]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, LED_128_Instance_addroundkey_out_49_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1 ( .s ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, LED_128_Instance_n31}), .b ({new_AGEMA_signal_1865, OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .a ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, LED_128_Instance_addroundkey_tmp[50]}), .c ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, LED_128_Instance_addroundkey_out_50_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1861, OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .a ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, LED_128_Instance_addroundkey_tmp[51]}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, LED_128_Instance_addroundkey_out_51_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1857, OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .a ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, LED_128_Instance_addroundkey_tmp[52]}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, LED_128_Instance_addroundkey_out_52_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1853, OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .a ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, LED_128_Instance_addroundkey_tmp[53]}), .c ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, LED_128_Instance_addroundkey_out_53_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1849, OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .a ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, LED_128_Instance_addroundkey_tmp[54]}), .c ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, LED_128_Instance_addroundkey_out_54_}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1845, OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .a ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, LED_128_Instance_addroundkey_tmp[55]}), .c ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, LED_128_Instance_addconst_out[55]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1841, OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .a ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, LED_128_Instance_addroundkey_tmp[56]}), .c ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, LED_128_Instance_addconst_out[56]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1837, OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, LED_128_Instance_addroundkey_tmp[57]}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, LED_128_Instance_addconst_out[57]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1833, OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .a ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, LED_128_Instance_addroundkey_tmp[58]}), .c ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, LED_128_Instance_addconst_out[58]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1829, OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .a ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, LED_128_Instance_addroundkey_tmp[59]}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, LED_128_Instance_addconst_out[59]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1821, OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .a ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, LED_128_Instance_addroundkey_tmp[60]}), .c ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, LED_128_Instance_addconst_out[60]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1817, OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .a ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, LED_128_Instance_addroundkey_tmp[61]}), .c ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, LED_128_Instance_addconst_out[61]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1813, OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, LED_128_Instance_addroundkey_tmp[62]}), .c ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, LED_128_Instance_addconst_out[62]}) ) ;
    mux2_masked_LMDPL LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1 ( .s ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, LED_128_Instance_MUX_addroundkey_out_n7}), .b ({new_AGEMA_signal_1809, OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .a ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, LED_128_Instance_addroundkey_tmp[63]}), .c ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, LED_128_Instance_addconst_out[63]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U28 ( .a ({LMDPL_pre1, 1'b0, roundconstant[5]}), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, LED_128_Instance_addroundkey_out_6_}), .c ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, LED_128_Instance_addconst_out[6]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U27 ( .a ({LMDPL_pre1, 1'b0, roundconstant[4]}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, LED_128_Instance_addroundkey_out_5_}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, LED_128_Instance_addconst_out[5]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U26 ( .a ({LMDPL_pre1, 1'b0, roundconstant[2]}), .b ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, LED_128_Instance_addroundkey_out_54_}), .c ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, LED_128_Instance_addconst_out[54]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U25 ( .a ({LMDPL_pre1, 1'b0, roundconstant[1]}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, LED_128_Instance_addroundkey_out_53_}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, LED_128_Instance_addconst_out[53]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U24 ( .a ({LMDPL_pre1, 1'b0, roundconstant[0]}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, LED_128_Instance_addroundkey_out_52_}), .c ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, LED_128_Instance_addconst_out[52]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U23 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, LED_128_Instance_addroundkey_out_51_}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, LED_128_Instance_addconst_out[51]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U22 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, LED_128_Instance_addroundkey_out_50_}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, LED_128_Instance_addconst_out[50]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U21 ( .a ({LMDPL_pre1, 1'b0, roundconstant[3]}), .b ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, LED_128_Instance_addroundkey_out_4_}), .c ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, LED_128_Instance_addconst_out[4]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_AddConstants_instance_U20 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, LED_128_Instance_addroundkey_out_49_}), .c ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, LED_128_Instance_addconst_out[49]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_AddConstants_instance_U19 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, LED_128_Instance_addroundkey_out_48_}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, LED_128_Instance_addconst_out[48]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U18 ( .a ({LMDPL_pre1, 1'b0, 1'b1}), .b ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, LED_128_Instance_addroundkey_out_3_}), .c ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, LED_128_Instance_addconst_out[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U17 ( .a ({LMDPL_pre1, 1'b0, roundconstant[5]}), .b ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, LED_128_Instance_addroundkey_out_38_}), .c ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, LED_128_Instance_addconst_out[38]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U16 ( .a ({LMDPL_pre1, 1'b0, roundconstant[4]}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, LED_128_Instance_addroundkey_out_37_}), .c ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, LED_128_Instance_addconst_out[37]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U15 ( .a ({LMDPL_pre1, 1'b0, roundconstant[3]}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, LED_128_Instance_addroundkey_out_36_}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, LED_128_Instance_addconst_out[36]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U14 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, LED_128_Instance_addroundkey_out_35_}), .c ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, LED_128_Instance_addconst_out[35]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U13 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, LED_128_Instance_addroundkey_out_34_}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, LED_128_Instance_addconst_out[34]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_AddConstants_instance_U12 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, LED_128_Instance_addroundkey_out_33_}), .c ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, LED_128_Instance_addconst_out[33]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U11 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, LED_128_Instance_addroundkey_out_32_}), .c ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, LED_128_Instance_addconst_out[32]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U10 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, LED_128_Instance_addroundkey_out_2_}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, LED_128_Instance_addconst_out[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U9 ( .a ({LMDPL_pre1, 1'b0, roundconstant[2]}), .b ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, LED_128_Instance_addroundkey_out_22_}), .c ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, LED_128_Instance_addconst_out[22]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U8 ( .a ({LMDPL_pre1, 1'b0, roundconstant[1]}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, LED_128_Instance_addroundkey_out_21_}), .c ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, LED_128_Instance_addconst_out[21]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U7 ( .a ({LMDPL_pre1, 1'b0, roundconstant[0]}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, LED_128_Instance_addroundkey_out_20_}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, LED_128_Instance_addconst_out[20]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U6 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, LED_128_Instance_addroundkey_out_1_}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, LED_128_Instance_addconst_out[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U5 ( .a ({LMDPL_pre1, 1'b0, 1'b1}), .b ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, LED_128_Instance_addroundkey_out_19_}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, LED_128_Instance_addconst_out[19]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U4 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, LED_128_Instance_addroundkey_out_18_}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, LED_128_Instance_addconst_out[18]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U3 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, LED_128_Instance_addroundkey_out_17_}), .c ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, LED_128_Instance_addconst_out[17]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_AddConstants_instance_U2 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, LED_128_Instance_addroundkey_out_16_}), .c ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, LED_128_Instance_addconst_out[16]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_AddConstants_instance_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, LED_128_Instance_addroundkey_out_0_}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, LED_128_Instance_addconst_out[0]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_0_U3 ( .x ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, LED_128_Instance_SBox_Instance_0_L0}), .y ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, LED_128_Instance_SBox_Instance_0_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_0_U2 ( .x ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, LED_128_Instance_addconst_out[3]}), .y ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, LED_128_Instance_SBox_Instance_0_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_0_U1 ( .x ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, LED_128_Instance_addconst_out[1]}), .y ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, LED_128_Instance_SBox_Instance_0_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR1_U1 ( .a ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, LED_128_Instance_addconst_out[2]}), .b ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, LED_128_Instance_addconst_out[1]}), .c ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, LED_128_Instance_SBox_Instance_0_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR2_U1 ( .a ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, LED_128_Instance_addconst_out[1]}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, LED_128_Instance_addconst_out[0]}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, LED_128_Instance_SBox_Instance_0_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR3_U1 ( .a ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, LED_128_Instance_SBox_Instance_0_L1}), .b ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, LED_128_Instance_addconst_out[3]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, LED_128_Instance_SBox_Instance_0_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_0_XOR16_U1 ( .a ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, LED_128_Instance_SBox_Instance_0_T0}), .b ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, LED_128_Instance_SBox_Instance_0_L2}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, LED_128_Instance_SBox_Instance_0_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR4_U1 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, LED_128_Instance_addconst_out[0]}), .c ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, LED_128_Instance_SBox_Instance_0_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR5_U1 ( .a ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, LED_128_Instance_SBox_Instance_0_L3}), .b ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, LED_128_Instance_SBox_Instance_0_L0}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, LED_128_Instance_SBox_Instance_0_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR6_U1 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, LED_128_Instance_addconst_out[1]}), .c ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, LED_128_Instance_SBox_Instance_0_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR7_U1 ( .a ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, LED_128_Instance_SBox_Instance_0_T0}), .b ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, LED_128_Instance_SBox_Instance_0_T2}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, LED_128_Instance_SBox_Instance_0_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_0_XOR8_U1 ( .a ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, LED_128_Instance_SBox_Instance_0_L4}), .b ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, LED_128_Instance_SBox_Instance_0_L5}), .c ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, LED_128_Instance_SBox_Instance_0_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR9_U1 ( .a ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, LED_128_Instance_SBox_Instance_0_L1}), .b ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, LED_128_Instance_addconst_out[2]}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, LED_128_Instance_SBox_Instance_0_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_0_AND1_U1 ( .a ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, LED_128_Instance_SBox_Instance_0_n1}), .b ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, LED_128_Instance_SBox_Instance_0_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[0]), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, LED_128_Instance_SBox_Instance_0_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_0_AND2_U1 ( .a ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, LED_128_Instance_SBox_Instance_0_Q2}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, LED_128_Instance_SBox_Instance_0_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[1]), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, LED_128_Instance_SBox_Instance_0_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_0_AND3_U1 ( .a ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, LED_128_Instance_SBox_Instance_0_n3}), .b ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, LED_128_Instance_addconst_out[2]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[2]), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, LED_128_Instance_SBox_Instance_0_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_0_AND4_U1 ( .a ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, LED_128_Instance_SBox_Instance_0_Q6}), .b ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, LED_128_Instance_SBox_Instance_0_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[3]), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, LED_128_Instance_SBox_Instance_0_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR10_U1 ( .a ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, LED_128_Instance_SBox_Instance_0_L5}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, LED_128_Instance_SBox_Instance_0_T3}), .c ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, LED_128_Instance_SBox_Instance_0_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR11_U1 ( .a ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, LED_128_Instance_addconst_out[0]}), .b ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, LED_128_Instance_SBox_Instance_0_L7}), .c ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, LED_128_Instance_subcells_out[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR12_U1 ( .a ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, LED_128_Instance_SBox_Instance_0_L5}), .b ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, LED_128_Instance_SBox_Instance_0_T1}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, LED_128_Instance_SBox_Instance_0_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR13_U1 ( .a ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, LED_128_Instance_SBox_Instance_0_L1}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, LED_128_Instance_SBox_Instance_0_L8}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, LED_128_Instance_subcells_out[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR14_U1 ( .a ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, LED_128_Instance_SBox_Instance_0_L4}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, LED_128_Instance_SBox_Instance_0_T3}), .c ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, LED_128_Instance_subcells_out[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR15_U1 ( .a ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, LED_128_Instance_SBox_Instance_0_L3}), .b ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, LED_128_Instance_SBox_Instance_0_T2}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, LED_128_Instance_subcells_out[0]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_1_U3 ( .x ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, LED_128_Instance_SBox_Instance_1_L0}), .y ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, LED_128_Instance_SBox_Instance_1_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_1_U2 ( .x ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, LED_128_Instance_addconst_out[7]}), .y ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, LED_128_Instance_SBox_Instance_1_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_1_U1 ( .x ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, LED_128_Instance_addconst_out[5]}), .y ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, LED_128_Instance_SBox_Instance_1_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR1_U1 ( .a ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, LED_128_Instance_addconst_out[6]}), .b ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, LED_128_Instance_addconst_out[5]}), .c ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, LED_128_Instance_SBox_Instance_1_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR2_U1 ( .a ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, LED_128_Instance_addconst_out[5]}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, LED_128_Instance_addconst_out[4]}), .c ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, LED_128_Instance_SBox_Instance_1_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR3_U1 ( .a ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, LED_128_Instance_SBox_Instance_1_L1}), .b ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, LED_128_Instance_addconst_out[7]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, LED_128_Instance_SBox_Instance_1_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_1_XOR16_U1 ( .a ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, LED_128_Instance_SBox_Instance_1_T0}), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, LED_128_Instance_SBox_Instance_1_L2}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, LED_128_Instance_SBox_Instance_1_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR4_U1 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, LED_128_Instance_addconst_out[4]}), .c ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, LED_128_Instance_SBox_Instance_1_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR5_U1 ( .a ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, LED_128_Instance_SBox_Instance_1_L3}), .b ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, LED_128_Instance_SBox_Instance_1_L0}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, LED_128_Instance_SBox_Instance_1_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR6_U1 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, LED_128_Instance_addconst_out[5]}), .c ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, LED_128_Instance_SBox_Instance_1_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR7_U1 ( .a ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, LED_128_Instance_SBox_Instance_1_T0}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, LED_128_Instance_SBox_Instance_1_T2}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, LED_128_Instance_SBox_Instance_1_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_1_XOR8_U1 ( .a ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, LED_128_Instance_SBox_Instance_1_L4}), .b ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, LED_128_Instance_SBox_Instance_1_L5}), .c ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, LED_128_Instance_SBox_Instance_1_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR9_U1 ( .a ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, LED_128_Instance_SBox_Instance_1_L1}), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, LED_128_Instance_addconst_out[6]}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, LED_128_Instance_SBox_Instance_1_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_1_AND1_U1 ( .a ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, LED_128_Instance_SBox_Instance_1_n1}), .b ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, LED_128_Instance_SBox_Instance_1_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[4]), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, LED_128_Instance_SBox_Instance_1_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_1_AND2_U1 ( .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, LED_128_Instance_SBox_Instance_1_Q2}), .b ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, LED_128_Instance_SBox_Instance_1_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[5]), .c ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, LED_128_Instance_SBox_Instance_1_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_1_AND3_U1 ( .a ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, LED_128_Instance_SBox_Instance_1_n3}), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, LED_128_Instance_addconst_out[6]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[6]), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, LED_128_Instance_SBox_Instance_1_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_1_AND4_U1 ( .a ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, LED_128_Instance_SBox_Instance_1_Q6}), .b ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, LED_128_Instance_SBox_Instance_1_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[7]), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, LED_128_Instance_SBox_Instance_1_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR10_U1 ( .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, LED_128_Instance_SBox_Instance_1_L5}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, LED_128_Instance_SBox_Instance_1_T3}), .c ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, LED_128_Instance_SBox_Instance_1_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR11_U1 ( .a ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, LED_128_Instance_addconst_out[4]}), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, LED_128_Instance_SBox_Instance_1_L7}), .c ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, LED_128_Instance_subcells_out[7]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR12_U1 ( .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, LED_128_Instance_SBox_Instance_1_L5}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, LED_128_Instance_SBox_Instance_1_T1}), .c ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, LED_128_Instance_SBox_Instance_1_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR13_U1 ( .a ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, LED_128_Instance_SBox_Instance_1_L1}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, LED_128_Instance_SBox_Instance_1_L8}), .c ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, LED_128_Instance_subcells_out[6]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR14_U1 ( .a ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, LED_128_Instance_SBox_Instance_1_L4}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, LED_128_Instance_SBox_Instance_1_T3}), .c ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, LED_128_Instance_subcells_out[5]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR15_U1 ( .a ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, LED_128_Instance_SBox_Instance_1_L3}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, LED_128_Instance_SBox_Instance_1_T2}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, LED_128_Instance_subcells_out[4]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_2_U3 ( .x ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, LED_128_Instance_SBox_Instance_2_L0}), .y ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, LED_128_Instance_SBox_Instance_2_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_2_U2 ( .x ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[11]}), .y ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, LED_128_Instance_SBox_Instance_2_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_2_U1 ( .x ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, LED_128_Instance_addconst_out[9]}), .y ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, LED_128_Instance_SBox_Instance_2_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR1_U1 ( .a ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, LED_128_Instance_addconst_out[10]}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, LED_128_Instance_addconst_out[9]}), .c ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, LED_128_Instance_SBox_Instance_2_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR2_U1 ( .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, LED_128_Instance_addconst_out[9]}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, LED_128_Instance_addconst_out[8]}), .c ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, LED_128_Instance_SBox_Instance_2_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR3_U1 ( .a ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, LED_128_Instance_SBox_Instance_2_L1}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[11]}), .c ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, LED_128_Instance_SBox_Instance_2_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_2_XOR16_U1 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, LED_128_Instance_SBox_Instance_2_T0}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, LED_128_Instance_SBox_Instance_2_L2}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, LED_128_Instance_SBox_Instance_2_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR4_U1 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, LED_128_Instance_addconst_out[8]}), .c ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, LED_128_Instance_SBox_Instance_2_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR5_U1 ( .a ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, LED_128_Instance_SBox_Instance_2_L3}), .b ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, LED_128_Instance_SBox_Instance_2_L0}), .c ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, LED_128_Instance_SBox_Instance_2_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR6_U1 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, LED_128_Instance_addconst_out[9]}), .c ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, LED_128_Instance_SBox_Instance_2_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR7_U1 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, LED_128_Instance_SBox_Instance_2_T0}), .b ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, LED_128_Instance_SBox_Instance_2_T2}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, LED_128_Instance_SBox_Instance_2_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_2_XOR8_U1 ( .a ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, LED_128_Instance_SBox_Instance_2_L4}), .b ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, LED_128_Instance_SBox_Instance_2_L5}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, LED_128_Instance_SBox_Instance_2_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR9_U1 ( .a ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, LED_128_Instance_SBox_Instance_2_L1}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, LED_128_Instance_addconst_out[10]}), .c ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, LED_128_Instance_SBox_Instance_2_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_2_AND1_U1 ( .a ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, LED_128_Instance_SBox_Instance_2_n1}), .b ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, LED_128_Instance_SBox_Instance_2_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[8]), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, LED_128_Instance_SBox_Instance_2_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_2_AND2_U1 ( .a ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, LED_128_Instance_SBox_Instance_2_Q2}), .b ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, LED_128_Instance_SBox_Instance_2_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[9]), .c ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, LED_128_Instance_SBox_Instance_2_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_2_AND3_U1 ( .a ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, LED_128_Instance_SBox_Instance_2_n3}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, LED_128_Instance_addconst_out[10]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[10]), .c ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, LED_128_Instance_SBox_Instance_2_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_2_AND4_U1 ( .a ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, LED_128_Instance_SBox_Instance_2_Q6}), .b ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, LED_128_Instance_SBox_Instance_2_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[11]), .c ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, LED_128_Instance_SBox_Instance_2_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR10_U1 ( .a ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, LED_128_Instance_SBox_Instance_2_L5}), .b ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, LED_128_Instance_SBox_Instance_2_T3}), .c ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, LED_128_Instance_SBox_Instance_2_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR11_U1 ( .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, LED_128_Instance_addconst_out[8]}), .b ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, LED_128_Instance_SBox_Instance_2_L7}), .c ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, LED_128_Instance_subcells_out[11]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR12_U1 ( .a ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, LED_128_Instance_SBox_Instance_2_L5}), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, LED_128_Instance_SBox_Instance_2_T1}), .c ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, LED_128_Instance_SBox_Instance_2_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR13_U1 ( .a ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, LED_128_Instance_SBox_Instance_2_L1}), .b ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, LED_128_Instance_SBox_Instance_2_L8}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, LED_128_Instance_subcells_out[10]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR14_U1 ( .a ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, LED_128_Instance_SBox_Instance_2_L4}), .b ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, LED_128_Instance_SBox_Instance_2_T3}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, LED_128_Instance_subcells_out[9]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR15_U1 ( .a ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, LED_128_Instance_SBox_Instance_2_L3}), .b ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, LED_128_Instance_SBox_Instance_2_T2}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, LED_128_Instance_subcells_out[8]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_3_U3 ( .x ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, LED_128_Instance_SBox_Instance_3_L0}), .y ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, LED_128_Instance_SBox_Instance_3_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_3_U2 ( .x ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, LED_128_Instance_addconst_out[15]}), .y ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, LED_128_Instance_SBox_Instance_3_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_3_U1 ( .x ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[13]}), .y ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, LED_128_Instance_SBox_Instance_3_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR1_U1 ( .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, LED_128_Instance_addconst_out[14]}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[13]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, LED_128_Instance_SBox_Instance_3_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR2_U1 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[13]}), .b ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, LED_128_Instance_addconst_out[12]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, LED_128_Instance_SBox_Instance_3_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR3_U1 ( .a ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, LED_128_Instance_SBox_Instance_3_L1}), .b ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, LED_128_Instance_addconst_out[15]}), .c ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, LED_128_Instance_SBox_Instance_3_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_3_XOR16_U1 ( .a ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, LED_128_Instance_SBox_Instance_3_T0}), .b ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, LED_128_Instance_SBox_Instance_3_L2}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, LED_128_Instance_SBox_Instance_3_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR4_U1 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, LED_128_Instance_addconst_out[12]}), .c ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, LED_128_Instance_SBox_Instance_3_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR5_U1 ( .a ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, LED_128_Instance_SBox_Instance_3_L3}), .b ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, LED_128_Instance_SBox_Instance_3_L0}), .c ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, LED_128_Instance_SBox_Instance_3_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR6_U1 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, LED_128_Instance_addconst_out[13]}), .c ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, LED_128_Instance_SBox_Instance_3_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR7_U1 ( .a ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, LED_128_Instance_SBox_Instance_3_T0}), .b ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, LED_128_Instance_SBox_Instance_3_T2}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, LED_128_Instance_SBox_Instance_3_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_3_XOR8_U1 ( .a ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, LED_128_Instance_SBox_Instance_3_L4}), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, LED_128_Instance_SBox_Instance_3_L5}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, LED_128_Instance_SBox_Instance_3_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR9_U1 ( .a ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, LED_128_Instance_SBox_Instance_3_L1}), .b ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, LED_128_Instance_addconst_out[14]}), .c ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, LED_128_Instance_SBox_Instance_3_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_3_AND1_U1 ( .a ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, LED_128_Instance_SBox_Instance_3_n1}), .b ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, LED_128_Instance_SBox_Instance_3_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[12]), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, LED_128_Instance_SBox_Instance_3_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_3_AND2_U1 ( .a ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, LED_128_Instance_SBox_Instance_3_Q2}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, LED_128_Instance_SBox_Instance_3_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[13]), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, LED_128_Instance_SBox_Instance_3_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_3_AND3_U1 ( .a ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, LED_128_Instance_SBox_Instance_3_n3}), .b ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, LED_128_Instance_addconst_out[14]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[14]), .c ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, LED_128_Instance_SBox_Instance_3_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_3_AND4_U1 ( .a ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, LED_128_Instance_SBox_Instance_3_Q6}), .b ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, LED_128_Instance_SBox_Instance_3_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[15]), .c ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, LED_128_Instance_SBox_Instance_3_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR10_U1 ( .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, LED_128_Instance_SBox_Instance_3_L5}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, LED_128_Instance_SBox_Instance_3_T3}), .c ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, LED_128_Instance_SBox_Instance_3_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR11_U1 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, LED_128_Instance_addconst_out[12]}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, LED_128_Instance_SBox_Instance_3_L7}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, LED_128_Instance_subcells_out[15]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR12_U1 ( .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, LED_128_Instance_SBox_Instance_3_L5}), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, LED_128_Instance_SBox_Instance_3_T1}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, LED_128_Instance_SBox_Instance_3_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR13_U1 ( .a ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, LED_128_Instance_SBox_Instance_3_L1}), .b ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, LED_128_Instance_SBox_Instance_3_L8}), .c ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, LED_128_Instance_subcells_out[14]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR14_U1 ( .a ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, LED_128_Instance_SBox_Instance_3_L4}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, LED_128_Instance_SBox_Instance_3_T3}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, LED_128_Instance_subcells_out[13]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR15_U1 ( .a ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, LED_128_Instance_SBox_Instance_3_L3}), .b ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, LED_128_Instance_SBox_Instance_3_T2}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, LED_128_Instance_subcells_out[12]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_4_U3 ( .x ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, LED_128_Instance_SBox_Instance_4_L0}), .y ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, LED_128_Instance_SBox_Instance_4_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_4_U2 ( .x ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, LED_128_Instance_addconst_out[19]}), .y ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, LED_128_Instance_SBox_Instance_4_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_4_U1 ( .x ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, LED_128_Instance_addconst_out[17]}), .y ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, LED_128_Instance_SBox_Instance_4_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR1_U1 ( .a ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, LED_128_Instance_addconst_out[18]}), .b ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, LED_128_Instance_addconst_out[17]}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, LED_128_Instance_SBox_Instance_4_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR2_U1 ( .a ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, LED_128_Instance_addconst_out[17]}), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, LED_128_Instance_addconst_out[16]}), .c ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, LED_128_Instance_SBox_Instance_4_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR3_U1 ( .a ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, LED_128_Instance_SBox_Instance_4_L1}), .b ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, LED_128_Instance_addconst_out[19]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, LED_128_Instance_SBox_Instance_4_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_4_XOR16_U1 ( .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, LED_128_Instance_SBox_Instance_4_T0}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, LED_128_Instance_SBox_Instance_4_L2}), .c ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, LED_128_Instance_SBox_Instance_4_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR4_U1 ( .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, LED_128_Instance_addconst_out[16]}), .c ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, LED_128_Instance_SBox_Instance_4_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR5_U1 ( .a ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, LED_128_Instance_SBox_Instance_4_L3}), .b ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, LED_128_Instance_SBox_Instance_4_L0}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, LED_128_Instance_SBox_Instance_4_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR6_U1 ( .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, LED_128_Instance_addconst_out[17]}), .c ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, LED_128_Instance_SBox_Instance_4_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR7_U1 ( .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, LED_128_Instance_SBox_Instance_4_T0}), .b ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, LED_128_Instance_SBox_Instance_4_T2}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, LED_128_Instance_SBox_Instance_4_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_4_XOR8_U1 ( .a ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, LED_128_Instance_SBox_Instance_4_L4}), .b ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, LED_128_Instance_SBox_Instance_4_L5}), .c ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, LED_128_Instance_SBox_Instance_4_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR9_U1 ( .a ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, LED_128_Instance_SBox_Instance_4_L1}), .b ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, LED_128_Instance_addconst_out[18]}), .c ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, LED_128_Instance_SBox_Instance_4_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_4_AND1_U1 ( .a ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, LED_128_Instance_SBox_Instance_4_n1}), .b ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, LED_128_Instance_SBox_Instance_4_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[16]), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, LED_128_Instance_SBox_Instance_4_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_4_AND2_U1 ( .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, LED_128_Instance_SBox_Instance_4_Q2}), .b ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, LED_128_Instance_SBox_Instance_4_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[17]), .c ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, LED_128_Instance_SBox_Instance_4_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_4_AND3_U1 ( .a ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, LED_128_Instance_SBox_Instance_4_n3}), .b ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, LED_128_Instance_addconst_out[18]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[18]), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, LED_128_Instance_SBox_Instance_4_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_4_AND4_U1 ( .a ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, LED_128_Instance_SBox_Instance_4_Q6}), .b ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, LED_128_Instance_SBox_Instance_4_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[19]), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, LED_128_Instance_SBox_Instance_4_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR10_U1 ( .a ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, LED_128_Instance_SBox_Instance_4_L5}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, LED_128_Instance_SBox_Instance_4_T3}), .c ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, LED_128_Instance_SBox_Instance_4_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR11_U1 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, LED_128_Instance_addconst_out[16]}), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, LED_128_Instance_SBox_Instance_4_L7}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, LED_128_Instance_subcells_out[19]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR12_U1 ( .a ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, LED_128_Instance_SBox_Instance_4_L5}), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, LED_128_Instance_SBox_Instance_4_T1}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, LED_128_Instance_SBox_Instance_4_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR13_U1 ( .a ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, LED_128_Instance_SBox_Instance_4_L1}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, LED_128_Instance_SBox_Instance_4_L8}), .c ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, LED_128_Instance_subcells_out[18]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR14_U1 ( .a ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, LED_128_Instance_SBox_Instance_4_L4}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, LED_128_Instance_SBox_Instance_4_T3}), .c ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, LED_128_Instance_subcells_out[17]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR15_U1 ( .a ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, LED_128_Instance_SBox_Instance_4_L3}), .b ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, LED_128_Instance_SBox_Instance_4_T2}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, LED_128_Instance_subcells_out[16]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_5_U3 ( .x ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, LED_128_Instance_SBox_Instance_5_L0}), .y ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, LED_128_Instance_SBox_Instance_5_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_5_U2 ( .x ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, LED_128_Instance_addconst_out[23]}), .y ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, LED_128_Instance_SBox_Instance_5_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_5_U1 ( .x ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, LED_128_Instance_addconst_out[21]}), .y ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, LED_128_Instance_SBox_Instance_5_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR1_U1 ( .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, LED_128_Instance_addconst_out[22]}), .b ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, LED_128_Instance_addconst_out[21]}), .c ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, LED_128_Instance_SBox_Instance_5_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR2_U1 ( .a ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, LED_128_Instance_addconst_out[21]}), .b ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, LED_128_Instance_addconst_out[20]}), .c ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, LED_128_Instance_SBox_Instance_5_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR3_U1 ( .a ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, LED_128_Instance_SBox_Instance_5_L1}), .b ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, LED_128_Instance_addconst_out[23]}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, LED_128_Instance_SBox_Instance_5_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_5_XOR16_U1 ( .a ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, LED_128_Instance_SBox_Instance_5_T0}), .b ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, LED_128_Instance_SBox_Instance_5_L2}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, LED_128_Instance_SBox_Instance_5_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR4_U1 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, LED_128_Instance_addconst_out[20]}), .c ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, LED_128_Instance_SBox_Instance_5_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR5_U1 ( .a ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, LED_128_Instance_SBox_Instance_5_L3}), .b ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, LED_128_Instance_SBox_Instance_5_L0}), .c ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, LED_128_Instance_SBox_Instance_5_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR6_U1 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, LED_128_Instance_addconst_out[21]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, LED_128_Instance_SBox_Instance_5_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR7_U1 ( .a ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, LED_128_Instance_SBox_Instance_5_T0}), .b ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, LED_128_Instance_SBox_Instance_5_T2}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, LED_128_Instance_SBox_Instance_5_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_5_XOR8_U1 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, LED_128_Instance_SBox_Instance_5_L4}), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, LED_128_Instance_SBox_Instance_5_L5}), .c ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, LED_128_Instance_SBox_Instance_5_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR9_U1 ( .a ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, LED_128_Instance_SBox_Instance_5_L1}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, LED_128_Instance_addconst_out[22]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, LED_128_Instance_SBox_Instance_5_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_5_AND1_U1 ( .a ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, LED_128_Instance_SBox_Instance_5_n1}), .b ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, LED_128_Instance_SBox_Instance_5_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[20]), .c ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, LED_128_Instance_SBox_Instance_5_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_5_AND2_U1 ( .a ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, LED_128_Instance_SBox_Instance_5_Q2}), .b ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, LED_128_Instance_SBox_Instance_5_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[21]), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, LED_128_Instance_SBox_Instance_5_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_5_AND3_U1 ( .a ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, LED_128_Instance_SBox_Instance_5_n3}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, LED_128_Instance_addconst_out[22]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[22]), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, LED_128_Instance_SBox_Instance_5_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_5_AND4_U1 ( .a ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, LED_128_Instance_SBox_Instance_5_Q6}), .b ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, LED_128_Instance_SBox_Instance_5_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[23]), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, LED_128_Instance_SBox_Instance_5_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR10_U1 ( .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, LED_128_Instance_SBox_Instance_5_L5}), .b ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, LED_128_Instance_SBox_Instance_5_T3}), .c ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, LED_128_Instance_SBox_Instance_5_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR11_U1 ( .a ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, LED_128_Instance_addconst_out[20]}), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, LED_128_Instance_SBox_Instance_5_L7}), .c ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, LED_128_Instance_subcells_out[23]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR12_U1 ( .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, LED_128_Instance_SBox_Instance_5_L5}), .b ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, LED_128_Instance_SBox_Instance_5_T1}), .c ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, LED_128_Instance_SBox_Instance_5_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR13_U1 ( .a ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, LED_128_Instance_SBox_Instance_5_L1}), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, LED_128_Instance_SBox_Instance_5_L8}), .c ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, LED_128_Instance_subcells_out[22]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR14_U1 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, LED_128_Instance_SBox_Instance_5_L4}), .b ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, LED_128_Instance_SBox_Instance_5_T3}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, LED_128_Instance_subcells_out[21]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR15_U1 ( .a ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, LED_128_Instance_SBox_Instance_5_L3}), .b ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, LED_128_Instance_SBox_Instance_5_T2}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, LED_128_Instance_subcells_out[20]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_6_U3 ( .x ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, LED_128_Instance_SBox_Instance_6_L0}), .y ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, LED_128_Instance_SBox_Instance_6_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_6_U2 ( .x ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, LED_128_Instance_addconst_out[27]}), .y ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, LED_128_Instance_SBox_Instance_6_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_6_U1 ( .x ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[25]}), .y ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, LED_128_Instance_SBox_Instance_6_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR1_U1 ( .a ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, LED_128_Instance_addconst_out[26]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[25]}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, LED_128_Instance_SBox_Instance_6_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR2_U1 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[25]}), .b ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, LED_128_Instance_addconst_out[24]}), .c ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, LED_128_Instance_SBox_Instance_6_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR3_U1 ( .a ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, LED_128_Instance_SBox_Instance_6_L1}), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, LED_128_Instance_addconst_out[27]}), .c ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, LED_128_Instance_SBox_Instance_6_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_6_XOR16_U1 ( .a ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, LED_128_Instance_SBox_Instance_6_T0}), .b ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, LED_128_Instance_SBox_Instance_6_L2}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, LED_128_Instance_SBox_Instance_6_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR4_U1 ( .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, LED_128_Instance_addconst_out[24]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, LED_128_Instance_SBox_Instance_6_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR5_U1 ( .a ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, LED_128_Instance_SBox_Instance_6_L3}), .b ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, LED_128_Instance_SBox_Instance_6_L0}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, LED_128_Instance_SBox_Instance_6_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR6_U1 ( .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, LED_128_Instance_addconst_out[25]}), .c ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, LED_128_Instance_SBox_Instance_6_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR7_U1 ( .a ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, LED_128_Instance_SBox_Instance_6_T0}), .b ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, LED_128_Instance_SBox_Instance_6_T2}), .c ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, LED_128_Instance_SBox_Instance_6_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_6_XOR8_U1 ( .a ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, LED_128_Instance_SBox_Instance_6_L4}), .b ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, LED_128_Instance_SBox_Instance_6_L5}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, LED_128_Instance_SBox_Instance_6_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR9_U1 ( .a ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, LED_128_Instance_SBox_Instance_6_L1}), .b ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, LED_128_Instance_addconst_out[26]}), .c ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, LED_128_Instance_SBox_Instance_6_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_6_AND1_U1 ( .a ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, LED_128_Instance_SBox_Instance_6_n1}), .b ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, LED_128_Instance_SBox_Instance_6_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[24]), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, LED_128_Instance_SBox_Instance_6_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_6_AND2_U1 ( .a ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, LED_128_Instance_SBox_Instance_6_Q2}), .b ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, LED_128_Instance_SBox_Instance_6_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[25]), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, LED_128_Instance_SBox_Instance_6_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_6_AND3_U1 ( .a ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, LED_128_Instance_SBox_Instance_6_n3}), .b ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, LED_128_Instance_addconst_out[26]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[26]), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, LED_128_Instance_SBox_Instance_6_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_6_AND4_U1 ( .a ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, LED_128_Instance_SBox_Instance_6_Q6}), .b ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, LED_128_Instance_SBox_Instance_6_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[27]), .c ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, LED_128_Instance_SBox_Instance_6_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR10_U1 ( .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, LED_128_Instance_SBox_Instance_6_L5}), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, LED_128_Instance_SBox_Instance_6_T3}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, LED_128_Instance_SBox_Instance_6_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR11_U1 ( .a ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, LED_128_Instance_addconst_out[24]}), .b ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, LED_128_Instance_SBox_Instance_6_L7}), .c ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, LED_128_Instance_subcells_out[27]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR12_U1 ( .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, LED_128_Instance_SBox_Instance_6_L5}), .b ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, LED_128_Instance_SBox_Instance_6_T1}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, LED_128_Instance_SBox_Instance_6_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR13_U1 ( .a ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, LED_128_Instance_SBox_Instance_6_L1}), .b ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, LED_128_Instance_SBox_Instance_6_L8}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, LED_128_Instance_subcells_out[26]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR14_U1 ( .a ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, LED_128_Instance_SBox_Instance_6_L4}), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, LED_128_Instance_SBox_Instance_6_T3}), .c ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, LED_128_Instance_subcells_out[25]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR15_U1 ( .a ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, LED_128_Instance_SBox_Instance_6_L3}), .b ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, LED_128_Instance_SBox_Instance_6_T2}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, LED_128_Instance_subcells_out[24]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_7_U3 ( .x ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, LED_128_Instance_SBox_Instance_7_L0}), .y ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, LED_128_Instance_SBox_Instance_7_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_7_U2 ( .x ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[31]}), .y ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, LED_128_Instance_SBox_Instance_7_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_7_U1 ( .x ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[29]}), .y ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, LED_128_Instance_SBox_Instance_7_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR1_U1 ( .a ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, LED_128_Instance_addconst_out[30]}), .b ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[29]}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, LED_128_Instance_SBox_Instance_7_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR2_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[29]}), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, LED_128_Instance_addconst_out[28]}), .c ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, LED_128_Instance_SBox_Instance_7_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR3_U1 ( .a ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, LED_128_Instance_SBox_Instance_7_L1}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[31]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, LED_128_Instance_SBox_Instance_7_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_7_XOR16_U1 ( .a ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, LED_128_Instance_SBox_Instance_7_T0}), .b ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, LED_128_Instance_SBox_Instance_7_L2}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, LED_128_Instance_SBox_Instance_7_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR4_U1 ( .a ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, LED_128_Instance_addconst_out[28]}), .c ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, LED_128_Instance_SBox_Instance_7_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR5_U1 ( .a ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, LED_128_Instance_SBox_Instance_7_L3}), .b ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, LED_128_Instance_SBox_Instance_7_L0}), .c ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, LED_128_Instance_SBox_Instance_7_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR6_U1 ( .a ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, LED_128_Instance_addconst_out[29]}), .c ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, LED_128_Instance_SBox_Instance_7_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR7_U1 ( .a ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, LED_128_Instance_SBox_Instance_7_T0}), .b ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, LED_128_Instance_SBox_Instance_7_T2}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, LED_128_Instance_SBox_Instance_7_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_7_XOR8_U1 ( .a ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, LED_128_Instance_SBox_Instance_7_L4}), .b ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, LED_128_Instance_SBox_Instance_7_L5}), .c ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, LED_128_Instance_SBox_Instance_7_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR9_U1 ( .a ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, LED_128_Instance_SBox_Instance_7_L1}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, LED_128_Instance_addconst_out[30]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, LED_128_Instance_SBox_Instance_7_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_7_AND1_U1 ( .a ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, LED_128_Instance_SBox_Instance_7_n1}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, LED_128_Instance_SBox_Instance_7_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[28]), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, LED_128_Instance_SBox_Instance_7_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_7_AND2_U1 ( .a ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, LED_128_Instance_SBox_Instance_7_Q2}), .b ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, LED_128_Instance_SBox_Instance_7_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[29]), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, LED_128_Instance_SBox_Instance_7_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_7_AND3_U1 ( .a ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, LED_128_Instance_SBox_Instance_7_n3}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, LED_128_Instance_addconst_out[30]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[30]), .c ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, LED_128_Instance_SBox_Instance_7_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_7_AND4_U1 ( .a ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, LED_128_Instance_SBox_Instance_7_Q6}), .b ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, LED_128_Instance_SBox_Instance_7_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[31]), .c ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, LED_128_Instance_SBox_Instance_7_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR10_U1 ( .a ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, LED_128_Instance_SBox_Instance_7_L5}), .b ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, LED_128_Instance_SBox_Instance_7_T3}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, LED_128_Instance_SBox_Instance_7_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR11_U1 ( .a ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, LED_128_Instance_addconst_out[28]}), .b ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, LED_128_Instance_SBox_Instance_7_L7}), .c ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, LED_128_Instance_subcells_out[31]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR12_U1 ( .a ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, LED_128_Instance_SBox_Instance_7_L5}), .b ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, LED_128_Instance_SBox_Instance_7_T1}), .c ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, LED_128_Instance_SBox_Instance_7_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR13_U1 ( .a ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, LED_128_Instance_SBox_Instance_7_L1}), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, LED_128_Instance_SBox_Instance_7_L8}), .c ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, LED_128_Instance_subcells_out[30]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR14_U1 ( .a ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, LED_128_Instance_SBox_Instance_7_L4}), .b ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, LED_128_Instance_SBox_Instance_7_T3}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, LED_128_Instance_subcells_out[29]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR15_U1 ( .a ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, LED_128_Instance_SBox_Instance_7_L3}), .b ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, LED_128_Instance_SBox_Instance_7_T2}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, LED_128_Instance_subcells_out[28]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_8_U3 ( .x ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, LED_128_Instance_SBox_Instance_8_L0}), .y ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, LED_128_Instance_SBox_Instance_8_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_8_U2 ( .x ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, LED_128_Instance_addconst_out[35]}), .y ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, LED_128_Instance_SBox_Instance_8_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_8_U1 ( .x ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, LED_128_Instance_addconst_out[33]}), .y ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, LED_128_Instance_SBox_Instance_8_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR1_U1 ( .a ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, LED_128_Instance_addconst_out[34]}), .b ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, LED_128_Instance_addconst_out[33]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, LED_128_Instance_SBox_Instance_8_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR2_U1 ( .a ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, LED_128_Instance_addconst_out[33]}), .b ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, LED_128_Instance_addconst_out[32]}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, LED_128_Instance_SBox_Instance_8_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR3_U1 ( .a ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, LED_128_Instance_SBox_Instance_8_L1}), .b ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, LED_128_Instance_addconst_out[35]}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, LED_128_Instance_SBox_Instance_8_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_8_XOR16_U1 ( .a ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, LED_128_Instance_SBox_Instance_8_T0}), .b ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, LED_128_Instance_SBox_Instance_8_L2}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, LED_128_Instance_SBox_Instance_8_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR4_U1 ( .a ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, LED_128_Instance_addconst_out[32]}), .c ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, LED_128_Instance_SBox_Instance_8_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR5_U1 ( .a ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, LED_128_Instance_SBox_Instance_8_L3}), .b ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, LED_128_Instance_SBox_Instance_8_L0}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, LED_128_Instance_SBox_Instance_8_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR6_U1 ( .a ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, LED_128_Instance_addconst_out[33]}), .c ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, LED_128_Instance_SBox_Instance_8_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR7_U1 ( .a ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, LED_128_Instance_SBox_Instance_8_T0}), .b ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, LED_128_Instance_SBox_Instance_8_T2}), .c ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, LED_128_Instance_SBox_Instance_8_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_8_XOR8_U1 ( .a ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, LED_128_Instance_SBox_Instance_8_L4}), .b ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, LED_128_Instance_SBox_Instance_8_L5}), .c ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, LED_128_Instance_SBox_Instance_8_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR9_U1 ( .a ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, LED_128_Instance_SBox_Instance_8_L1}), .b ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, LED_128_Instance_addconst_out[34]}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, LED_128_Instance_SBox_Instance_8_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_8_AND1_U1 ( .a ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, LED_128_Instance_SBox_Instance_8_n1}), .b ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, LED_128_Instance_SBox_Instance_8_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[32]), .c ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, LED_128_Instance_SBox_Instance_8_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_8_AND2_U1 ( .a ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, LED_128_Instance_SBox_Instance_8_Q2}), .b ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, LED_128_Instance_SBox_Instance_8_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[33]), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, LED_128_Instance_SBox_Instance_8_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_8_AND3_U1 ( .a ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, LED_128_Instance_SBox_Instance_8_n3}), .b ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, LED_128_Instance_addconst_out[34]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[34]), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, LED_128_Instance_SBox_Instance_8_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_8_AND4_U1 ( .a ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, LED_128_Instance_SBox_Instance_8_Q6}), .b ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, LED_128_Instance_SBox_Instance_8_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[35]), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, LED_128_Instance_SBox_Instance_8_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR10_U1 ( .a ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, LED_128_Instance_SBox_Instance_8_L5}), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, LED_128_Instance_SBox_Instance_8_T3}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, LED_128_Instance_SBox_Instance_8_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR11_U1 ( .a ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, LED_128_Instance_addconst_out[32]}), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, LED_128_Instance_SBox_Instance_8_L7}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, LED_128_Instance_subcells_out[35]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR12_U1 ( .a ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, LED_128_Instance_SBox_Instance_8_L5}), .b ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, LED_128_Instance_SBox_Instance_8_T1}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, LED_128_Instance_SBox_Instance_8_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR13_U1 ( .a ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, LED_128_Instance_SBox_Instance_8_L1}), .b ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, LED_128_Instance_SBox_Instance_8_L8}), .c ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, LED_128_Instance_subcells_out[34]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR14_U1 ( .a ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, LED_128_Instance_SBox_Instance_8_L4}), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, LED_128_Instance_SBox_Instance_8_T3}), .c ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, LED_128_Instance_subcells_out[33]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR15_U1 ( .a ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, LED_128_Instance_SBox_Instance_8_L3}), .b ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, LED_128_Instance_SBox_Instance_8_T2}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, LED_128_Instance_subcells_out[32]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_9_U3 ( .x ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, LED_128_Instance_SBox_Instance_9_L0}), .y ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, LED_128_Instance_SBox_Instance_9_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_9_U2 ( .x ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, LED_128_Instance_addconst_out[39]}), .y ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, LED_128_Instance_SBox_Instance_9_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_9_U1 ( .x ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, LED_128_Instance_addconst_out[37]}), .y ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, LED_128_Instance_SBox_Instance_9_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR1_U1 ( .a ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, LED_128_Instance_addconst_out[38]}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, LED_128_Instance_addconst_out[37]}), .c ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, LED_128_Instance_SBox_Instance_9_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR2_U1 ( .a ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, LED_128_Instance_addconst_out[37]}), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, LED_128_Instance_addconst_out[36]}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, LED_128_Instance_SBox_Instance_9_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR3_U1 ( .a ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, LED_128_Instance_SBox_Instance_9_L1}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, LED_128_Instance_addconst_out[39]}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, LED_128_Instance_SBox_Instance_9_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_9_XOR16_U1 ( .a ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, LED_128_Instance_SBox_Instance_9_T0}), .b ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, LED_128_Instance_SBox_Instance_9_L2}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, LED_128_Instance_SBox_Instance_9_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR4_U1 ( .a ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, LED_128_Instance_addconst_out[36]}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, LED_128_Instance_SBox_Instance_9_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR5_U1 ( .a ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, LED_128_Instance_SBox_Instance_9_L3}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, LED_128_Instance_SBox_Instance_9_L0}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, LED_128_Instance_SBox_Instance_9_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR6_U1 ( .a ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, LED_128_Instance_addconst_out[37]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, LED_128_Instance_SBox_Instance_9_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR7_U1 ( .a ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, LED_128_Instance_SBox_Instance_9_T0}), .b ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, LED_128_Instance_SBox_Instance_9_T2}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, LED_128_Instance_SBox_Instance_9_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_9_XOR8_U1 ( .a ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, LED_128_Instance_SBox_Instance_9_L4}), .b ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, LED_128_Instance_SBox_Instance_9_L5}), .c ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, LED_128_Instance_SBox_Instance_9_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR9_U1 ( .a ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, LED_128_Instance_SBox_Instance_9_L1}), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, LED_128_Instance_addconst_out[38]}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, LED_128_Instance_SBox_Instance_9_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_9_AND1_U1 ( .a ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, LED_128_Instance_SBox_Instance_9_n1}), .b ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, LED_128_Instance_SBox_Instance_9_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[36]), .c ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, LED_128_Instance_SBox_Instance_9_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_9_AND2_U1 ( .a ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, LED_128_Instance_SBox_Instance_9_Q2}), .b ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, LED_128_Instance_SBox_Instance_9_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[37]), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, LED_128_Instance_SBox_Instance_9_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_9_AND3_U1 ( .a ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, LED_128_Instance_SBox_Instance_9_n3}), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, LED_128_Instance_addconst_out[38]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[38]), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, LED_128_Instance_SBox_Instance_9_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_9_AND4_U1 ( .a ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, LED_128_Instance_SBox_Instance_9_Q6}), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, LED_128_Instance_SBox_Instance_9_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[39]), .c ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, LED_128_Instance_SBox_Instance_9_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR10_U1 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, LED_128_Instance_SBox_Instance_9_L5}), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, LED_128_Instance_SBox_Instance_9_T3}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, LED_128_Instance_SBox_Instance_9_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR11_U1 ( .a ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, LED_128_Instance_addconst_out[36]}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, LED_128_Instance_SBox_Instance_9_L7}), .c ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, LED_128_Instance_subcells_out[39]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR12_U1 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, LED_128_Instance_SBox_Instance_9_L5}), .b ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, LED_128_Instance_SBox_Instance_9_T1}), .c ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, LED_128_Instance_SBox_Instance_9_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR13_U1 ( .a ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, LED_128_Instance_SBox_Instance_9_L1}), .b ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, LED_128_Instance_SBox_Instance_9_L8}), .c ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, LED_128_Instance_subcells_out[38]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR14_U1 ( .a ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, LED_128_Instance_SBox_Instance_9_L4}), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, LED_128_Instance_SBox_Instance_9_T3}), .c ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, LED_128_Instance_subcells_out[37]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR15_U1 ( .a ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, LED_128_Instance_SBox_Instance_9_L3}), .b ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, LED_128_Instance_SBox_Instance_9_T2}), .c ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, LED_128_Instance_subcells_out[36]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_10_U3 ( .x ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, LED_128_Instance_SBox_Instance_10_L0}), .y ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, LED_128_Instance_SBox_Instance_10_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_10_U2 ( .x ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, LED_128_Instance_addconst_out[43]}), .y ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, LED_128_Instance_SBox_Instance_10_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_10_U1 ( .x ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, LED_128_Instance_addconst_out[41]}), .y ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, LED_128_Instance_SBox_Instance_10_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR1_U1 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, LED_128_Instance_addconst_out[42]}), .b ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, LED_128_Instance_addconst_out[41]}), .c ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, LED_128_Instance_SBox_Instance_10_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR2_U1 ( .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, LED_128_Instance_addconst_out[41]}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, LED_128_Instance_addconst_out[40]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, LED_128_Instance_SBox_Instance_10_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR3_U1 ( .a ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, LED_128_Instance_SBox_Instance_10_L1}), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, LED_128_Instance_addconst_out[43]}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, LED_128_Instance_SBox_Instance_10_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_10_XOR16_U1 ( .a ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, LED_128_Instance_SBox_Instance_10_T0}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, LED_128_Instance_SBox_Instance_10_L2}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, LED_128_Instance_SBox_Instance_10_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR4_U1 ( .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, LED_128_Instance_addconst_out[40]}), .c ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, LED_128_Instance_SBox_Instance_10_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR5_U1 ( .a ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, LED_128_Instance_SBox_Instance_10_L3}), .b ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, LED_128_Instance_SBox_Instance_10_L0}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, LED_128_Instance_SBox_Instance_10_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR6_U1 ( .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, LED_128_Instance_addconst_out[41]}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, LED_128_Instance_SBox_Instance_10_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR7_U1 ( .a ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, LED_128_Instance_SBox_Instance_10_T0}), .b ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, LED_128_Instance_SBox_Instance_10_T2}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, LED_128_Instance_SBox_Instance_10_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_10_XOR8_U1 ( .a ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, LED_128_Instance_SBox_Instance_10_L4}), .b ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, LED_128_Instance_SBox_Instance_10_L5}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, LED_128_Instance_SBox_Instance_10_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR9_U1 ( .a ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, LED_128_Instance_SBox_Instance_10_L1}), .b ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, LED_128_Instance_addconst_out[42]}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, LED_128_Instance_SBox_Instance_10_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_10_AND1_U1 ( .a ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, LED_128_Instance_SBox_Instance_10_n1}), .b ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, LED_128_Instance_SBox_Instance_10_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[40]), .c ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, LED_128_Instance_SBox_Instance_10_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_10_AND2_U1 ( .a ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, LED_128_Instance_SBox_Instance_10_Q2}), .b ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, LED_128_Instance_SBox_Instance_10_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[41]), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, LED_128_Instance_SBox_Instance_10_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_10_AND3_U1 ( .a ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, LED_128_Instance_SBox_Instance_10_n3}), .b ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, LED_128_Instance_addconst_out[42]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[42]), .c ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, LED_128_Instance_SBox_Instance_10_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_10_AND4_U1 ( .a ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, LED_128_Instance_SBox_Instance_10_Q6}), .b ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, LED_128_Instance_SBox_Instance_10_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[43]), .c ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, LED_128_Instance_SBox_Instance_10_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR10_U1 ( .a ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, LED_128_Instance_SBox_Instance_10_L5}), .b ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, LED_128_Instance_SBox_Instance_10_T3}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, LED_128_Instance_SBox_Instance_10_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR11_U1 ( .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, LED_128_Instance_addconst_out[40]}), .b ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, LED_128_Instance_SBox_Instance_10_L7}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[43]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR12_U1 ( .a ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, LED_128_Instance_SBox_Instance_10_L5}), .b ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, LED_128_Instance_SBox_Instance_10_T1}), .c ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, LED_128_Instance_SBox_Instance_10_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR13_U1 ( .a ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, LED_128_Instance_SBox_Instance_10_L1}), .b ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, LED_128_Instance_SBox_Instance_10_L8}), .c ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, LED_128_Instance_subcells_out[42]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR14_U1 ( .a ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, LED_128_Instance_SBox_Instance_10_L4}), .b ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, LED_128_Instance_SBox_Instance_10_T3}), .c ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, LED_128_Instance_subcells_out[41]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR15_U1 ( .a ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, LED_128_Instance_SBox_Instance_10_L3}), .b ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, LED_128_Instance_SBox_Instance_10_T2}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, LED_128_Instance_subcells_out[40]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_11_U3 ( .x ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, LED_128_Instance_SBox_Instance_11_L0}), .y ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, LED_128_Instance_SBox_Instance_11_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_11_U2 ( .x ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, LED_128_Instance_addconst_out[47]}), .y ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, LED_128_Instance_SBox_Instance_11_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_11_U1 ( .x ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, LED_128_Instance_addconst_out[45]}), .y ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, LED_128_Instance_SBox_Instance_11_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR1_U1 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, LED_128_Instance_addconst_out[46]}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, LED_128_Instance_addconst_out[45]}), .c ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, LED_128_Instance_SBox_Instance_11_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR2_U1 ( .a ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, LED_128_Instance_addconst_out[45]}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, LED_128_Instance_addconst_out[44]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, LED_128_Instance_SBox_Instance_11_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR3_U1 ( .a ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, LED_128_Instance_SBox_Instance_11_L1}), .b ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, LED_128_Instance_addconst_out[47]}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, LED_128_Instance_SBox_Instance_11_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_11_XOR16_U1 ( .a ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, LED_128_Instance_SBox_Instance_11_T0}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, LED_128_Instance_SBox_Instance_11_L2}), .c ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, LED_128_Instance_SBox_Instance_11_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR4_U1 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, LED_128_Instance_addconst_out[44]}), .c ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, LED_128_Instance_SBox_Instance_11_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR5_U1 ( .a ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, LED_128_Instance_SBox_Instance_11_L3}), .b ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, LED_128_Instance_SBox_Instance_11_L0}), .c ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, LED_128_Instance_SBox_Instance_11_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR6_U1 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, LED_128_Instance_addconst_out[45]}), .c ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, LED_128_Instance_SBox_Instance_11_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR7_U1 ( .a ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, LED_128_Instance_SBox_Instance_11_T0}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, LED_128_Instance_SBox_Instance_11_T2}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, LED_128_Instance_SBox_Instance_11_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_11_XOR8_U1 ( .a ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, LED_128_Instance_SBox_Instance_11_L4}), .b ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, LED_128_Instance_SBox_Instance_11_L5}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, LED_128_Instance_SBox_Instance_11_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR9_U1 ( .a ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, LED_128_Instance_SBox_Instance_11_L1}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, LED_128_Instance_addconst_out[46]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, LED_128_Instance_SBox_Instance_11_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_11_AND1_U1 ( .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, LED_128_Instance_SBox_Instance_11_n1}), .b ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, LED_128_Instance_SBox_Instance_11_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[44]), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, LED_128_Instance_SBox_Instance_11_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_11_AND2_U1 ( .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, LED_128_Instance_SBox_Instance_11_Q2}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, LED_128_Instance_SBox_Instance_11_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[45]), .c ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, LED_128_Instance_SBox_Instance_11_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_11_AND3_U1 ( .a ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, LED_128_Instance_SBox_Instance_11_n3}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, LED_128_Instance_addconst_out[46]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[46]), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, LED_128_Instance_SBox_Instance_11_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_11_AND4_U1 ( .a ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, LED_128_Instance_SBox_Instance_11_Q6}), .b ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, LED_128_Instance_SBox_Instance_11_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[47]), .c ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, LED_128_Instance_SBox_Instance_11_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR10_U1 ( .a ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, LED_128_Instance_SBox_Instance_11_L5}), .b ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, LED_128_Instance_SBox_Instance_11_T3}), .c ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, LED_128_Instance_SBox_Instance_11_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR11_U1 ( .a ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, LED_128_Instance_addconst_out[44]}), .b ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, LED_128_Instance_SBox_Instance_11_L7}), .c ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, LED_128_Instance_subcells_out[47]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR12_U1 ( .a ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, LED_128_Instance_SBox_Instance_11_L5}), .b ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, LED_128_Instance_SBox_Instance_11_T1}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, LED_128_Instance_SBox_Instance_11_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR13_U1 ( .a ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, LED_128_Instance_SBox_Instance_11_L1}), .b ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, LED_128_Instance_SBox_Instance_11_L8}), .c ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, LED_128_Instance_subcells_out[46]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR14_U1 ( .a ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, LED_128_Instance_SBox_Instance_11_L4}), .b ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, LED_128_Instance_SBox_Instance_11_T3}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, LED_128_Instance_subcells_out[45]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR15_U1 ( .a ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, LED_128_Instance_SBox_Instance_11_L3}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, LED_128_Instance_SBox_Instance_11_T2}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, LED_128_Instance_subcells_out[44]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_12_U3 ( .x ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, LED_128_Instance_SBox_Instance_12_L0}), .y ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, LED_128_Instance_SBox_Instance_12_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_12_U2 ( .x ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, LED_128_Instance_addconst_out[51]}), .y ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, LED_128_Instance_SBox_Instance_12_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_12_U1 ( .x ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, LED_128_Instance_addconst_out[49]}), .y ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, LED_128_Instance_SBox_Instance_12_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR1_U1 ( .a ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, LED_128_Instance_addconst_out[50]}), .b ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, LED_128_Instance_addconst_out[49]}), .c ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, LED_128_Instance_SBox_Instance_12_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR2_U1 ( .a ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, LED_128_Instance_addconst_out[49]}), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, LED_128_Instance_addconst_out[48]}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, LED_128_Instance_SBox_Instance_12_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR3_U1 ( .a ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, LED_128_Instance_SBox_Instance_12_L1}), .b ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, LED_128_Instance_addconst_out[51]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, LED_128_Instance_SBox_Instance_12_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_12_XOR16_U1 ( .a ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, LED_128_Instance_SBox_Instance_12_T0}), .b ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, LED_128_Instance_SBox_Instance_12_L2}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, LED_128_Instance_SBox_Instance_12_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR4_U1 ( .a ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, LED_128_Instance_addconst_out[48]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, LED_128_Instance_SBox_Instance_12_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR5_U1 ( .a ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, LED_128_Instance_SBox_Instance_12_L3}), .b ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, LED_128_Instance_SBox_Instance_12_L0}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, LED_128_Instance_SBox_Instance_12_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR6_U1 ( .a ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, LED_128_Instance_addconst_out[49]}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, LED_128_Instance_SBox_Instance_12_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR7_U1 ( .a ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, LED_128_Instance_SBox_Instance_12_T0}), .b ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, LED_128_Instance_SBox_Instance_12_T2}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, LED_128_Instance_SBox_Instance_12_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_12_XOR8_U1 ( .a ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, LED_128_Instance_SBox_Instance_12_L4}), .b ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, LED_128_Instance_SBox_Instance_12_L5}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, LED_128_Instance_SBox_Instance_12_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR9_U1 ( .a ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, LED_128_Instance_SBox_Instance_12_L1}), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, LED_128_Instance_addconst_out[50]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, LED_128_Instance_SBox_Instance_12_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_12_AND1_U1 ( .a ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, LED_128_Instance_SBox_Instance_12_n1}), .b ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, LED_128_Instance_SBox_Instance_12_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[48]), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, LED_128_Instance_SBox_Instance_12_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_12_AND2_U1 ( .a ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, LED_128_Instance_SBox_Instance_12_Q2}), .b ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, LED_128_Instance_SBox_Instance_12_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[49]), .c ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, LED_128_Instance_SBox_Instance_12_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_12_AND3_U1 ( .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, LED_128_Instance_SBox_Instance_12_n3}), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, LED_128_Instance_addconst_out[50]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[50]), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, LED_128_Instance_SBox_Instance_12_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_12_AND4_U1 ( .a ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, LED_128_Instance_SBox_Instance_12_Q6}), .b ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, LED_128_Instance_SBox_Instance_12_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[51]), .c ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, LED_128_Instance_SBox_Instance_12_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR10_U1 ( .a ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, LED_128_Instance_SBox_Instance_12_L5}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, LED_128_Instance_SBox_Instance_12_T3}), .c ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, LED_128_Instance_SBox_Instance_12_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR11_U1 ( .a ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, LED_128_Instance_addconst_out[48]}), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, LED_128_Instance_SBox_Instance_12_L7}), .c ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, LED_128_Instance_subcells_out[51]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR12_U1 ( .a ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, LED_128_Instance_SBox_Instance_12_L5}), .b ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, LED_128_Instance_SBox_Instance_12_T1}), .c ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, LED_128_Instance_SBox_Instance_12_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR13_U1 ( .a ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, LED_128_Instance_SBox_Instance_12_L1}), .b ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, LED_128_Instance_SBox_Instance_12_L8}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, LED_128_Instance_subcells_out[50]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR14_U1 ( .a ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, LED_128_Instance_SBox_Instance_12_L4}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, LED_128_Instance_SBox_Instance_12_T3}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, LED_128_Instance_subcells_out[49]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR15_U1 ( .a ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, LED_128_Instance_SBox_Instance_12_L3}), .b ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, LED_128_Instance_SBox_Instance_12_T2}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, LED_128_Instance_subcells_out[48]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_13_U3 ( .x ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, LED_128_Instance_SBox_Instance_13_L0}), .y ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, LED_128_Instance_SBox_Instance_13_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_13_U2 ( .x ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, LED_128_Instance_addconst_out[55]}), .y ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, LED_128_Instance_SBox_Instance_13_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_13_U1 ( .x ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, LED_128_Instance_addconst_out[53]}), .y ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, LED_128_Instance_SBox_Instance_13_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR1_U1 ( .a ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, LED_128_Instance_addconst_out[54]}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, LED_128_Instance_addconst_out[53]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, LED_128_Instance_SBox_Instance_13_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR2_U1 ( .a ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, LED_128_Instance_addconst_out[53]}), .b ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, LED_128_Instance_addconst_out[52]}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, LED_128_Instance_SBox_Instance_13_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR3_U1 ( .a ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, LED_128_Instance_SBox_Instance_13_L1}), .b ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, LED_128_Instance_addconst_out[55]}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, LED_128_Instance_SBox_Instance_13_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_13_XOR16_U1 ( .a ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, LED_128_Instance_SBox_Instance_13_T0}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, LED_128_Instance_SBox_Instance_13_L2}), .c ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, LED_128_Instance_SBox_Instance_13_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR4_U1 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, LED_128_Instance_addconst_out[52]}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, LED_128_Instance_SBox_Instance_13_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR5_U1 ( .a ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, LED_128_Instance_SBox_Instance_13_L3}), .b ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, LED_128_Instance_SBox_Instance_13_L0}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, LED_128_Instance_SBox_Instance_13_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR6_U1 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, LED_128_Instance_addconst_out[53]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, LED_128_Instance_SBox_Instance_13_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR7_U1 ( .a ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, LED_128_Instance_SBox_Instance_13_T0}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, LED_128_Instance_SBox_Instance_13_T2}), .c ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, LED_128_Instance_SBox_Instance_13_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_13_XOR8_U1 ( .a ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, LED_128_Instance_SBox_Instance_13_L4}), .b ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, LED_128_Instance_SBox_Instance_13_L5}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, LED_128_Instance_SBox_Instance_13_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR9_U1 ( .a ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, LED_128_Instance_SBox_Instance_13_L1}), .b ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, LED_128_Instance_addconst_out[54]}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, LED_128_Instance_SBox_Instance_13_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_13_AND1_U1 ( .a ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, LED_128_Instance_SBox_Instance_13_n1}), .b ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, LED_128_Instance_SBox_Instance_13_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[52]), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, LED_128_Instance_SBox_Instance_13_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_13_AND2_U1 ( .a ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, LED_128_Instance_SBox_Instance_13_Q2}), .b ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, LED_128_Instance_SBox_Instance_13_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[53]), .c ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, LED_128_Instance_SBox_Instance_13_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_13_AND3_U1 ( .a ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, LED_128_Instance_SBox_Instance_13_n3}), .b ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, LED_128_Instance_addconst_out[54]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[54]), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, LED_128_Instance_SBox_Instance_13_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_13_AND4_U1 ( .a ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, LED_128_Instance_SBox_Instance_13_Q6}), .b ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, LED_128_Instance_SBox_Instance_13_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[55]), .c ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, LED_128_Instance_SBox_Instance_13_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR10_U1 ( .a ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, LED_128_Instance_SBox_Instance_13_L5}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, LED_128_Instance_SBox_Instance_13_T3}), .c ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, LED_128_Instance_SBox_Instance_13_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR11_U1 ( .a ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, LED_128_Instance_addconst_out[52]}), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, LED_128_Instance_SBox_Instance_13_L7}), .c ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, LED_128_Instance_subcells_out[55]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR12_U1 ( .a ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, LED_128_Instance_SBox_Instance_13_L5}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, LED_128_Instance_SBox_Instance_13_T1}), .c ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, LED_128_Instance_SBox_Instance_13_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR13_U1 ( .a ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, LED_128_Instance_SBox_Instance_13_L1}), .b ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, LED_128_Instance_SBox_Instance_13_L8}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, LED_128_Instance_subcells_out[54]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR14_U1 ( .a ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, LED_128_Instance_SBox_Instance_13_L4}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, LED_128_Instance_SBox_Instance_13_T3}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, LED_128_Instance_subcells_out[53]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR15_U1 ( .a ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, LED_128_Instance_SBox_Instance_13_L3}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, LED_128_Instance_SBox_Instance_13_T2}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, LED_128_Instance_subcells_out[52]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_14_U3 ( .x ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, LED_128_Instance_SBox_Instance_14_L0}), .y ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, LED_128_Instance_SBox_Instance_14_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_14_U2 ( .x ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, LED_128_Instance_addconst_out[59]}), .y ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, LED_128_Instance_SBox_Instance_14_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_14_U1 ( .x ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, LED_128_Instance_addconst_out[57]}), .y ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, LED_128_Instance_SBox_Instance_14_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR1_U1 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, LED_128_Instance_addconst_out[58]}), .b ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, LED_128_Instance_addconst_out[57]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, LED_128_Instance_SBox_Instance_14_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR2_U1 ( .a ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, LED_128_Instance_addconst_out[57]}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, LED_128_Instance_addconst_out[56]}), .c ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, LED_128_Instance_SBox_Instance_14_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR3_U1 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, LED_128_Instance_SBox_Instance_14_L1}), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, LED_128_Instance_addconst_out[59]}), .c ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, LED_128_Instance_SBox_Instance_14_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_14_XOR16_U1 ( .a ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, LED_128_Instance_SBox_Instance_14_T0}), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, LED_128_Instance_SBox_Instance_14_L2}), .c ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, LED_128_Instance_SBox_Instance_14_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR4_U1 ( .a ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, LED_128_Instance_addconst_out[56]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, LED_128_Instance_SBox_Instance_14_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR5_U1 ( .a ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, LED_128_Instance_SBox_Instance_14_L3}), .b ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, LED_128_Instance_SBox_Instance_14_L0}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, LED_128_Instance_SBox_Instance_14_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR6_U1 ( .a ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, LED_128_Instance_addconst_out[57]}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, LED_128_Instance_SBox_Instance_14_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR7_U1 ( .a ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, LED_128_Instance_SBox_Instance_14_T0}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, LED_128_Instance_SBox_Instance_14_T2}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, LED_128_Instance_SBox_Instance_14_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_14_XOR8_U1 ( .a ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, LED_128_Instance_SBox_Instance_14_L4}), .b ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, LED_128_Instance_SBox_Instance_14_L5}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, LED_128_Instance_SBox_Instance_14_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR9_U1 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, LED_128_Instance_SBox_Instance_14_L1}), .b ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, LED_128_Instance_addconst_out[58]}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, LED_128_Instance_SBox_Instance_14_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_14_AND1_U1 ( .a ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, LED_128_Instance_SBox_Instance_14_n1}), .b ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, LED_128_Instance_SBox_Instance_14_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[56]), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, LED_128_Instance_SBox_Instance_14_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_14_AND2_U1 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, LED_128_Instance_SBox_Instance_14_Q2}), .b ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, LED_128_Instance_SBox_Instance_14_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[57]), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, LED_128_Instance_SBox_Instance_14_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_14_AND3_U1 ( .a ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, LED_128_Instance_SBox_Instance_14_n3}), .b ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, LED_128_Instance_addconst_out[58]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[58]), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, LED_128_Instance_SBox_Instance_14_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_14_AND4_U1 ( .a ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, LED_128_Instance_SBox_Instance_14_Q6}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, LED_128_Instance_SBox_Instance_14_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[59]), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, LED_128_Instance_SBox_Instance_14_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR10_U1 ( .a ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, LED_128_Instance_SBox_Instance_14_L5}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, LED_128_Instance_SBox_Instance_14_T3}), .c ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, LED_128_Instance_SBox_Instance_14_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR11_U1 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, LED_128_Instance_addconst_out[56]}), .b ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, LED_128_Instance_SBox_Instance_14_L7}), .c ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, LED_128_Instance_subcells_out[59]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR12_U1 ( .a ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, LED_128_Instance_SBox_Instance_14_L5}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, LED_128_Instance_SBox_Instance_14_T1}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, LED_128_Instance_SBox_Instance_14_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR13_U1 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, LED_128_Instance_SBox_Instance_14_L1}), .b ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, LED_128_Instance_SBox_Instance_14_L8}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, LED_128_Instance_subcells_out[58]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR14_U1 ( .a ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, LED_128_Instance_SBox_Instance_14_L4}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, LED_128_Instance_SBox_Instance_14_T3}), .c ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, LED_128_Instance_subcells_out[57]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR15_U1 ( .a ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, LED_128_Instance_SBox_Instance_14_L3}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, LED_128_Instance_SBox_Instance_14_T2}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, LED_128_Instance_subcells_out[56]}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_15_U3 ( .x ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, LED_128_Instance_SBox_Instance_15_L0}), .y ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, LED_128_Instance_SBox_Instance_15_n1}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_15_U2 ( .x ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, LED_128_Instance_addconst_out[63]}), .y ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, LED_128_Instance_SBox_Instance_15_n2}) ) ;
    not_LMDPL LED_128_Instance_SBox_Instance_15_U1 ( .x ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, LED_128_Instance_addconst_out[61]}), .y ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, LED_128_Instance_SBox_Instance_15_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR1_U1 ( .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, LED_128_Instance_addconst_out[62]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, LED_128_Instance_addconst_out[61]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, LED_128_Instance_SBox_Instance_15_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR2_U1 ( .a ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, LED_128_Instance_addconst_out[61]}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, LED_128_Instance_addconst_out[60]}), .c ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, LED_128_Instance_SBox_Instance_15_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR3_U1 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, LED_128_Instance_SBox_Instance_15_L1}), .b ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, LED_128_Instance_addconst_out[63]}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, LED_128_Instance_SBox_Instance_15_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_15_XOR16_U1 ( .a ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, LED_128_Instance_SBox_Instance_15_T0}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, LED_128_Instance_SBox_Instance_15_L2}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, LED_128_Instance_SBox_Instance_15_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR4_U1 ( .a ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, LED_128_Instance_addconst_out[60]}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, LED_128_Instance_SBox_Instance_15_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR5_U1 ( .a ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, LED_128_Instance_SBox_Instance_15_L3}), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, LED_128_Instance_SBox_Instance_15_L0}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, LED_128_Instance_SBox_Instance_15_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR6_U1 ( .a ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, LED_128_Instance_addconst_out[61]}), .c ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, LED_128_Instance_SBox_Instance_15_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR7_U1 ( .a ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, LED_128_Instance_SBox_Instance_15_T0}), .b ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, LED_128_Instance_SBox_Instance_15_T2}), .c ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, LED_128_Instance_SBox_Instance_15_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_SBox_Instance_15_XOR8_U1 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, LED_128_Instance_SBox_Instance_15_L4}), .b ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, LED_128_Instance_SBox_Instance_15_L5}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, LED_128_Instance_SBox_Instance_15_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR9_U1 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, LED_128_Instance_SBox_Instance_15_L1}), .b ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, LED_128_Instance_addconst_out[62]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, LED_128_Instance_SBox_Instance_15_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_15_AND1_U1 ( .a ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, LED_128_Instance_SBox_Instance_15_n1}), .b ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, LED_128_Instance_SBox_Instance_15_n2}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[60]), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, LED_128_Instance_SBox_Instance_15_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_15_AND2_U1 ( .a ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, LED_128_Instance_SBox_Instance_15_Q2}), .b ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, LED_128_Instance_SBox_Instance_15_Q3}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[61]), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, LED_128_Instance_SBox_Instance_15_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_15_AND3_U1 ( .a ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, LED_128_Instance_SBox_Instance_15_n3}), .b ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, LED_128_Instance_addconst_out[62]}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[62]), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, LED_128_Instance_SBox_Instance_15_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) LED_128_Instance_SBox_Instance_15_AND4_U1 ( .a ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, LED_128_Instance_SBox_Instance_15_Q6}), .b ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, LED_128_Instance_SBox_Instance_15_Q7}), .mid_rst (mid_rst), .clk (CLK), .r (Fresh[63]), .c ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, LED_128_Instance_SBox_Instance_15_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR10_U1 ( .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, LED_128_Instance_SBox_Instance_15_L5}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, LED_128_Instance_SBox_Instance_15_T3}), .c ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, LED_128_Instance_SBox_Instance_15_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR11_U1 ( .a ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, LED_128_Instance_addconst_out[60]}), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, LED_128_Instance_SBox_Instance_15_L7}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, LED_128_Instance_subcells_out[63]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR12_U1 ( .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, LED_128_Instance_SBox_Instance_15_L5}), .b ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, LED_128_Instance_SBox_Instance_15_T1}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, LED_128_Instance_SBox_Instance_15_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR13_U1 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, LED_128_Instance_SBox_Instance_15_L1}), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, LED_128_Instance_SBox_Instance_15_L8}), .c ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, LED_128_Instance_subcells_out[62]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR14_U1 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, LED_128_Instance_SBox_Instance_15_L4}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, LED_128_Instance_SBox_Instance_15_T3}), .c ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, LED_128_Instance_subcells_out[61]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR15_U1 ( .a ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, LED_128_Instance_SBox_Instance_15_L3}), .b ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, LED_128_Instance_SBox_Instance_15_T2}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, LED_128_Instance_subcells_out[60]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U54 ( .a ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, LED_128_Instance_MCS_Instance_0_n38}), .b ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, LED_128_Instance_MCS_Instance_0_n37}), .c ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, LED_128_Instance_mixcolumns_out[51]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U53 ( .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, LED_128_Instance_MCS_Instance_0_n37}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U52 ( .a ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, LED_128_Instance_mixcolumns_out[34]}), .b ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, LED_128_Instance_mixcolumns_out[18]}), .c ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, LED_128_Instance_MCS_Instance_0_n38}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U51 ( .a ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, LED_128_Instance_MCS_Instance_0_n36}), .b ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, LED_128_Instance_mixcolumns_out[34]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U50 ( .a ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, LED_128_Instance_MCS_Instance_0_n34}), .c ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, LED_128_Instance_MCS_Instance_0_n36}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U49 ( .a ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, LED_128_Instance_MCS_Instance_0_n33}), .b ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, LED_128_Instance_mixcolumns_out[33]}), .c ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, LED_128_Instance_mixcolumns_out[50]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U48 ( .a ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[2]}), .b ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, LED_128_Instance_MCS_Instance_0_n33}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U47 ( .a ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, LED_128_Instance_MCS_Instance_0_n32}), .b ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, LED_128_Instance_MCS_Instance_0_n31}), .c ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, LED_128_Instance_mixcolumns_out[49]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U46 ( .a ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, LED_128_Instance_MCS_Instance_0_n30}), .b ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, LED_128_Instance_MCS_Instance_0_n29}), .c ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, LED_128_Instance_MCS_Instance_0_n32}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U45 ( .a ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, LED_128_Instance_mixcolumns_out[1]}), .c ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, LED_128_Instance_MCS_Instance_0_n29}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U44 ( .a ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, LED_128_Instance_mixcolumns_out[32]}), .b ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, LED_128_Instance_MCS_Instance_0_n28}), .c ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, LED_128_Instance_MCS_Instance_0_n30}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U43 ( .a ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, LED_128_Instance_MCS_Instance_0_n27}), .b ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, LED_128_Instance_MCS_Instance_0_n26}), .c ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, LED_128_Instance_mixcolumns_out[32]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U42 ( .a ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, LED_128_Instance_mixcolumns_out[3]}), .c ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, LED_128_Instance_MCS_Instance_0_n26}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U41 ( .a ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, LED_128_Instance_subcells_out[60]}), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, LED_128_Instance_mixcolumns_out[19]}), .c ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, LED_128_Instance_MCS_Instance_0_n27}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U40 ( .a ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, LED_128_Instance_MCS_Instance_0_n25}), .b ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, LED_128_Instance_mixcolumns_out[0]}), .c ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, LED_128_Instance_mixcolumns_out[48]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U39 ( .a ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, LED_128_Instance_mixcolumns_out[19]}), .b ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, LED_128_Instance_MCS_Instance_0_n28}), .c ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, LED_128_Instance_MCS_Instance_0_n25}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U38 ( .a ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, LED_128_Instance_mixcolumns_out[35]}), .c ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, LED_128_Instance_MCS_Instance_0_n28}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U37 ( .a ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, LED_128_Instance_MCS_Instance_0_n24}), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, LED_128_Instance_MCS_Instance_0_n23}), .c ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, LED_128_Instance_mixcolumns_out[35]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U36 ( .a ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, LED_128_Instance_subcells_out[41]}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, LED_128_Instance_MCS_Instance_0_n23}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U35 ( .a ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, LED_128_Instance_mixcolumns_out[18]}), .b ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[2]}), .c ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, LED_128_Instance_MCS_Instance_0_n24}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U34 ( .a ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, LED_128_Instance_MCS_Instance_0_n22}), .b ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, LED_128_Instance_MCS_Instance_0_n21}), .c ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, LED_128_Instance_mixcolumns_out[18]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U33 ( .a ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, LED_128_Instance_MCS_Instance_0_n20}), .b ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, LED_128_Instance_MCS_Instance_0_n21}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U32 ( .a ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, LED_128_Instance_mixcolumns_out[1]}), .b ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, LED_128_Instance_subcells_out[20]}), .c ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, LED_128_Instance_MCS_Instance_0_n22}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U31 ( .a ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, LED_128_Instance_MCS_Instance_0_n19}), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, LED_128_Instance_MCS_Instance_0_n18}), .c ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, LED_128_Instance_mixcolumns_out[1]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U30 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, LED_128_Instance_subcells_out[40]}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, LED_128_Instance_MCS_Instance_0_n18}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U29 ( .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, LED_128_Instance_MCS_Instance_0_n17}), .b ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, LED_128_Instance_MCS_Instance_0_n34}), .c ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, LED_128_Instance_MCS_Instance_0_n19}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U28 ( .a ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, LED_128_Instance_MCS_Instance_0_n16}), .b ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, LED_128_Instance_subcells_out[2]}), .c ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, LED_128_Instance_MCS_Instance_0_n34}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U27 ( .a ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, LED_128_Instance_subcells_out[21]}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, LED_128_Instance_subcells_out[3]}), .c ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, LED_128_Instance_MCS_Instance_0_n16}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U26 ( .a ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, LED_128_Instance_MCS_Instance_0_n15}), .b ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, LED_128_Instance_MCS_Instance_0_n31}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, LED_128_Instance_mixcolumns_out[33]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U25 ( .a ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, LED_128_Instance_mixcolumns_out[16]}), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, LED_128_Instance_mixcolumns_out[19]}), .c ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, LED_128_Instance_MCS_Instance_0_n31}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U24 ( .a ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, LED_128_Instance_MCS_Instance_0_n14}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, LED_128_Instance_MCS_Instance_0_n13}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, LED_128_Instance_MCS_Instance_0_n15}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U23 ( .a ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, LED_128_Instance_MCS_Instance_0_n13}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U22 ( .a ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, LED_128_Instance_MCS_Instance_0_n12}), .b ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, LED_128_Instance_MCS_Instance_0_n14}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U21 ( .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, LED_128_Instance_MCS_Instance_0_n11}), .b ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, LED_128_Instance_MCS_Instance_0_n10}), .c ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, LED_128_Instance_mixcolumns_out[16]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U20 ( .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, LED_128_Instance_subcells_out[63]}), .c ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, LED_128_Instance_MCS_Instance_0_n10}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U19 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, LED_128_Instance_subcells_out[40]}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, LED_128_Instance_subcells_out[22]}), .c ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, LED_128_Instance_MCS_Instance_0_n11}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U18 ( .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, LED_128_Instance_MCS_Instance_0_n9}), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, LED_128_Instance_MCS_Instance_0_n8}), .c ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, LED_128_Instance_mixcolumns_out[19]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U17 ( .a ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, LED_128_Instance_MCS_Instance_0_n8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U16 ( .a ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[2]}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, LED_128_Instance_subcells_out[21]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, LED_128_Instance_MCS_Instance_0_n9}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U15 ( .a ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, LED_128_Instance_MCS_Instance_0_n7}), .b ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, LED_128_Instance_MCS_Instance_0_n6}), .c ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, LED_128_Instance_mixcolumns_out[2]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U14 ( .a ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, LED_128_Instance_MCS_Instance_0_n5}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, LED_128_Instance_subcells_out[3]}), .c ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, LED_128_Instance_MCS_Instance_0_n6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U13 ( .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, LED_128_Instance_subcells_out[0]}), .b ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, LED_128_Instance_MCS_Instance_0_n7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U12 ( .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, LED_128_Instance_MCS_Instance_0_n17}), .b ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, LED_128_Instance_mixcolumns_out[17]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U11 ( .a ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, LED_128_Instance_MCS_Instance_0_n4}), .b ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, LED_128_Instance_MCS_Instance_0_n12}), .c ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, LED_128_Instance_MCS_Instance_0_n35}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U10 ( .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, LED_128_Instance_mixcolumns_out[0]}), .c ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, LED_128_Instance_MCS_Instance_0_n12}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U9 ( .a ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, LED_128_Instance_subcells_out[23]}), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, LED_128_Instance_MCS_Instance_0_n5}), .c ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, LED_128_Instance_MCS_Instance_0_n4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U8 ( .a ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, LED_128_Instance_subcells_out[22]}), .b ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, LED_128_Instance_subcells_out[41]}), .c ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, LED_128_Instance_MCS_Instance_0_n5}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U7 ( .a ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, LED_128_Instance_subcells_out[60]}), .c ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, LED_128_Instance_MCS_Instance_0_n17}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U6 ( .a ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, LED_128_Instance_MCS_Instance_0_n3}), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, LED_128_Instance_MCS_Instance_0_n2}), .c ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, LED_128_Instance_mixcolumns_out[0]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U5 ( .a ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, LED_128_Instance_MCS_Instance_0_n2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U4 ( .a ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, LED_128_Instance_subcells_out[2]}), .b ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, LED_128_Instance_subcells_out[20]}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, LED_128_Instance_MCS_Instance_0_n3}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U3 ( .a ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, LED_128_Instance_MCS_Instance_0_n1}), .b ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, LED_128_Instance_subcells_out[62]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, LED_128_Instance_mixcolumns_out[3]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_0_U2 ( .a ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, LED_128_Instance_MCS_Instance_0_n20}), .b ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, LED_128_Instance_subcells_out[1]}), .c ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, LED_128_Instance_MCS_Instance_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_0_U1 ( .a ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, LED_128_Instance_subcells_out[23]}), .c ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, LED_128_Instance_MCS_Instance_0_n20}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U54 ( .a ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, LED_128_Instance_MCS_Instance_1_n38}), .b ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, LED_128_Instance_MCS_Instance_1_n37}), .c ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, LED_128_Instance_mixcolumns_out[55]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U53 ( .a ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, LED_128_Instance_MCS_Instance_1_n37}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U52 ( .a ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, LED_128_Instance_mixcolumns_out[38]}), .b ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, LED_128_Instance_mixcolumns_out[22]}), .c ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, LED_128_Instance_MCS_Instance_1_n38}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U51 ( .a ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, LED_128_Instance_MCS_Instance_1_n36}), .b ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, LED_128_Instance_mixcolumns_out[38]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U50 ( .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, LED_128_Instance_MCS_Instance_1_n34}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, LED_128_Instance_MCS_Instance_1_n36}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U49 ( .a ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, LED_128_Instance_MCS_Instance_1_n33}), .b ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, LED_128_Instance_mixcolumns_out[37]}), .c ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, LED_128_Instance_mixcolumns_out[54]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U48 ( .a ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, LED_128_Instance_mixcolumns_out[6]}), .b ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, LED_128_Instance_MCS_Instance_1_n33}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U47 ( .a ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, LED_128_Instance_MCS_Instance_1_n32}), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, LED_128_Instance_MCS_Instance_1_n31}), .c ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, LED_128_Instance_mixcolumns_out[53]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U46 ( .a ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, LED_128_Instance_MCS_Instance_1_n30}), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, LED_128_Instance_MCS_Instance_1_n29}), .c ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, LED_128_Instance_MCS_Instance_1_n32}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U45 ( .a ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, LED_128_Instance_mixcolumns_out[5]}), .c ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, LED_128_Instance_MCS_Instance_1_n29}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U44 ( .a ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, LED_128_Instance_mixcolumns_out[36]}), .b ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, LED_128_Instance_MCS_Instance_1_n28}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, LED_128_Instance_MCS_Instance_1_n30}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U43 ( .a ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, LED_128_Instance_MCS_Instance_1_n27}), .b ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, LED_128_Instance_MCS_Instance_1_n26}), .c ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, LED_128_Instance_mixcolumns_out[36]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U42 ( .a ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, LED_128_Instance_mixcolumns_out[7]}), .c ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, LED_128_Instance_MCS_Instance_1_n26}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U41 ( .a ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, LED_128_Instance_subcells_out[48]}), .b ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, LED_128_Instance_mixcolumns_out[23]}), .c ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, LED_128_Instance_MCS_Instance_1_n27}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U40 ( .a ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, LED_128_Instance_MCS_Instance_1_n25}), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, LED_128_Instance_mixcolumns_out[4]}), .c ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, LED_128_Instance_mixcolumns_out[52]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U39 ( .a ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, LED_128_Instance_mixcolumns_out[23]}), .b ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, LED_128_Instance_MCS_Instance_1_n28}), .c ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, LED_128_Instance_MCS_Instance_1_n25}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U38 ( .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, LED_128_Instance_mixcolumns_out[39]}), .c ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, LED_128_Instance_MCS_Instance_1_n28}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U37 ( .a ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, LED_128_Instance_MCS_Instance_1_n24}), .b ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, LED_128_Instance_MCS_Instance_1_n23}), .c ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, LED_128_Instance_mixcolumns_out[39]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U36 ( .a ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, LED_128_Instance_subcells_out[45]}), .c ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, LED_128_Instance_MCS_Instance_1_n23}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U35 ( .a ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, LED_128_Instance_mixcolumns_out[22]}), .b ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, LED_128_Instance_mixcolumns_out[6]}), .c ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, LED_128_Instance_MCS_Instance_1_n24}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U34 ( .a ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, LED_128_Instance_MCS_Instance_1_n22}), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, LED_128_Instance_MCS_Instance_1_n21}), .c ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, LED_128_Instance_mixcolumns_out[22]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U33 ( .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, LED_128_Instance_MCS_Instance_1_n20}), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, LED_128_Instance_MCS_Instance_1_n21}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U32 ( .a ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, LED_128_Instance_mixcolumns_out[5]}), .b ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, LED_128_Instance_subcells_out[24]}), .c ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, LED_128_Instance_MCS_Instance_1_n22}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U31 ( .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, LED_128_Instance_MCS_Instance_1_n19}), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, LED_128_Instance_MCS_Instance_1_n18}), .c ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, LED_128_Instance_mixcolumns_out[5]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U30 ( .a ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, LED_128_Instance_subcells_out[44]}), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, LED_128_Instance_MCS_Instance_1_n18}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U29 ( .a ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, LED_128_Instance_MCS_Instance_1_n17}), .b ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, LED_128_Instance_MCS_Instance_1_n34}), .c ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, LED_128_Instance_MCS_Instance_1_n19}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U28 ( .a ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, LED_128_Instance_MCS_Instance_1_n16}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, LED_128_Instance_subcells_out[6]}), .c ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, LED_128_Instance_MCS_Instance_1_n34}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U27 ( .a ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, LED_128_Instance_subcells_out[25]}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, LED_128_Instance_subcells_out[7]}), .c ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, LED_128_Instance_MCS_Instance_1_n16}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U26 ( .a ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, LED_128_Instance_MCS_Instance_1_n15}), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, LED_128_Instance_MCS_Instance_1_n31}), .c ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, LED_128_Instance_mixcolumns_out[37]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U25 ( .a ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, LED_128_Instance_mixcolumns_out[20]}), .b ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, LED_128_Instance_mixcolumns_out[23]}), .c ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, LED_128_Instance_MCS_Instance_1_n31}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U24 ( .a ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, LED_128_Instance_MCS_Instance_1_n14}), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, LED_128_Instance_MCS_Instance_1_n13}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, LED_128_Instance_MCS_Instance_1_n15}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U23 ( .a ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, LED_128_Instance_MCS_Instance_1_n13}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U22 ( .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, LED_128_Instance_MCS_Instance_1_n12}), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, LED_128_Instance_MCS_Instance_1_n14}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U21 ( .a ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, LED_128_Instance_MCS_Instance_1_n11}), .b ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, LED_128_Instance_MCS_Instance_1_n10}), .c ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, LED_128_Instance_mixcolumns_out[20]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U20 ( .a ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, LED_128_Instance_subcells_out[51]}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, LED_128_Instance_MCS_Instance_1_n10}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U19 ( .a ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, LED_128_Instance_subcells_out[44]}), .b ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, LED_128_Instance_subcells_out[26]}), .c ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, LED_128_Instance_MCS_Instance_1_n11}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U18 ( .a ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, LED_128_Instance_MCS_Instance_1_n9}), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, LED_128_Instance_MCS_Instance_1_n8}), .c ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, LED_128_Instance_mixcolumns_out[23]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U17 ( .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, LED_128_Instance_MCS_Instance_1_n8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U16 ( .a ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, LED_128_Instance_mixcolumns_out[6]}), .b ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, LED_128_Instance_subcells_out[25]}), .c ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, LED_128_Instance_MCS_Instance_1_n9}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U15 ( .a ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, LED_128_Instance_MCS_Instance_1_n7}), .b ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, LED_128_Instance_MCS_Instance_1_n6}), .c ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, LED_128_Instance_mixcolumns_out[6]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U14 ( .a ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, LED_128_Instance_MCS_Instance_1_n5}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, LED_128_Instance_subcells_out[7]}), .c ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, LED_128_Instance_MCS_Instance_1_n6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U13 ( .a ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, LED_128_Instance_subcells_out[4]}), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, LED_128_Instance_MCS_Instance_1_n7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U12 ( .a ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, LED_128_Instance_MCS_Instance_1_n17}), .b ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, LED_128_Instance_mixcolumns_out[21]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U11 ( .a ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, LED_128_Instance_MCS_Instance_1_n4}), .b ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, LED_128_Instance_MCS_Instance_1_n12}), .c ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, LED_128_Instance_MCS_Instance_1_n35}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U10 ( .a ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, LED_128_Instance_mixcolumns_out[4]}), .c ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, LED_128_Instance_MCS_Instance_1_n12}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U9 ( .a ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, LED_128_Instance_subcells_out[27]}), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, LED_128_Instance_MCS_Instance_1_n5}), .c ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, LED_128_Instance_MCS_Instance_1_n4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U8 ( .a ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, LED_128_Instance_subcells_out[26]}), .b ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, LED_128_Instance_subcells_out[45]}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, LED_128_Instance_MCS_Instance_1_n5}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U7 ( .a ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, LED_128_Instance_subcells_out[48]}), .c ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, LED_128_Instance_MCS_Instance_1_n17}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U6 ( .a ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, LED_128_Instance_MCS_Instance_1_n3}), .b ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, LED_128_Instance_MCS_Instance_1_n2}), .c ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, LED_128_Instance_mixcolumns_out[4]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U5 ( .a ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, LED_128_Instance_MCS_Instance_1_n2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U4 ( .a ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, LED_128_Instance_subcells_out[6]}), .b ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, LED_128_Instance_subcells_out[24]}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, LED_128_Instance_MCS_Instance_1_n3}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U3 ( .a ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, LED_128_Instance_MCS_Instance_1_n1}), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, LED_128_Instance_subcells_out[50]}), .c ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, LED_128_Instance_mixcolumns_out[7]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_1_U2 ( .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, LED_128_Instance_MCS_Instance_1_n20}), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, LED_128_Instance_subcells_out[5]}), .c ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, LED_128_Instance_MCS_Instance_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_1_U1 ( .a ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, LED_128_Instance_subcells_out[27]}), .c ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, LED_128_Instance_MCS_Instance_1_n20}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U54 ( .a ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, LED_128_Instance_MCS_Instance_2_n38}), .b ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, LED_128_Instance_MCS_Instance_2_n37}), .c ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, LED_128_Instance_mixcolumns_out[59]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U53 ( .a ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, LED_128_Instance_MCS_Instance_2_n37}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U52 ( .a ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, LED_128_Instance_mixcolumns_out[42]}), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, LED_128_Instance_mixcolumns_out[26]}), .c ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, LED_128_Instance_MCS_Instance_2_n38}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U51 ( .a ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, LED_128_Instance_MCS_Instance_2_n36}), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, LED_128_Instance_mixcolumns_out[42]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U50 ( .a ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, LED_128_Instance_MCS_Instance_2_n34}), .c ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, LED_128_Instance_MCS_Instance_2_n36}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U49 ( .a ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, LED_128_Instance_MCS_Instance_2_n33}), .b ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, LED_128_Instance_mixcolumns_out[41]}), .c ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, LED_128_Instance_mixcolumns_out[58]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U48 ( .a ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, LED_128_Instance_mixcolumns_out[10]}), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, LED_128_Instance_MCS_Instance_2_n33}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U47 ( .a ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, LED_128_Instance_MCS_Instance_2_n32}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, LED_128_Instance_MCS_Instance_2_n31}), .c ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, LED_128_Instance_mixcolumns_out[57]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U46 ( .a ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, LED_128_Instance_MCS_Instance_2_n30}), .b ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, LED_128_Instance_MCS_Instance_2_n29}), .c ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, LED_128_Instance_MCS_Instance_2_n32}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U45 ( .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, LED_128_Instance_mixcolumns_out[9]}), .c ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, LED_128_Instance_MCS_Instance_2_n29}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U44 ( .a ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, LED_128_Instance_mixcolumns_out[40]}), .b ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, LED_128_Instance_MCS_Instance_2_n28}), .c ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, LED_128_Instance_MCS_Instance_2_n30}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U43 ( .a ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, LED_128_Instance_MCS_Instance_2_n27}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, LED_128_Instance_MCS_Instance_2_n26}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, LED_128_Instance_mixcolumns_out[40]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U42 ( .a ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, LED_128_Instance_mixcolumns_out[11]}), .c ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, LED_128_Instance_MCS_Instance_2_n26}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U41 ( .a ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, LED_128_Instance_subcells_out[52]}), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, LED_128_Instance_mixcolumns_out[27]}), .c ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, LED_128_Instance_MCS_Instance_2_n27}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U40 ( .a ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, LED_128_Instance_MCS_Instance_2_n25}), .b ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, LED_128_Instance_mixcolumns_out[8]}), .c ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, LED_128_Instance_mixcolumns_out[56]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U39 ( .a ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, LED_128_Instance_mixcolumns_out[27]}), .b ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, LED_128_Instance_MCS_Instance_2_n28}), .c ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, LED_128_Instance_MCS_Instance_2_n25}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U38 ( .a ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, LED_128_Instance_mixcolumns_out[43]}), .c ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, LED_128_Instance_MCS_Instance_2_n28}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U37 ( .a ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, LED_128_Instance_MCS_Instance_2_n24}), .b ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, LED_128_Instance_MCS_Instance_2_n23}), .c ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, LED_128_Instance_mixcolumns_out[43]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U36 ( .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, LED_128_Instance_subcells_out[33]}), .c ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, LED_128_Instance_MCS_Instance_2_n23}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U35 ( .a ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, LED_128_Instance_mixcolumns_out[26]}), .b ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, LED_128_Instance_mixcolumns_out[10]}), .c ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, LED_128_Instance_MCS_Instance_2_n24}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U34 ( .a ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, LED_128_Instance_MCS_Instance_2_n22}), .b ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, LED_128_Instance_MCS_Instance_2_n21}), .c ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, LED_128_Instance_mixcolumns_out[26]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U33 ( .a ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, LED_128_Instance_MCS_Instance_2_n20}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, LED_128_Instance_MCS_Instance_2_n21}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U32 ( .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, LED_128_Instance_mixcolumns_out[9]}), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, LED_128_Instance_subcells_out[28]}), .c ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, LED_128_Instance_MCS_Instance_2_n22}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U31 ( .a ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, LED_128_Instance_MCS_Instance_2_n19}), .b ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, LED_128_Instance_MCS_Instance_2_n18}), .c ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, LED_128_Instance_mixcolumns_out[9]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U30 ( .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, LED_128_Instance_subcells_out[32]}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, LED_128_Instance_MCS_Instance_2_n18}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U29 ( .a ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, LED_128_Instance_MCS_Instance_2_n17}), .b ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, LED_128_Instance_MCS_Instance_2_n34}), .c ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, LED_128_Instance_MCS_Instance_2_n19}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U28 ( .a ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, LED_128_Instance_MCS_Instance_2_n16}), .b ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, LED_128_Instance_subcells_out[10]}), .c ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, LED_128_Instance_MCS_Instance_2_n34}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U27 ( .a ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, LED_128_Instance_subcells_out[29]}), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, LED_128_Instance_subcells_out[11]}), .c ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, LED_128_Instance_MCS_Instance_2_n16}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U26 ( .a ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, LED_128_Instance_MCS_Instance_2_n15}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, LED_128_Instance_MCS_Instance_2_n31}), .c ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, LED_128_Instance_mixcolumns_out[41]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U25 ( .a ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, LED_128_Instance_mixcolumns_out[24]}), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, LED_128_Instance_mixcolumns_out[27]}), .c ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, LED_128_Instance_MCS_Instance_2_n31}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U24 ( .a ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, LED_128_Instance_MCS_Instance_2_n14}), .b ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, LED_128_Instance_MCS_Instance_2_n13}), .c ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, LED_128_Instance_MCS_Instance_2_n15}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U23 ( .a ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, LED_128_Instance_MCS_Instance_2_n13}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U22 ( .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, LED_128_Instance_MCS_Instance_2_n12}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, LED_128_Instance_MCS_Instance_2_n14}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U21 ( .a ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, LED_128_Instance_MCS_Instance_2_n11}), .b ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, LED_128_Instance_MCS_Instance_2_n10}), .c ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, LED_128_Instance_mixcolumns_out[24]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U20 ( .a ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, LED_128_Instance_subcells_out[55]}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, LED_128_Instance_MCS_Instance_2_n10}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U19 ( .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, LED_128_Instance_subcells_out[32]}), .b ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, LED_128_Instance_subcells_out[30]}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, LED_128_Instance_MCS_Instance_2_n11}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U18 ( .a ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, LED_128_Instance_MCS_Instance_2_n9}), .b ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, LED_128_Instance_MCS_Instance_2_n8}), .c ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, LED_128_Instance_mixcolumns_out[27]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U17 ( .a ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, LED_128_Instance_MCS_Instance_2_n8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U16 ( .a ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, LED_128_Instance_mixcolumns_out[10]}), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, LED_128_Instance_subcells_out[29]}), .c ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, LED_128_Instance_MCS_Instance_2_n9}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U15 ( .a ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, LED_128_Instance_MCS_Instance_2_n7}), .b ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, LED_128_Instance_MCS_Instance_2_n6}), .c ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, LED_128_Instance_mixcolumns_out[10]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U14 ( .a ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, LED_128_Instance_MCS_Instance_2_n5}), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, LED_128_Instance_subcells_out[11]}), .c ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, LED_128_Instance_MCS_Instance_2_n6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U13 ( .a ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, LED_128_Instance_subcells_out[8]}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, LED_128_Instance_MCS_Instance_2_n7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U12 ( .a ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, LED_128_Instance_MCS_Instance_2_n17}), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, LED_128_Instance_mixcolumns_out[25]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U11 ( .a ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, LED_128_Instance_MCS_Instance_2_n4}), .b ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, LED_128_Instance_MCS_Instance_2_n12}), .c ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, LED_128_Instance_MCS_Instance_2_n35}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U10 ( .a ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, LED_128_Instance_mixcolumns_out[8]}), .c ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, LED_128_Instance_MCS_Instance_2_n12}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U9 ( .a ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, LED_128_Instance_subcells_out[31]}), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, LED_128_Instance_MCS_Instance_2_n5}), .c ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, LED_128_Instance_MCS_Instance_2_n4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U8 ( .a ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, LED_128_Instance_subcells_out[30]}), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, LED_128_Instance_subcells_out[33]}), .c ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, LED_128_Instance_MCS_Instance_2_n5}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U7 ( .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, LED_128_Instance_subcells_out[52]}), .c ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, LED_128_Instance_MCS_Instance_2_n17}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U6 ( .a ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, LED_128_Instance_MCS_Instance_2_n3}), .b ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, LED_128_Instance_MCS_Instance_2_n2}), .c ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, LED_128_Instance_mixcolumns_out[8]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U5 ( .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, LED_128_Instance_MCS_Instance_2_n2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U4 ( .a ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, LED_128_Instance_subcells_out[10]}), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, LED_128_Instance_subcells_out[28]}), .c ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, LED_128_Instance_MCS_Instance_2_n3}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U3 ( .a ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, LED_128_Instance_MCS_Instance_2_n1}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, LED_128_Instance_subcells_out[54]}), .c ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, LED_128_Instance_mixcolumns_out[11]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_2_U2 ( .a ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, LED_128_Instance_MCS_Instance_2_n20}), .b ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, LED_128_Instance_subcells_out[9]}), .c ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, LED_128_Instance_MCS_Instance_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_2_U1 ( .a ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, LED_128_Instance_subcells_out[31]}), .c ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, LED_128_Instance_MCS_Instance_2_n20}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U54 ( .a ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, LED_128_Instance_MCS_Instance_3_n38}), .b ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, LED_128_Instance_MCS_Instance_3_n37}), .c ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, LED_128_Instance_mixcolumns_out[63]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U53 ( .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, LED_128_Instance_MCS_Instance_3_n37}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U52 ( .a ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, LED_128_Instance_mixcolumns_out[46]}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, LED_128_Instance_mixcolumns_out[30]}), .c ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, LED_128_Instance_MCS_Instance_3_n38}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U51 ( .a ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, LED_128_Instance_MCS_Instance_3_n36}), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, LED_128_Instance_mixcolumns_out[46]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U50 ( .a ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, LED_128_Instance_MCS_Instance_3_n34}), .c ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, LED_128_Instance_MCS_Instance_3_n36}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U49 ( .a ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, LED_128_Instance_MCS_Instance_3_n33}), .b ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, LED_128_Instance_mixcolumns_out[45]}), .c ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, LED_128_Instance_mixcolumns_out[62]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U48 ( .a ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, LED_128_Instance_mixcolumns_out[14]}), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, LED_128_Instance_MCS_Instance_3_n33}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U47 ( .a ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, LED_128_Instance_MCS_Instance_3_n32}), .b ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, LED_128_Instance_MCS_Instance_3_n31}), .c ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, LED_128_Instance_mixcolumns_out[61]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U46 ( .a ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, LED_128_Instance_MCS_Instance_3_n30}), .b ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, LED_128_Instance_MCS_Instance_3_n29}), .c ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, LED_128_Instance_MCS_Instance_3_n32}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U45 ( .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, LED_128_Instance_mixcolumns_out[13]}), .c ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, LED_128_Instance_MCS_Instance_3_n29}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U44 ( .a ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, LED_128_Instance_mixcolumns_out[44]}), .b ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, LED_128_Instance_MCS_Instance_3_n28}), .c ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, LED_128_Instance_MCS_Instance_3_n30}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U43 ( .a ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, LED_128_Instance_MCS_Instance_3_n27}), .b ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, LED_128_Instance_MCS_Instance_3_n26}), .c ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, LED_128_Instance_mixcolumns_out[44]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U42 ( .a ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, LED_128_Instance_mixcolumns_out[15]}), .c ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, LED_128_Instance_MCS_Instance_3_n26}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U41 ( .a ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, LED_128_Instance_subcells_out[56]}), .b ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, LED_128_Instance_mixcolumns_out[31]}), .c ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, LED_128_Instance_MCS_Instance_3_n27}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U40 ( .a ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, LED_128_Instance_MCS_Instance_3_n25}), .b ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, LED_128_Instance_mixcolumns_out[12]}), .c ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, LED_128_Instance_mixcolumns_out[60]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U39 ( .a ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, LED_128_Instance_mixcolumns_out[31]}), .b ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, LED_128_Instance_MCS_Instance_3_n28}), .c ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, LED_128_Instance_MCS_Instance_3_n25}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U38 ( .a ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, LED_128_Instance_mixcolumns_out[47]}), .c ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, LED_128_Instance_MCS_Instance_3_n28}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U37 ( .a ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, LED_128_Instance_MCS_Instance_3_n24}), .b ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, LED_128_Instance_MCS_Instance_3_n23}), .c ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, LED_128_Instance_mixcolumns_out[47]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U36 ( .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, LED_128_Instance_subcells_out[37]}), .c ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, LED_128_Instance_MCS_Instance_3_n23}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U35 ( .a ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, LED_128_Instance_mixcolumns_out[30]}), .b ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, LED_128_Instance_mixcolumns_out[14]}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, LED_128_Instance_MCS_Instance_3_n24}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U34 ( .a ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, LED_128_Instance_MCS_Instance_3_n22}), .b ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, LED_128_Instance_MCS_Instance_3_n21}), .c ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, LED_128_Instance_mixcolumns_out[30]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U33 ( .a ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, LED_128_Instance_MCS_Instance_3_n20}), .b ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, LED_128_Instance_MCS_Instance_3_n21}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U32 ( .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, LED_128_Instance_mixcolumns_out[13]}), .b ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, LED_128_Instance_subcells_out[16]}), .c ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, LED_128_Instance_MCS_Instance_3_n22}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U31 ( .a ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, LED_128_Instance_MCS_Instance_3_n19}), .b ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, LED_128_Instance_MCS_Instance_3_n18}), .c ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, LED_128_Instance_mixcolumns_out[13]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U30 ( .a ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, LED_128_Instance_subcells_out[36]}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, LED_128_Instance_MCS_Instance_3_n18}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U29 ( .a ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, LED_128_Instance_MCS_Instance_3_n17}), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, LED_128_Instance_MCS_Instance_3_n34}), .c ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, LED_128_Instance_MCS_Instance_3_n19}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U28 ( .a ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, LED_128_Instance_MCS_Instance_3_n16}), .b ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, LED_128_Instance_subcells_out[14]}), .c ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, LED_128_Instance_MCS_Instance_3_n34}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U27 ( .a ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, LED_128_Instance_subcells_out[17]}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, LED_128_Instance_subcells_out[15]}), .c ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, LED_128_Instance_MCS_Instance_3_n16}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U26 ( .a ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, LED_128_Instance_MCS_Instance_3_n15}), .b ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, LED_128_Instance_MCS_Instance_3_n31}), .c ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, LED_128_Instance_mixcolumns_out[45]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U25 ( .a ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, LED_128_Instance_mixcolumns_out[28]}), .b ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, LED_128_Instance_mixcolumns_out[31]}), .c ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, LED_128_Instance_MCS_Instance_3_n31}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U24 ( .a ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, LED_128_Instance_MCS_Instance_3_n14}), .b ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, LED_128_Instance_MCS_Instance_3_n13}), .c ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, LED_128_Instance_MCS_Instance_3_n15}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U23 ( .a ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, LED_128_Instance_MCS_Instance_3_n13}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U22 ( .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, LED_128_Instance_MCS_Instance_3_n12}), .b ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, LED_128_Instance_MCS_Instance_3_n14}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U21 ( .a ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, LED_128_Instance_MCS_Instance_3_n11}), .b ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, LED_128_Instance_MCS_Instance_3_n10}), .c ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, LED_128_Instance_mixcolumns_out[28]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U20 ( .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, LED_128_Instance_subcells_out[59]}), .c ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, LED_128_Instance_MCS_Instance_3_n10}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U19 ( .a ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, LED_128_Instance_subcells_out[36]}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, LED_128_Instance_subcells_out[18]}), .c ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, LED_128_Instance_MCS_Instance_3_n11}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U18 ( .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, LED_128_Instance_MCS_Instance_3_n9}), .b ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, LED_128_Instance_MCS_Instance_3_n8}), .c ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, LED_128_Instance_mixcolumns_out[31]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U17 ( .a ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, LED_128_Instance_MCS_Instance_3_n8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U16 ( .a ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, LED_128_Instance_mixcolumns_out[14]}), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, LED_128_Instance_subcells_out[17]}), .c ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, LED_128_Instance_MCS_Instance_3_n9}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U15 ( .a ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, LED_128_Instance_MCS_Instance_3_n7}), .b ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, LED_128_Instance_MCS_Instance_3_n6}), .c ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, LED_128_Instance_mixcolumns_out[14]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U14 ( .a ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, LED_128_Instance_MCS_Instance_3_n5}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, LED_128_Instance_subcells_out[15]}), .c ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, LED_128_Instance_MCS_Instance_3_n6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U13 ( .a ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, LED_128_Instance_subcells_out[12]}), .b ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, LED_128_Instance_MCS_Instance_3_n7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U12 ( .a ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, LED_128_Instance_MCS_Instance_3_n17}), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, LED_128_Instance_mixcolumns_out[29]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U11 ( .a ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, LED_128_Instance_MCS_Instance_3_n4}), .b ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, LED_128_Instance_MCS_Instance_3_n12}), .c ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, LED_128_Instance_MCS_Instance_3_n35}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U10 ( .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, LED_128_Instance_mixcolumns_out[12]}), .c ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, LED_128_Instance_MCS_Instance_3_n12}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U9 ( .a ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, LED_128_Instance_subcells_out[19]}), .b ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, LED_128_Instance_MCS_Instance_3_n5}), .c ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, LED_128_Instance_MCS_Instance_3_n4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U8 ( .a ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, LED_128_Instance_subcells_out[18]}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, LED_128_Instance_subcells_out[37]}), .c ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, LED_128_Instance_MCS_Instance_3_n5}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U7 ( .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, LED_128_Instance_subcells_out[56]}), .c ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, LED_128_Instance_MCS_Instance_3_n17}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U6 ( .a ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, LED_128_Instance_MCS_Instance_3_n3}), .b ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, LED_128_Instance_MCS_Instance_3_n2}), .c ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, LED_128_Instance_mixcolumns_out[12]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U5 ( .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, LED_128_Instance_MCS_Instance_3_n2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U4 ( .a ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, LED_128_Instance_subcells_out[14]}), .b ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, LED_128_Instance_subcells_out[16]}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, LED_128_Instance_MCS_Instance_3_n3}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U3 ( .a ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, LED_128_Instance_MCS_Instance_3_n1}), .b ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, LED_128_Instance_subcells_out[58]}), .c ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, LED_128_Instance_mixcolumns_out[15]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) LED_128_Instance_MCS_Instance_3_U2 ( .a ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, LED_128_Instance_MCS_Instance_3_n20}), .b ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, LED_128_Instance_subcells_out[13]}), .c ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, LED_128_Instance_MCS_Instance_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) LED_128_Instance_MCS_Instance_3_U1 ( .a ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, LED_128_Instance_subcells_out[19]}), .c ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, LED_128_Instance_MCS_Instance_3_n20}) ) ;
    INV_X1 LED_128_Instance_ks_reg_0__U1 ( .A (LED_128_Instance_ks_reg_0__Q), .ZN (LED_128_Instance_n4) ) ;
    INV_X1 LED_128_Instance_ks_reg_1__U1 ( .A (LED_128_Instance_n26), .ZN (LED_128_Instance_n8) ) ;
    INV_X1 LED_128_Instance_ks_reg_2__U1 ( .A (LED_128_Instance_n25), .ZN (LED_128_Instance_n1) ) ;
    INV_X1 LED_128_Instance_ks_reg_3__U1 ( .A (LED_128_Instance_n2), .ZN (LED_128_Instance_n24) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_0__U1 ( .A (roundconstant[0]), .ZN (LED_128_Instance_n6) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_1__U1 ( .A (roundconstant[1]), .ZN (LED_128_Instance_n29) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_2__U1 ( .A (roundconstant[2]), .ZN (LED_128_Instance_n5) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_3__U1 ( .A (roundconstant[3]), .ZN (LED_128_Instance_n30) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_4__U1 ( .A (roundconstant[4]), .ZN (LED_128_Instance_n28) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_5__U1 ( .A (roundconstant[5]), .ZN (LED_128_Instance_n27) ) ;
    Precharger_reg new_AGEMA_gate_1128 ( .D (LED_128_Instance_n12), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_1333, new_AGEMA_signal_1332}) ) ;
    Precharger_reg new_AGEMA_gate_1129 ( .D (LED_128_Instance_MUX_current_roundkey_n9), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_1465, new_AGEMA_signal_1464}) ) ;
    Precharger_reg new_AGEMA_gate_1130 ( .D (LED_128_Instance_MUX_current_roundkey_n8), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_1551, new_AGEMA_signal_1550}) ) ;
    Precharger_reg new_AGEMA_gate_1131 ( .D (LED_128_Instance_MUX_current_roundkey_n7), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_1559, new_AGEMA_signal_1558}) ) ;
    Precharger_reg new_AGEMA_gate_1132 ( .D (LED_128_Instance_n31), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_1777, new_AGEMA_signal_1776}) ) ;
    Precharger_reg new_AGEMA_gate_1133 ( .D (LED_128_Instance_MUX_addroundkey_out_n7), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_1997, new_AGEMA_signal_1996}) ) ;
    Precharger_reg new_AGEMA_gate_1134 ( .D (LED_128_Instance_MUX_addroundkey_out_n8), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_2025, new_AGEMA_signal_2024}) ) ;
    Precharger_reg new_AGEMA_gate_1135 ( .D (LED_128_Instance_MUX_state0_n9), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_3033, new_AGEMA_signal_3032}) ) ;
    Precharger_reg new_AGEMA_gate_1136 ( .D (LED_128_Instance_MUX_state0_n8), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_3075, new_AGEMA_signal_3074}) ) ;
    Precharger_reg new_AGEMA_gate_1137 ( .D (LED_128_Instance_MUX_state0_n10), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_3079, new_AGEMA_signal_3078}) ) ;
    Precharger_reg new_AGEMA_gate_1138 ( .D (IN_reset), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_3097, new_AGEMA_signal_3096}) ) ;
    Precharger_reg new_AGEMA_gate_1139 ( .D (LED_128_Instance_n22), .mid_rst (mid_rst), .clk (CLK), .Q ({new_AGEMA_signal_3491, new_AGEMA_signal_3490}) ) ;
    ClockController_LMDPL ClockControllerInst ( .clk (CLK), .Po_rst (Po_rst), .pre1 (LMDPL_pre1), .pre2 (LMDPL_pre2), .mid_rst (mid_rst) ) ;
    Precharger PrechargeCell_0 ( .D (IN_plaintext_s1[63]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3649, new_AGEMA_signal_3648}) ) ;
    Precharger PrechargeCell_1 ( .D (IN_plaintext_s1[62]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3645, new_AGEMA_signal_3644}) ) ;
    Precharger PrechargeCell_2 ( .D (IN_plaintext_s1[61]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3721, new_AGEMA_signal_3720}) ) ;
    Precharger PrechargeCell_3 ( .D (IN_plaintext_s1[60]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3697, new_AGEMA_signal_3696}) ) ;
    Precharger PrechargeCell_4 ( .D (IN_plaintext_s1[59]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3609, new_AGEMA_signal_3608}) ) ;
    Precharger PrechargeCell_5 ( .D (IN_plaintext_s1[58]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3605, new_AGEMA_signal_3604}) ) ;
    Precharger PrechargeCell_6 ( .D (IN_plaintext_s1[57]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3717, new_AGEMA_signal_3716}) ) ;
    Precharger PrechargeCell_7 ( .D (IN_plaintext_s1[56]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3693, new_AGEMA_signal_3692}) ) ;
    Precharger PrechargeCell_8 ( .D (IN_plaintext_s1[55]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3641, new_AGEMA_signal_3640}) ) ;
    Precharger PrechargeCell_9 ( .D (IN_plaintext_s1[54]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3601, new_AGEMA_signal_3600}) ) ;
    Precharger PrechargeCell_10 ( .D (IN_plaintext_s1[53]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3729, new_AGEMA_signal_3728}) ) ;
    Precharger PrechargeCell_11 ( .D (IN_plaintext_s1[52]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3713, new_AGEMA_signal_3712}) ) ;
    Precharger PrechargeCell_12 ( .D (IN_plaintext_s1[51]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3637, new_AGEMA_signal_3636}) ) ;
    Precharger PrechargeCell_13 ( .D (IN_plaintext_s1[50]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3633, new_AGEMA_signal_3632}) ) ;
    Precharger PrechargeCell_14 ( .D (IN_plaintext_s1[49]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3725, new_AGEMA_signal_3724}) ) ;
    Precharger PrechargeCell_15 ( .D (IN_plaintext_s1[48]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3709, new_AGEMA_signal_3708}) ) ;
    Precharger PrechargeCell_16 ( .D (IN_plaintext_s1[47]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3597, new_AGEMA_signal_3596}) ) ;
    Precharger PrechargeCell_17 ( .D (IN_plaintext_s1[46]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3549, new_AGEMA_signal_3548}) ) ;
    Precharger PrechargeCell_18 ( .D (IN_plaintext_s1[45]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3593, new_AGEMA_signal_3592}) ) ;
    Precharger PrechargeCell_19 ( .D (IN_plaintext_s1[44]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3545, new_AGEMA_signal_3544}) ) ;
    Precharger PrechargeCell_20 ( .D (IN_plaintext_s1[43]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3589, new_AGEMA_signal_3588}) ) ;
    Precharger PrechargeCell_21 ( .D (IN_plaintext_s1[42]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3461, new_AGEMA_signal_3460}) ) ;
    Precharger PrechargeCell_22 ( .D (IN_plaintext_s1[41]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3541, new_AGEMA_signal_3540}) ) ;
    Precharger PrechargeCell_23 ( .D (IN_plaintext_s1[40]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3537, new_AGEMA_signal_3536}) ) ;
    Precharger PrechargeCell_24 ( .D (IN_plaintext_s1[39]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3629, new_AGEMA_signal_3628}) ) ;
    Precharger PrechargeCell_25 ( .D (IN_plaintext_s1[38]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3457, new_AGEMA_signal_3456}) ) ;
    Precharger PrechargeCell_26 ( .D (IN_plaintext_s1[37]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3533, new_AGEMA_signal_3532}) ) ;
    Precharger PrechargeCell_27 ( .D (IN_plaintext_s1[36]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3529, new_AGEMA_signal_3528}) ) ;
    Precharger PrechargeCell_28 ( .D (IN_plaintext_s1[35]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3625, new_AGEMA_signal_3624}) ) ;
    Precharger PrechargeCell_29 ( .D (IN_plaintext_s1[34]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3525, new_AGEMA_signal_3524}) ) ;
    Precharger PrechargeCell_30 ( .D (IN_plaintext_s1[33]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3585, new_AGEMA_signal_3584}) ) ;
    Precharger PrechargeCell_31 ( .D (IN_plaintext_s1[32]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3521, new_AGEMA_signal_3520}) ) ;
    Precharger PrechargeCell_32 ( .D (IN_plaintext_s1[31]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3363, new_AGEMA_signal_3362}) ) ;
    Precharger PrechargeCell_33 ( .D (IN_plaintext_s1[30]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3453, new_AGEMA_signal_3452}) ) ;
    Precharger PrechargeCell_34 ( .D (IN_plaintext_s1[29]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3517, new_AGEMA_signal_3516}) ) ;
    Precharger PrechargeCell_35 ( .D (IN_plaintext_s1[28]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3449, new_AGEMA_signal_3448}) ) ;
    Precharger PrechargeCell_36 ( .D (IN_plaintext_s1[27]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3359, new_AGEMA_signal_3358}) ) ;
    Precharger PrechargeCell_37 ( .D (IN_plaintext_s1[26]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3445, new_AGEMA_signal_3444}) ) ;
    Precharger PrechargeCell_38 ( .D (IN_plaintext_s1[25]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3441, new_AGEMA_signal_3440}) ) ;
    Precharger PrechargeCell_39 ( .D (IN_plaintext_s1[24]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3355, new_AGEMA_signal_3354}) ) ;
    Precharger PrechargeCell_40 ( .D (IN_plaintext_s1[23]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3351, new_AGEMA_signal_3350}) ) ;
    Precharger PrechargeCell_41 ( .D (IN_plaintext_s1[22]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3513, new_AGEMA_signal_3512}) ) ;
    Precharger PrechargeCell_42 ( .D (IN_plaintext_s1[21]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3437, new_AGEMA_signal_3436}) ) ;
    Precharger PrechargeCell_43 ( .D (IN_plaintext_s1[20]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3347, new_AGEMA_signal_3346}) ) ;
    Precharger PrechargeCell_44 ( .D (IN_plaintext_s1[19]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3343, new_AGEMA_signal_3342}) ) ;
    Precharger PrechargeCell_45 ( .D (IN_plaintext_s1[18]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3509, new_AGEMA_signal_3508}) ) ;
    Precharger PrechargeCell_46 ( .D (IN_plaintext_s1[17]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3505, new_AGEMA_signal_3504}) ) ;
    Precharger PrechargeCell_47 ( .D (IN_plaintext_s1[16]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3433, new_AGEMA_signal_3432}) ) ;
    Precharger PrechargeCell_48 ( .D (IN_plaintext_s1[15]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3263, new_AGEMA_signal_3262}) ) ;
    Precharger PrechargeCell_49 ( .D (IN_plaintext_s1[14]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3183, new_AGEMA_signal_3182}) ) ;
    Precharger PrechargeCell_50 ( .D (IN_plaintext_s1[13]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3259, new_AGEMA_signal_3258}) ) ;
    Precharger PrechargeCell_51 ( .D (IN_plaintext_s1[12]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3179, new_AGEMA_signal_3178}) ) ;
    Precharger PrechargeCell_52 ( .D (IN_plaintext_s1[11]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3175, new_AGEMA_signal_3174}) ) ;
    Precharger PrechargeCell_53 ( .D (IN_plaintext_s1[10]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3171, new_AGEMA_signal_3170}) ) ;
    Precharger PrechargeCell_54 ( .D (IN_plaintext_s1[9]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3255, new_AGEMA_signal_3254}) ) ;
    Precharger PrechargeCell_55 ( .D (IN_plaintext_s1[8]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3167, new_AGEMA_signal_3166}) ) ;
    Precharger PrechargeCell_56 ( .D (IN_plaintext_s1[7]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3163, new_AGEMA_signal_3162}) ) ;
    Precharger PrechargeCell_57 ( .D (IN_plaintext_s1[6]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3159, new_AGEMA_signal_3158}) ) ;
    Precharger PrechargeCell_58 ( .D (IN_plaintext_s1[5]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3339, new_AGEMA_signal_3338}) ) ;
    Precharger PrechargeCell_59 ( .D (IN_plaintext_s1[4]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3155, new_AGEMA_signal_3154}) ) ;
    Precharger PrechargeCell_60 ( .D (IN_plaintext_s1[3]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3251, new_AGEMA_signal_3250}) ) ;
    Precharger PrechargeCell_61 ( .D (IN_plaintext_s1[2]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3151, new_AGEMA_signal_3150}) ) ;
    Precharger PrechargeCell_62 ( .D (IN_plaintext_s1[1]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3335, new_AGEMA_signal_3334}) ) ;
    Precharger PrechargeCell_63 ( .D (IN_plaintext_s1[0]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3099, new_AGEMA_signal_3098}) ) ;
    Precharger PrechargeCell_64 ( .D (IN_key_s1[127]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1771, new_AGEMA_signal_1770}) ) ;
    Precharger PrechargeCell_65 ( .D (IN_key_s1[126]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1765, new_AGEMA_signal_1764}) ) ;
    Precharger PrechargeCell_66 ( .D (IN_key_s1[125]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1759, new_AGEMA_signal_1758}) ) ;
    Precharger PrechargeCell_67 ( .D (IN_key_s1[124]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1753, new_AGEMA_signal_1752}) ) ;
    Precharger PrechargeCell_68 ( .D (IN_key_s1[123]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1747, new_AGEMA_signal_1746}) ) ;
    Precharger PrechargeCell_69 ( .D (IN_key_s1[122]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1741, new_AGEMA_signal_1740}) ) ;
    Precharger PrechargeCell_70 ( .D (IN_key_s1[121]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1735, new_AGEMA_signal_1734}) ) ;
    Precharger PrechargeCell_71 ( .D (IN_key_s1[120]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1729, new_AGEMA_signal_1728}) ) ;
    Precharger PrechargeCell_72 ( .D (IN_key_s1[119]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1723, new_AGEMA_signal_1722}) ) ;
    Precharger PrechargeCell_73 ( .D (IN_key_s1[118]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1717, new_AGEMA_signal_1716}) ) ;
    Precharger PrechargeCell_74 ( .D (IN_key_s1[117]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1711, new_AGEMA_signal_1710}) ) ;
    Precharger PrechargeCell_75 ( .D (IN_key_s1[116]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1705, new_AGEMA_signal_1704}) ) ;
    Precharger PrechargeCell_76 ( .D (IN_key_s1[115]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1699, new_AGEMA_signal_1698}) ) ;
    Precharger PrechargeCell_77 ( .D (IN_key_s1[114]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1693, new_AGEMA_signal_1692}) ) ;
    Precharger PrechargeCell_78 ( .D (IN_key_s1[113]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1687, new_AGEMA_signal_1686}) ) ;
    Precharger PrechargeCell_79 ( .D (IN_key_s1[112]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1681, new_AGEMA_signal_1680}) ) ;
    Precharger PrechargeCell_80 ( .D (IN_key_s1[111]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1675, new_AGEMA_signal_1674}) ) ;
    Precharger PrechargeCell_81 ( .D (IN_key_s1[110]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1669, new_AGEMA_signal_1668}) ) ;
    Precharger PrechargeCell_82 ( .D (IN_key_s1[109]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1663, new_AGEMA_signal_1662}) ) ;
    Precharger PrechargeCell_83 ( .D (IN_key_s1[108]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1657, new_AGEMA_signal_1656}) ) ;
    Precharger PrechargeCell_84 ( .D (IN_key_s1[107]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1651, new_AGEMA_signal_1650}) ) ;
    Precharger PrechargeCell_85 ( .D (IN_key_s1[106]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1645, new_AGEMA_signal_1644}) ) ;
    Precharger PrechargeCell_86 ( .D (IN_key_s1[105]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1639, new_AGEMA_signal_1638}) ) ;
    Precharger PrechargeCell_87 ( .D (IN_key_s1[104]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1633, new_AGEMA_signal_1632}) ) ;
    Precharger PrechargeCell_88 ( .D (IN_key_s1[103]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1407, new_AGEMA_signal_1406}) ) ;
    Precharger PrechargeCell_89 ( .D (IN_key_s1[102]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1627, new_AGEMA_signal_1626}) ) ;
    Precharger PrechargeCell_90 ( .D (IN_key_s1[101]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1621, new_AGEMA_signal_1620}) ) ;
    Precharger PrechargeCell_91 ( .D (IN_key_s1[100]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1401, new_AGEMA_signal_1400}) ) ;
    Precharger PrechargeCell_92 ( .D (IN_key_s1[99]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1395, new_AGEMA_signal_1394}) ) ;
    Precharger PrechargeCell_93 ( .D (IN_key_s1[98]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1389, new_AGEMA_signal_1388}) ) ;
    Precharger PrechargeCell_94 ( .D (IN_key_s1[97]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1615, new_AGEMA_signal_1614}) ) ;
    Precharger PrechargeCell_95 ( .D (IN_key_s1[96]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1383, new_AGEMA_signal_1382}) ) ;
    Precharger PrechargeCell_96 ( .D (IN_key_s1[95]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1609, new_AGEMA_signal_1608}) ) ;
    Precharger PrechargeCell_97 ( .D (IN_key_s1[94]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1603, new_AGEMA_signal_1602}) ) ;
    Precharger PrechargeCell_98 ( .D (IN_key_s1[93]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1597, new_AGEMA_signal_1596}) ) ;
    Precharger PrechargeCell_99 ( .D (IN_key_s1[92]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1377, new_AGEMA_signal_1376}) ) ;
    Precharger PrechargeCell_100 ( .D (IN_key_s1[91]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1591, new_AGEMA_signal_1590}) ) ;
    Precharger PrechargeCell_101 ( .D (IN_key_s1[90]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1371, new_AGEMA_signal_1370}) ) ;
    Precharger PrechargeCell_102 ( .D (IN_key_s1[89]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1585, new_AGEMA_signal_1584}) ) ;
    Precharger PrechargeCell_103 ( .D (IN_key_s1[88]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1365, new_AGEMA_signal_1364}) ) ;
    Precharger PrechargeCell_104 ( .D (IN_key_s1[87]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1579, new_AGEMA_signal_1578}) ) ;
    Precharger PrechargeCell_105 ( .D (IN_key_s1[86]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1359, new_AGEMA_signal_1358}) ) ;
    Precharger PrechargeCell_106 ( .D (IN_key_s1[85]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1573, new_AGEMA_signal_1572}) ) ;
    Precharger PrechargeCell_107 ( .D (IN_key_s1[84]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1567, new_AGEMA_signal_1566}) ) ;
    Precharger PrechargeCell_108 ( .D (IN_key_s1[83]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1353, new_AGEMA_signal_1352}) ) ;
    Precharger PrechargeCell_109 ( .D (IN_key_s1[82]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1561, new_AGEMA_signal_1560}) ) ;
    Precharger PrechargeCell_110 ( .D (IN_key_s1[81]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1553, new_AGEMA_signal_1552}) ) ;
    Precharger PrechargeCell_111 ( .D (IN_key_s1[80]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1347, new_AGEMA_signal_1346}) ) ;
    Precharger PrechargeCell_112 ( .D (IN_key_s1[79]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1545, new_AGEMA_signal_1544}) ) ;
    Precharger PrechargeCell_113 ( .D (IN_key_s1[78]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1539, new_AGEMA_signal_1538}) ) ;
    Precharger PrechargeCell_114 ( .D (IN_key_s1[77]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1533, new_AGEMA_signal_1532}) ) ;
    Precharger PrechargeCell_115 ( .D (IN_key_s1[76]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1527, new_AGEMA_signal_1526}) ) ;
    Precharger PrechargeCell_116 ( .D (IN_key_s1[75]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1521, new_AGEMA_signal_1520}) ) ;
    Precharger PrechargeCell_117 ( .D (IN_key_s1[74]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1515, new_AGEMA_signal_1514}) ) ;
    Precharger PrechargeCell_118 ( .D (IN_key_s1[73]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1509, new_AGEMA_signal_1508}) ) ;
    Precharger PrechargeCell_119 ( .D (IN_key_s1[72]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1503, new_AGEMA_signal_1502}) ) ;
    Precharger PrechargeCell_120 ( .D (IN_key_s1[71]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1497, new_AGEMA_signal_1496}) ) ;
    Precharger PrechargeCell_121 ( .D (IN_key_s1[70]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1491, new_AGEMA_signal_1490}) ) ;
    Precharger PrechargeCell_122 ( .D (IN_key_s1[69]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1485, new_AGEMA_signal_1484}) ) ;
    Precharger PrechargeCell_123 ( .D (IN_key_s1[68]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1479, new_AGEMA_signal_1478}) ) ;
    Precharger PrechargeCell_124 ( .D (IN_key_s1[67]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1341, new_AGEMA_signal_1340}) ) ;
    Precharger PrechargeCell_125 ( .D (IN_key_s1[66]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1473, new_AGEMA_signal_1472}) ) ;
    Precharger PrechargeCell_126 ( .D (IN_key_s1[65]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1467, new_AGEMA_signal_1466}) ) ;
    Precharger PrechargeCell_127 ( .D (IN_key_s1[64]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1335, new_AGEMA_signal_1334}) ) ;
    Precharger PrechargeCell_128 ( .D (IN_key_s1[63]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1773, new_AGEMA_signal_1772}) ) ;
    Precharger PrechargeCell_129 ( .D (IN_key_s1[62]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1767, new_AGEMA_signal_1766}) ) ;
    Precharger PrechargeCell_130 ( .D (IN_key_s1[61]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1761, new_AGEMA_signal_1760}) ) ;
    Precharger PrechargeCell_131 ( .D (IN_key_s1[60]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1755, new_AGEMA_signal_1754}) ) ;
    Precharger PrechargeCell_132 ( .D (IN_key_s1[59]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1749, new_AGEMA_signal_1748}) ) ;
    Precharger PrechargeCell_133 ( .D (IN_key_s1[58]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1743, new_AGEMA_signal_1742}) ) ;
    Precharger PrechargeCell_134 ( .D (IN_key_s1[57]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1737, new_AGEMA_signal_1736}) ) ;
    Precharger PrechargeCell_135 ( .D (IN_key_s1[56]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1731, new_AGEMA_signal_1730}) ) ;
    Precharger PrechargeCell_136 ( .D (IN_key_s1[55]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1725, new_AGEMA_signal_1724}) ) ;
    Precharger PrechargeCell_137 ( .D (IN_key_s1[54]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1719, new_AGEMA_signal_1718}) ) ;
    Precharger PrechargeCell_138 ( .D (IN_key_s1[53]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1713, new_AGEMA_signal_1712}) ) ;
    Precharger PrechargeCell_139 ( .D (IN_key_s1[52]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1707, new_AGEMA_signal_1706}) ) ;
    Precharger PrechargeCell_140 ( .D (IN_key_s1[51]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1701, new_AGEMA_signal_1700}) ) ;
    Precharger PrechargeCell_141 ( .D (IN_key_s1[50]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1695, new_AGEMA_signal_1694}) ) ;
    Precharger PrechargeCell_142 ( .D (IN_key_s1[49]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1689, new_AGEMA_signal_1688}) ) ;
    Precharger PrechargeCell_143 ( .D (IN_key_s1[48]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1683, new_AGEMA_signal_1682}) ) ;
    Precharger PrechargeCell_144 ( .D (IN_key_s1[47]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1677, new_AGEMA_signal_1676}) ) ;
    Precharger PrechargeCell_145 ( .D (IN_key_s1[46]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1671, new_AGEMA_signal_1670}) ) ;
    Precharger PrechargeCell_146 ( .D (IN_key_s1[45]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1665, new_AGEMA_signal_1664}) ) ;
    Precharger PrechargeCell_147 ( .D (IN_key_s1[44]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1659, new_AGEMA_signal_1658}) ) ;
    Precharger PrechargeCell_148 ( .D (IN_key_s1[43]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1653, new_AGEMA_signal_1652}) ) ;
    Precharger PrechargeCell_149 ( .D (IN_key_s1[42]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1647, new_AGEMA_signal_1646}) ) ;
    Precharger PrechargeCell_150 ( .D (IN_key_s1[41]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1641, new_AGEMA_signal_1640}) ) ;
    Precharger PrechargeCell_151 ( .D (IN_key_s1[40]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1635, new_AGEMA_signal_1634}) ) ;
    Precharger PrechargeCell_152 ( .D (IN_key_s1[39]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1409, new_AGEMA_signal_1408}) ) ;
    Precharger PrechargeCell_153 ( .D (IN_key_s1[38]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1629, new_AGEMA_signal_1628}) ) ;
    Precharger PrechargeCell_154 ( .D (IN_key_s1[37]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1623, new_AGEMA_signal_1622}) ) ;
    Precharger PrechargeCell_155 ( .D (IN_key_s1[36]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1403, new_AGEMA_signal_1402}) ) ;
    Precharger PrechargeCell_156 ( .D (IN_key_s1[35]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1397, new_AGEMA_signal_1396}) ) ;
    Precharger PrechargeCell_157 ( .D (IN_key_s1[34]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1391, new_AGEMA_signal_1390}) ) ;
    Precharger PrechargeCell_158 ( .D (IN_key_s1[33]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1617, new_AGEMA_signal_1616}) ) ;
    Precharger PrechargeCell_159 ( .D (IN_key_s1[32]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1385, new_AGEMA_signal_1384}) ) ;
    Precharger PrechargeCell_160 ( .D (IN_key_s1[31]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1611, new_AGEMA_signal_1610}) ) ;
    Precharger PrechargeCell_161 ( .D (IN_key_s1[30]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1605, new_AGEMA_signal_1604}) ) ;
    Precharger PrechargeCell_162 ( .D (IN_key_s1[29]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1599, new_AGEMA_signal_1598}) ) ;
    Precharger PrechargeCell_163 ( .D (IN_key_s1[28]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1379, new_AGEMA_signal_1378}) ) ;
    Precharger PrechargeCell_164 ( .D (IN_key_s1[27]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1593, new_AGEMA_signal_1592}) ) ;
    Precharger PrechargeCell_165 ( .D (IN_key_s1[26]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1373, new_AGEMA_signal_1372}) ) ;
    Precharger PrechargeCell_166 ( .D (IN_key_s1[25]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1587, new_AGEMA_signal_1586}) ) ;
    Precharger PrechargeCell_167 ( .D (IN_key_s1[24]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1367, new_AGEMA_signal_1366}) ) ;
    Precharger PrechargeCell_168 ( .D (IN_key_s1[23]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1581, new_AGEMA_signal_1580}) ) ;
    Precharger PrechargeCell_169 ( .D (IN_key_s1[22]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1361, new_AGEMA_signal_1360}) ) ;
    Precharger PrechargeCell_170 ( .D (IN_key_s1[21]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1575, new_AGEMA_signal_1574}) ) ;
    Precharger PrechargeCell_171 ( .D (IN_key_s1[20]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1569, new_AGEMA_signal_1568}) ) ;
    Precharger PrechargeCell_172 ( .D (IN_key_s1[19]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1355, new_AGEMA_signal_1354}) ) ;
    Precharger PrechargeCell_173 ( .D (IN_key_s1[18]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1563, new_AGEMA_signal_1562}) ) ;
    Precharger PrechargeCell_174 ( .D (IN_key_s1[17]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1555, new_AGEMA_signal_1554}) ) ;
    Precharger PrechargeCell_175 ( .D (IN_key_s1[16]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1349, new_AGEMA_signal_1348}) ) ;
    Precharger PrechargeCell_176 ( .D (IN_key_s1[15]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1547, new_AGEMA_signal_1546}) ) ;
    Precharger PrechargeCell_177 ( .D (IN_key_s1[14]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1541, new_AGEMA_signal_1540}) ) ;
    Precharger PrechargeCell_178 ( .D (IN_key_s1[13]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1535, new_AGEMA_signal_1534}) ) ;
    Precharger PrechargeCell_179 ( .D (IN_key_s1[12]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1529, new_AGEMA_signal_1528}) ) ;
    Precharger PrechargeCell_180 ( .D (IN_key_s1[11]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1523, new_AGEMA_signal_1522}) ) ;
    Precharger PrechargeCell_181 ( .D (IN_key_s1[10]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1517, new_AGEMA_signal_1516}) ) ;
    Precharger PrechargeCell_182 ( .D (IN_key_s1[9]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1511, new_AGEMA_signal_1510}) ) ;
    Precharger PrechargeCell_183 ( .D (IN_key_s1[8]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1505, new_AGEMA_signal_1504}) ) ;
    Precharger PrechargeCell_184 ( .D (IN_key_s1[7]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1499, new_AGEMA_signal_1498}) ) ;
    Precharger PrechargeCell_185 ( .D (IN_key_s1[6]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1493, new_AGEMA_signal_1492}) ) ;
    Precharger PrechargeCell_186 ( .D (IN_key_s1[5]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1487, new_AGEMA_signal_1486}) ) ;
    Precharger PrechargeCell_187 ( .D (IN_key_s1[4]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1481, new_AGEMA_signal_1480}) ) ;
    Precharger PrechargeCell_188 ( .D (IN_key_s1[3]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1343, new_AGEMA_signal_1342}) ) ;
    Precharger PrechargeCell_189 ( .D (IN_key_s1[2]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1475, new_AGEMA_signal_1474}) ) ;
    Precharger PrechargeCell_190 ( .D (IN_key_s1[1]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1469, new_AGEMA_signal_1468}) ) ;
    Precharger PrechargeCell_191 ( .D (IN_key_s1[0]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1337, new_AGEMA_signal_1336}) ) ;

    /* register cells */
    reg_sr_LMDPL LED_128_Instance_ks_reg_0__FF_FF ( .D (LED_128_Instance_N10), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (LED_128_Instance_ks_reg_0__Q), .QN () ) ;
    reg_sr_LMDPL LED_128_Instance_ks_reg_1__FF_FF ( .D (LED_128_Instance_N11), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (LED_128_Instance_n26), .QN () ) ;
    reg_sr_LMDPL LED_128_Instance_ks_reg_2__FF_FF ( .D (LED_128_Instance_N12), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (LED_128_Instance_n25), .QN () ) ;
    reg_sr_LMDPL LED_128_Instance_ks_reg_3__FF_FF ( .D (LED_128_Instance_N13), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (LED_128_Instance_n2), .QN () ) ;
    reg_sr_LMDPL LED_128_Instance_roundconstant_reg_0__FF_FF ( .D (LED_128_Instance_N4), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (roundconstant[0]), .QN () ) ;
    reg_sr_LMDPL LED_128_Instance_roundconstant_reg_1__FF_FF ( .D (LED_128_Instance_N5), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (roundconstant[1]), .QN () ) ;
    reg_sr_LMDPL LED_128_Instance_roundconstant_reg_2__FF_FF ( .D (LED_128_Instance_N6), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (roundconstant[2]), .QN () ) ;
    reg_sr_LMDPL LED_128_Instance_roundconstant_reg_3__FF_FF ( .D (LED_128_Instance_N7), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (roundconstant[3]), .QN () ) ;
    reg_sr_LMDPL LED_128_Instance_roundconstant_reg_4__FF_FF ( .D (LED_128_Instance_N8), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (roundconstant[4]), .QN () ) ;
    reg_sr_LMDPL LED_128_Instance_roundconstant_reg_5__FF_FF ( .D (LED_128_Instance_N9), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (roundconstant[5]), .QN () ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_0__FF_FF ( .D ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, LED_128_Instance_state1[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1461, OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_1__FF_FF ( .D ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, LED_128_Instance_state1[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1961, OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_2__FF_FF ( .D ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, LED_128_Instance_state1[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1933, OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_3__FF_FF ( .D ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, LED_128_Instance_state1[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1413, OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_4__FF_FF ( .D ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, LED_128_Instance_state1[4]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1869, OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_5__FF_FF ( .D ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, LED_128_Instance_state1[5]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1825, OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_6__FF_FF ( .D ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, LED_128_Instance_state1[6]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1805, OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_7__FF_FF ( .D ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, LED_128_Instance_state1[7]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1801, OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_8__FF_FF ( .D ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, LED_128_Instance_state1[8]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1797, OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_9__FF_FF ( .D ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, LED_128_Instance_state1[9]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1793, OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_10__FF_FF ( .D ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, LED_128_Instance_state1[10]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1993, OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_11__FF_FF ( .D ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, LED_128_Instance_state1[11]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1989, OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_12__FF_FF ( .D ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, LED_128_Instance_state1[12]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1985, OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_13__FF_FF ( .D ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, LED_128_Instance_state1[13]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1981, OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_14__FF_FF ( .D ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, LED_128_Instance_state1[14]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1977, OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_15__FF_FF ( .D ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, LED_128_Instance_state1[15]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1973, OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_16__FF_FF ( .D ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, LED_128_Instance_state1[16]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1457, OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_17__FF_FF ( .D ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, LED_128_Instance_state1[17]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1969, OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_18__FF_FF ( .D ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, LED_128_Instance_state1[18]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1965, OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_19__FF_FF ( .D ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, LED_128_Instance_state1[19]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1453, OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_20__FF_FF ( .D ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, LED_128_Instance_state1[20]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1957, OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_21__FF_FF ( .D ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, LED_128_Instance_state1[21]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1953, OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_22__FF_FF ( .D ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, LED_128_Instance_state1[22]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1449, OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_23__FF_FF ( .D ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, LED_128_Instance_state1[23]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1949, OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_24__FF_FF ( .D ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, LED_128_Instance_state1[24]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1445, OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_25__FF_FF ( .D ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, LED_128_Instance_state1[25]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1945, OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_26__FF_FF ( .D ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, LED_128_Instance_state1[26]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1441, OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_27__FF_FF ( .D ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, LED_128_Instance_state1[27]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1941, OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_28__FF_FF ( .D ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, LED_128_Instance_state1[28]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1437, OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_29__FF_FF ( .D ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, LED_128_Instance_state1[29]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1937, OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_30__FF_FF ( .D ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, LED_128_Instance_state1[30]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1929, OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_31__FF_FF ( .D ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, LED_128_Instance_state1[31]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1925, OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_32__FF_FF ( .D ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, LED_128_Instance_state1[32]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1433, OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_33__FF_FF ( .D ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, LED_128_Instance_state1[33]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1921, OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_34__FF_FF ( .D ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, LED_128_Instance_state1[34]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1429, OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_35__FF_FF ( .D ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, LED_128_Instance_state1[35]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1425, OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_36__FF_FF ( .D ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, LED_128_Instance_state1[36]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1421, OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_37__FF_FF ( .D ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, LED_128_Instance_state1[37]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1917, OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_38__FF_FF ( .D ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, LED_128_Instance_state1[38]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1913, OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_39__FF_FF ( .D ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, LED_128_Instance_state1[39]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1417, OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_40__FF_FF ( .D ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, LED_128_Instance_state1[40]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1909, OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_41__FF_FF ( .D ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, LED_128_Instance_state1[41]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1905, OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_42__FF_FF ( .D ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, LED_128_Instance_state1[42]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1901, OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_43__FF_FF ( .D ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, LED_128_Instance_state1[43]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1897, OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_44__FF_FF ( .D ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, LED_128_Instance_state1[44]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1893, OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_45__FF_FF ( .D ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, LED_128_Instance_state1[45]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1889, OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_46__FF_FF ( .D ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, LED_128_Instance_state1[46]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1885, OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_47__FF_FF ( .D ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, LED_128_Instance_state1[47]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1881, OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_48__FF_FF ( .D ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, LED_128_Instance_state1[48]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1877, OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_49__FF_FF ( .D ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, LED_128_Instance_state1[49]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1873, OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_50__FF_FF ( .D ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, LED_128_Instance_state1[50]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1865, OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_51__FF_FF ( .D ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, LED_128_Instance_state1[51]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1861, OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_52__FF_FF ( .D ({new_AGEMA_signal_3715, new_AGEMA_signal_3714, LED_128_Instance_state1[52]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1857, OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_53__FF_FF ( .D ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, LED_128_Instance_state1[53]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1853, OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_54__FF_FF ( .D ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, LED_128_Instance_state1[54]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1849, OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_55__FF_FF ( .D ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, LED_128_Instance_state1[55]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1845, OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_56__FF_FF ( .D ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, LED_128_Instance_state1[56]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1841, OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_57__FF_FF ( .D ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, LED_128_Instance_state1[57]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1837, OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_58__FF_FF ( .D ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, LED_128_Instance_state1[58]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1833, OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_59__FF_FF ( .D ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, LED_128_Instance_state1[59]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1829, OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_60__FF_FF ( .D ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, LED_128_Instance_state1[60]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1821, OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_61__FF_FF ( .D ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, LED_128_Instance_state1[61]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1817, OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_62__FF_FF ( .D ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, LED_128_Instance_state1[62]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1813, OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    reg_LMDPL LED_128_Instance_cipherstate_reg_63__FF_FF ( .D ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, LED_128_Instance_state1[63]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (CLK), .Q ({new_AGEMA_signal_1809, OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    reg_sr_LMDPL internal_done_reg_FF_FF ( .D (n15), .clk (CLK), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (OUT_done), .QN () ) ;
endmodule
