/* modified netlist. Source: module CRAFT in file Designs/CRAFT_round-based/AGEMA/CRAFT.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module CRAFT_HPC2_BDDsylvan_ClockGating_d1 (plaintext_s0, key_s0, clk, rst, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input [127:0] key_s1 ;
    input [63:0] plaintext_s1 ;
    input [271:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    output Synch ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1277 ;
    wire signal_1280 ;
    wire signal_1283 ;
    wire signal_1286 ;
    wire signal_1289 ;
    wire signal_1292 ;
    wire signal_1295 ;
    wire signal_1298 ;
    wire signal_1301 ;
    wire signal_1304 ;
    wire signal_1307 ;
    wire signal_1310 ;
    wire signal_1313 ;
    wire signal_1316 ;
    wire signal_1319 ;
    wire signal_1322 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1564 ;
    wire signal_1566 ;
    wire signal_1568 ;
    wire signal_1570 ;
    wire signal_1572 ;
    wire signal_1574 ;
    wire signal_1576 ;
    wire signal_1578 ;
    wire signal_1580 ;
    wire signal_1582 ;
    wire signal_1584 ;
    wire signal_1586 ;
    wire signal_1588 ;
    wire signal_1590 ;
    wire signal_1592 ;
    wire signal_1594 ;
    wire signal_1597 ;
    wire signal_1600 ;
    wire signal_1603 ;
    wire signal_1606 ;
    wire signal_1609 ;
    wire signal_1612 ;
    wire signal_1615 ;
    wire signal_1618 ;
    wire signal_1621 ;
    wire signal_1624 ;
    wire signal_1627 ;
    wire signal_1630 ;
    wire signal_1633 ;
    wire signal_1636 ;
    wire signal_1639 ;
    wire signal_1642 ;
    wire signal_1645 ;
    wire signal_1648 ;
    wire signal_1651 ;
    wire signal_1654 ;
    wire signal_1657 ;
    wire signal_1660 ;
    wire signal_1663 ;
    wire signal_1666 ;
    wire signal_1669 ;
    wire signal_1672 ;
    wire signal_1675 ;
    wire signal_1678 ;
    wire signal_1681 ;
    wire signal_1684 ;
    wire signal_1687 ;
    wire signal_1690 ;
    wire signal_1693 ;
    wire signal_1696 ;
    wire signal_1699 ;
    wire signal_1702 ;
    wire signal_1705 ;
    wire signal_1708 ;
    wire signal_1711 ;
    wire signal_1714 ;
    wire signal_1717 ;
    wire signal_1720 ;
    wire signal_1723 ;
    wire signal_1726 ;
    wire signal_1729 ;
    wire signal_1732 ;
    wire signal_1735 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1788 ;
    wire signal_1790 ;
    wire signal_1792 ;
    wire signal_1794 ;
    wire signal_1796 ;
    wire signal_1798 ;
    wire signal_1800 ;
    wire signal_1802 ;
    wire signal_1804 ;
    wire signal_1806 ;
    wire signal_1808 ;
    wire signal_1810 ;
    wire signal_1812 ;
    wire signal_1814 ;
    wire signal_1816 ;
    wire signal_1818 ;
    wire signal_1820 ;
    wire signal_1822 ;
    wire signal_1824 ;
    wire signal_1826 ;
    wire signal_1828 ;
    wire signal_1830 ;
    wire signal_1832 ;
    wire signal_1834 ;
    wire signal_1836 ;
    wire signal_1838 ;
    wire signal_1840 ;
    wire signal_1842 ;
    wire signal_1844 ;
    wire signal_1846 ;
    wire signal_1848 ;
    wire signal_1850 ;
    wire signal_1852 ;
    wire signal_1854 ;
    wire signal_1856 ;
    wire signal_1858 ;
    wire signal_1860 ;
    wire signal_1862 ;
    wire signal_1864 ;
    wire signal_1866 ;
    wire signal_1868 ;
    wire signal_1870 ;
    wire signal_1872 ;
    wire signal_1874 ;
    wire signal_1876 ;
    wire signal_1878 ;
    wire signal_1880 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2371 ;

    /* cells in depth 0 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_177 ( .a ({signal_1684, signal_894}), .b ({1'b0, signal_266}), .c ({signal_1895, signal_333}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_180 ( .a ({signal_1687, signal_893}), .b ({1'b0, signal_1014}), .c ({signal_1896, signal_335}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_183 ( .a ({signal_1690, signal_892}), .b ({1'b0, signal_1013}), .c ({signal_1897, signal_337}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_186 ( .a ({signal_1693, signal_891}), .b ({1'b0, 1'b0}), .c ({signal_1898, signal_339}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_189 ( .a ({signal_1696, signal_890}), .b ({1'b0, signal_265}), .c ({signal_1899, signal_341}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_192 ( .a ({signal_1699, signal_889}), .b ({1'b0, signal_1011}), .c ({signal_1900, signal_343}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_195 ( .a ({signal_1702, signal_888}), .b ({1'b0, signal_1010}), .c ({signal_1901, signal_345}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_198 ( .a ({signal_1705, signal_887}), .b ({1'b0, signal_1009}), .c ({signal_1902, signal_347}) ) ;
    INV_X1 cell_712 ( .A (signal_1000), .ZN (signal_692) ) ;
    INV_X1 cell_713 ( .A (signal_692), .ZN (signal_693) ) ;
    INV_X1 cell_714 ( .A (signal_692), .ZN (signal_694) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_715 ( .s (signal_1000), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1277, signal_934}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_716 ( .s (signal_693), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1597, signal_933}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_717 ( .s (signal_1000), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1280, signal_932}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_718 ( .s (signal_693), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1600, signal_931}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_719 ( .s (signal_693), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1603, signal_930}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_720 ( .s (signal_693), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({signal_1606, signal_929}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_721 ( .s (signal_693), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({signal_1609, signal_928}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_722 ( .s (signal_693), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({signal_1612, signal_927}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_723 ( .s (signal_693), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1615, signal_926}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_724 ( .s (signal_693), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1618, signal_925}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_725 ( .s (signal_693), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1621, signal_924}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_726 ( .s (signal_693), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1624, signal_923}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_727 ( .s (signal_693), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({signal_1627, signal_922}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_728 ( .s (signal_693), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1630, signal_921}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_729 ( .s (signal_693), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1633, signal_920}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_730 ( .s (signal_693), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1636, signal_919}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_731 ( .s (signal_693), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({signal_1639, signal_918}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_732 ( .s (signal_693), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({signal_1642, signal_917}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_733 ( .s (signal_693), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({signal_1645, signal_916}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_734 ( .s (signal_693), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({signal_1648, signal_915}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_735 ( .s (signal_693), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({signal_1651, signal_914}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_736 ( .s (signal_693), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({signal_1654, signal_913}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_737 ( .s (signal_1000), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({signal_1283, signal_912}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_738 ( .s (signal_1000), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({signal_1286, signal_911}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_739 ( .s (signal_1000), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({signal_1289, signal_910}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_740 ( .s (signal_1000), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({signal_1292, signal_909}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_741 ( .s (signal_1000), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1295, signal_908}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_742 ( .s (signal_1000), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({signal_1298, signal_907}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_743 ( .s (signal_694), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({signal_1657, signal_906}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_744 ( .s (signal_694), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({signal_1660, signal_905}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_745 ( .s (signal_694), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({signal_1663, signal_904}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_746 ( .s (signal_694), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({signal_1666, signal_903}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_747 ( .s (signal_694), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({signal_1669, signal_902}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_748 ( .s (signal_1000), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({signal_1301, signal_901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_749 ( .s (signal_694), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({signal_1672, signal_900}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_750 ( .s (signal_694), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({signal_1675, signal_899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_751 ( .s (signal_1000), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({signal_1304, signal_898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_752 ( .s (signal_694), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({signal_1678, signal_897}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_753 ( .s (signal_694), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({signal_1681, signal_896}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_754 ( .s (signal_1000), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({signal_1307, signal_895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_755 ( .s (signal_694), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({signal_1684, signal_894}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_756 ( .s (signal_694), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({signal_1687, signal_893}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_757 ( .s (signal_694), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({signal_1690, signal_892}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_758 ( .s (signal_694), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({signal_1693, signal_891}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_759 ( .s (signal_694), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({signal_1696, signal_890}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_760 ( .s (signal_694), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({signal_1699, signal_889}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_761 ( .s (signal_694), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({signal_1702, signal_888}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_762 ( .s (signal_694), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({signal_1705, signal_887}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_763 ( .s (signal_694), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({signal_1708, signal_886}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_764 ( .s (signal_694), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({signal_1711, signal_885}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_765 ( .s (signal_694), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({signal_1714, signal_884}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_766 ( .s (signal_694), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({signal_1717, signal_883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_767 ( .s (signal_694), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({signal_1720, signal_882}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_768 ( .s (signal_1000), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({signal_1310, signal_881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_769 ( .s (signal_1000), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({signal_1313, signal_880}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_770 ( .s (signal_694), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({signal_1723, signal_879}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_771 ( .s (signal_1000), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({signal_1316, signal_878}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_772 ( .s (signal_694), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({signal_1726, signal_877}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_773 ( .s (signal_694), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({signal_1729, signal_876}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_774 ( .s (signal_1000), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({signal_1319, signal_875}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_775 ( .s (signal_694), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({signal_1732, signal_874}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_776 ( .s (signal_694), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({signal_1735, signal_873}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_777 ( .s (signal_1000), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({signal_1322, signal_872}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_778 ( .s (signal_694), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({signal_1738, signal_871}) ) ;
    MUX2_X1 cell_779 ( .S (rst), .A (signal_1007), .B (1'b1), .Z (signal_266) ) ;
    MUX2_X1 cell_780 ( .S (rst), .A (signal_1006), .B (1'b0), .Z (signal_1014) ) ;
    MUX2_X1 cell_781 ( .S (rst), .A (signal_1005), .B (1'b0), .Z (signal_1013) ) ;
    MUX2_X1 cell_782 ( .S (rst), .A (signal_1004), .B (1'b1), .Z (signal_265) ) ;
    MUX2_X1 cell_783 ( .S (rst), .A (signal_1003), .B (1'b0), .Z (signal_1011) ) ;
    MUX2_X1 cell_784 ( .S (rst), .A (signal_1002), .B (1'b0), .Z (signal_1010) ) ;
    MUX2_X1 cell_785 ( .S (rst), .A (signal_1001), .B (1'b0), .Z (signal_1009) ) ;
    XOR2_X1 cell_786 ( .A (signal_265), .B (signal_1011), .Z (signal_1008) ) ;
    XOR2_X1 cell_787 ( .A (signal_1014), .B (signal_266), .Z (signal_1012) ) ;
    AND2_X1 cell_802 ( .A1 (signal_1009), .A2 (signal_702), .ZN (signal_267) ) ;
    NOR2_X1 cell_803 ( .A1 (signal_703), .A2 (signal_704), .ZN (signal_702) ) ;
    NAND2_X1 cell_804 ( .A1 (signal_705), .A2 (signal_706), .ZN (signal_704) ) ;
    NOR2_X1 cell_805 ( .A1 (signal_1011), .A2 (signal_1010), .ZN (signal_706) ) ;
    NOR2_X1 cell_806 ( .A1 (signal_1014), .A2 (signal_265), .ZN (signal_705) ) ;
    NAND2_X1 cell_807 ( .A1 (signal_266), .A2 (signal_1013), .ZN (signal_703) ) ;
    MUX2_X1 cell_808 ( .S (rst), .A (signal_1016), .B (1'b0), .Z (signal_1000) ) ;
    MUX2_X1 cell_809 ( .S (rst), .A (signal_1015), .B (1'b0), .Z (signal_999) ) ;
    XNOR2_X1 cell_810 ( .A (signal_707), .B (signal_999), .ZN (signal_1017) ) ;
    XNOR2_X1 cell_811 ( .A (signal_1000), .B (1'b0), .ZN (signal_707) ) ;
    INV_X1 cell_812 ( .A (signal_1000), .ZN (signal_1018) ) ;
    ClockGatingController #(9) cell_1091 ( .clk (clk), .rst (rst), .GatedClk (signal_2371), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_819 ( .s ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[0]), .c ({signal_1228, signal_1019}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_820 ( .s ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[1]), .c ({signal_1229, signal_1020}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_821 ( .s ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[2]), .c ({signal_1231, signal_1021}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_822 ( .s ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[3]), .c ({signal_1232, signal_1022}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_823 ( .s ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[4]), .c ({signal_1234, signal_1023}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_824 ( .s ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[5]), .c ({signal_1235, signal_1024}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_825 ( .s ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[6]), .c ({signal_1237, signal_1025}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_826 ( .s ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[7]), .c ({signal_1238, signal_1026}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_827 ( .s ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[8]), .c ({signal_1240, signal_1027}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_828 ( .s ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[9]), .c ({signal_1241, signal_1028}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_829 ( .s ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[10]), .c ({signal_1243, signal_1029}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_830 ( .s ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[11]), .c ({signal_1244, signal_1030}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_831 ( .s ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[12]), .c ({signal_1246, signal_1031}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_832 ( .s ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[13]), .c ({signal_1247, signal_1032}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_833 ( .s ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[14]), .c ({signal_1249, signal_1033}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_834 ( .s ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[15]), .c ({signal_1250, signal_1034}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_835 ( .s ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[16]), .c ({signal_1252, signal_1035}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_836 ( .s ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[17]), .c ({signal_1253, signal_1036}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_837 ( .s ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[18]), .c ({signal_1255, signal_1037}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_838 ( .s ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[19]), .c ({signal_1256, signal_1038}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_839 ( .s ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[20]), .c ({signal_1258, signal_1039}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_840 ( .s ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[21]), .c ({signal_1259, signal_1040}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_841 ( .s ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[22]), .c ({signal_1261, signal_1041}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_842 ( .s ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[23]), .c ({signal_1262, signal_1042}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_843 ( .s ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[24]), .c ({signal_1264, signal_1043}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_844 ( .s ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[25]), .c ({signal_1265, signal_1044}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_845 ( .s ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[26]), .c ({signal_1267, signal_1045}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_846 ( .s ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[27]), .c ({signal_1268, signal_1046}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_847 ( .s ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[28]), .c ({signal_1270, signal_1047}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_848 ( .s ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[29]), .c ({signal_1271, signal_1048}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_849 ( .s ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[30]), .c ({signal_1273, signal_1049}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_850 ( .s ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[31]), .c ({signal_1274, signal_1050}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_851 ( .s ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({1'b0, 1'b1}), .a ({signal_1228, signal_1019}), .clk (clk), .r (Fresh[32]), .c ({signal_1324, signal_1051}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_852 ( .s ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_1229, signal_1020}), .a ({signal_1228, signal_1019}), .clk (clk), .r (Fresh[33]), .c ({signal_1325, signal_1052}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_853 ( .s ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_1228, signal_1019}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[34]), .c ({signal_1326, signal_1053}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_854 ( .s ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({1'b0, 1'b0}), .a ({signal_1228, signal_1019}), .clk (clk), .r (Fresh[35]), .c ({signal_1327, signal_1054}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_855 ( .s ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_1229, signal_1020}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[36]), .c ({signal_1328, signal_1055}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_856 ( .s ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({1'b0, 1'b1}), .a ({signal_1231, signal_1021}), .clk (clk), .r (Fresh[37]), .c ({signal_1330, signal_1056}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_857 ( .s ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({signal_1232, signal_1022}), .a ({signal_1231, signal_1021}), .clk (clk), .r (Fresh[38]), .c ({signal_1331, signal_1057}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_858 ( .s ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({signal_1231, signal_1021}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[39]), .c ({signal_1332, signal_1058}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_859 ( .s ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({1'b0, 1'b0}), .a ({signal_1231, signal_1021}), .clk (clk), .r (Fresh[40]), .c ({signal_1333, signal_1059}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_860 ( .s ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({signal_1232, signal_1022}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[41]), .c ({signal_1334, signal_1060}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_861 ( .s ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({1'b0, 1'b1}), .a ({signal_1234, signal_1023}), .clk (clk), .r (Fresh[42]), .c ({signal_1336, signal_1061}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_862 ( .s ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({signal_1235, signal_1024}), .a ({signal_1234, signal_1023}), .clk (clk), .r (Fresh[43]), .c ({signal_1337, signal_1062}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_863 ( .s ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({signal_1234, signal_1023}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[44]), .c ({signal_1338, signal_1063}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_864 ( .s ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({1'b0, 1'b0}), .a ({signal_1234, signal_1023}), .clk (clk), .r (Fresh[45]), .c ({signal_1339, signal_1064}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_865 ( .s ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({signal_1235, signal_1024}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[46]), .c ({signal_1340, signal_1065}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_866 ( .s ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({1'b0, 1'b1}), .a ({signal_1237, signal_1025}), .clk (clk), .r (Fresh[47]), .c ({signal_1342, signal_1066}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_867 ( .s ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({signal_1238, signal_1026}), .a ({signal_1237, signal_1025}), .clk (clk), .r (Fresh[48]), .c ({signal_1343, signal_1067}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_868 ( .s ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({signal_1237, signal_1025}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[49]), .c ({signal_1344, signal_1068}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_869 ( .s ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({1'b0, 1'b0}), .a ({signal_1237, signal_1025}), .clk (clk), .r (Fresh[50]), .c ({signal_1345, signal_1069}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_870 ( .s ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({signal_1238, signal_1026}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[51]), .c ({signal_1346, signal_1070}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_871 ( .s ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({1'b0, 1'b1}), .a ({signal_1240, signal_1027}), .clk (clk), .r (Fresh[52]), .c ({signal_1348, signal_1071}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_872 ( .s ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({signal_1241, signal_1028}), .a ({signal_1240, signal_1027}), .clk (clk), .r (Fresh[53]), .c ({signal_1349, signal_1072}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_873 ( .s ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({signal_1240, signal_1027}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[54]), .c ({signal_1350, signal_1073}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_874 ( .s ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({1'b0, 1'b0}), .a ({signal_1240, signal_1027}), .clk (clk), .r (Fresh[55]), .c ({signal_1351, signal_1074}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_875 ( .s ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({signal_1241, signal_1028}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[56]), .c ({signal_1352, signal_1075}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_876 ( .s ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({1'b0, 1'b1}), .a ({signal_1243, signal_1029}), .clk (clk), .r (Fresh[57]), .c ({signal_1354, signal_1076}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_877 ( .s ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({signal_1244, signal_1030}), .a ({signal_1243, signal_1029}), .clk (clk), .r (Fresh[58]), .c ({signal_1355, signal_1077}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_878 ( .s ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({signal_1243, signal_1029}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[59]), .c ({signal_1356, signal_1078}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_879 ( .s ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({1'b0, 1'b0}), .a ({signal_1243, signal_1029}), .clk (clk), .r (Fresh[60]), .c ({signal_1357, signal_1079}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_880 ( .s ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({signal_1244, signal_1030}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[61]), .c ({signal_1358, signal_1080}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_881 ( .s ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({1'b0, 1'b1}), .a ({signal_1246, signal_1031}), .clk (clk), .r (Fresh[62]), .c ({signal_1360, signal_1081}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_882 ( .s ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({signal_1247, signal_1032}), .a ({signal_1246, signal_1031}), .clk (clk), .r (Fresh[63]), .c ({signal_1361, signal_1082}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_883 ( .s ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({signal_1246, signal_1031}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[64]), .c ({signal_1362, signal_1083}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_884 ( .s ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({1'b0, 1'b0}), .a ({signal_1246, signal_1031}), .clk (clk), .r (Fresh[65]), .c ({signal_1363, signal_1084}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_885 ( .s ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({signal_1247, signal_1032}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[66]), .c ({signal_1364, signal_1085}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_886 ( .s ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({1'b0, 1'b1}), .a ({signal_1249, signal_1033}), .clk (clk), .r (Fresh[67]), .c ({signal_1366, signal_1086}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_887 ( .s ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({signal_1250, signal_1034}), .a ({signal_1249, signal_1033}), .clk (clk), .r (Fresh[68]), .c ({signal_1367, signal_1087}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_888 ( .s ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({signal_1249, signal_1033}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[69]), .c ({signal_1368, signal_1088}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_889 ( .s ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({1'b0, 1'b0}), .a ({signal_1249, signal_1033}), .clk (clk), .r (Fresh[70]), .c ({signal_1369, signal_1089}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_890 ( .s ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({signal_1250, signal_1034}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[71]), .c ({signal_1370, signal_1090}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_891 ( .s ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({1'b0, 1'b1}), .a ({signal_1252, signal_1035}), .clk (clk), .r (Fresh[72]), .c ({signal_1372, signal_1091}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_892 ( .s ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({signal_1253, signal_1036}), .a ({signal_1252, signal_1035}), .clk (clk), .r (Fresh[73]), .c ({signal_1373, signal_1092}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_893 ( .s ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({signal_1252, signal_1035}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[74]), .c ({signal_1374, signal_1093}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_894 ( .s ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({1'b0, 1'b0}), .a ({signal_1252, signal_1035}), .clk (clk), .r (Fresh[75]), .c ({signal_1375, signal_1094}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_895 ( .s ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({signal_1253, signal_1036}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[76]), .c ({signal_1376, signal_1095}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_896 ( .s ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({1'b0, 1'b1}), .a ({signal_1255, signal_1037}), .clk (clk), .r (Fresh[77]), .c ({signal_1378, signal_1096}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_897 ( .s ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_1256, signal_1038}), .a ({signal_1255, signal_1037}), .clk (clk), .r (Fresh[78]), .c ({signal_1379, signal_1097}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_898 ( .s ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_1255, signal_1037}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[79]), .c ({signal_1380, signal_1098}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_899 ( .s ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({1'b0, 1'b0}), .a ({signal_1255, signal_1037}), .clk (clk), .r (Fresh[80]), .c ({signal_1381, signal_1099}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_900 ( .s ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_1256, signal_1038}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[81]), .c ({signal_1382, signal_1100}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_901 ( .s ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({1'b0, 1'b1}), .a ({signal_1258, signal_1039}), .clk (clk), .r (Fresh[82]), .c ({signal_1384, signal_1101}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_902 ( .s ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({signal_1259, signal_1040}), .a ({signal_1258, signal_1039}), .clk (clk), .r (Fresh[83]), .c ({signal_1385, signal_1102}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_903 ( .s ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({signal_1258, signal_1039}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[84]), .c ({signal_1386, signal_1103}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_904 ( .s ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({1'b0, 1'b0}), .a ({signal_1258, signal_1039}), .clk (clk), .r (Fresh[85]), .c ({signal_1387, signal_1104}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_905 ( .s ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({signal_1259, signal_1040}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[86]), .c ({signal_1388, signal_1105}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_906 ( .s ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({1'b0, 1'b1}), .a ({signal_1261, signal_1041}), .clk (clk), .r (Fresh[87]), .c ({signal_1390, signal_1106}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_907 ( .s ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({signal_1262, signal_1042}), .a ({signal_1261, signal_1041}), .clk (clk), .r (Fresh[88]), .c ({signal_1391, signal_1107}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_908 ( .s ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({signal_1261, signal_1041}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[89]), .c ({signal_1392, signal_1108}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_909 ( .s ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({1'b0, 1'b0}), .a ({signal_1261, signal_1041}), .clk (clk), .r (Fresh[90]), .c ({signal_1393, signal_1109}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_910 ( .s ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({signal_1262, signal_1042}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[91]), .c ({signal_1394, signal_1110}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_911 ( .s ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({1'b0, 1'b1}), .a ({signal_1264, signal_1043}), .clk (clk), .r (Fresh[92]), .c ({signal_1396, signal_1111}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_912 ( .s ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({signal_1265, signal_1044}), .a ({signal_1264, signal_1043}), .clk (clk), .r (Fresh[93]), .c ({signal_1397, signal_1112}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_913 ( .s ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({signal_1264, signal_1043}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[94]), .c ({signal_1398, signal_1113}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_914 ( .s ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({1'b0, 1'b0}), .a ({signal_1264, signal_1043}), .clk (clk), .r (Fresh[95]), .c ({signal_1399, signal_1114}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_915 ( .s ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({signal_1265, signal_1044}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[96]), .c ({signal_1400, signal_1115}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_916 ( .s ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({1'b0, 1'b1}), .a ({signal_1267, signal_1045}), .clk (clk), .r (Fresh[97]), .c ({signal_1402, signal_1116}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_917 ( .s ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({signal_1268, signal_1046}), .a ({signal_1267, signal_1045}), .clk (clk), .r (Fresh[98]), .c ({signal_1403, signal_1117}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_918 ( .s ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({signal_1267, signal_1045}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[99]), .c ({signal_1404, signal_1118}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_919 ( .s ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({1'b0, 1'b0}), .a ({signal_1267, signal_1045}), .clk (clk), .r (Fresh[100]), .c ({signal_1405, signal_1119}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_920 ( .s ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({signal_1268, signal_1046}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[101]), .c ({signal_1406, signal_1120}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_921 ( .s ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({1'b0, 1'b1}), .a ({signal_1270, signal_1047}), .clk (clk), .r (Fresh[102]), .c ({signal_1408, signal_1121}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_922 ( .s ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({signal_1271, signal_1048}), .a ({signal_1270, signal_1047}), .clk (clk), .r (Fresh[103]), .c ({signal_1409, signal_1122}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_923 ( .s ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({signal_1270, signal_1047}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[104]), .c ({signal_1410, signal_1123}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_924 ( .s ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({1'b0, 1'b0}), .a ({signal_1270, signal_1047}), .clk (clk), .r (Fresh[105]), .c ({signal_1411, signal_1124}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_925 ( .s ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({signal_1271, signal_1048}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[106]), .c ({signal_1412, signal_1125}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_926 ( .s ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({1'b0, 1'b1}), .a ({signal_1273, signal_1049}), .clk (clk), .r (Fresh[107]), .c ({signal_1414, signal_1126}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_927 ( .s ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({signal_1274, signal_1050}), .a ({signal_1273, signal_1049}), .clk (clk), .r (Fresh[108]), .c ({signal_1415, signal_1127}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_928 ( .s ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({signal_1273, signal_1049}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[109]), .c ({signal_1416, signal_1128}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_929 ( .s ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_1273, signal_1049}), .clk (clk), .r (Fresh[110]), .c ({signal_1417, signal_1129}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_930 ( .s ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({signal_1274, signal_1050}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[111]), .c ({signal_1418, signal_1130}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1 ( .s (rst), .b ({signal_1423, signal_773}), .a ({plaintext_s1[1], plaintext_s0[1]}), .c ({signal_1564, signal_869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_5 ( .s (rst), .b ({signal_1432, signal_769}), .a ({plaintext_s1[5], plaintext_s0[5]}), .c ({signal_1566, signal_865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_9 ( .s (rst), .b ({signal_1441, signal_765}), .a ({plaintext_s1[9], plaintext_s0[9]}), .c ({signal_1568, signal_861}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_13 ( .s (rst), .b ({signal_1450, signal_761}), .a ({plaintext_s1[13], plaintext_s0[13]}), .c ({signal_1570, signal_857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_17 ( .s (rst), .b ({signal_1459, signal_757}), .a ({plaintext_s1[17], plaintext_s0[17]}), .c ({signal_1572, signal_853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_21 ( .s (rst), .b ({signal_1468, signal_753}), .a ({plaintext_s1[21], plaintext_s0[21]}), .c ({signal_1574, signal_849}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_25 ( .s (rst), .b ({signal_1477, signal_749}), .a ({plaintext_s1[25], plaintext_s0[25]}), .c ({signal_1576, signal_845}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_29 ( .s (rst), .b ({signal_1486, signal_745}), .a ({plaintext_s1[29], plaintext_s0[29]}), .c ({signal_1578, signal_841}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_33 ( .s (rst), .b ({signal_1495, signal_741}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({signal_1580, signal_805}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_37 ( .s (rst), .b ({signal_1504, signal_737}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({signal_1582, signal_801}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_41 ( .s (rst), .b ({signal_1513, signal_733}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({signal_1584, signal_797}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_45 ( .s (rst), .b ({signal_1522, signal_729}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({signal_1586, signal_793}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_49 ( .s (rst), .b ({signal_1531, signal_725}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({signal_1588, signal_789}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_53 ( .s (rst), .b ({signal_1540, signal_721}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({signal_1590, signal_785}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_57 ( .s (rst), .b ({signal_1549, signal_717}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({signal_1592, signal_781}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_61 ( .s (rst), .b ({signal_1558, signal_713}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({signal_1594, signal_777}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_69 ( .a ({signal_1884, signal_271}), .b ({signal_1883, signal_272}), .c ({signal_1914, signal_821}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_70 ( .a ({signal_1572, signal_853}), .b ({signal_1564, signal_869}), .c ({signal_1883, signal_272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_71 ( .a ({1'b0, 1'b0}), .b ({signal_1588, signal_789}), .c ({signal_1884, signal_271}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_72 ( .a ({signal_1885, signal_273}), .b ({signal_1564, signal_869}), .c ({signal_1915, signal_837}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_73 ( .a ({1'b0, 1'b0}), .b ({signal_1580, signal_805}), .c ({signal_1885, signal_273}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_89 ( .a ({signal_1887, signal_283}), .b ({signal_1886, signal_284}), .c ({signal_1925, signal_817}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_90 ( .a ({signal_1574, signal_849}), .b ({signal_1566, signal_865}), .c ({signal_1886, signal_284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_91 ( .a ({1'b0, 1'b0}), .b ({signal_1590, signal_785}), .c ({signal_1887, signal_283}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_92 ( .a ({signal_1888, signal_285}), .b ({signal_1566, signal_865}), .c ({signal_1926, signal_833}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_93 ( .a ({1'b0, 1'b0}), .b ({signal_1582, signal_801}), .c ({signal_1888, signal_285}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_109 ( .a ({signal_1890, signal_295}), .b ({signal_1889, signal_296}), .c ({signal_1936, signal_813}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_110 ( .a ({signal_1576, signal_845}), .b ({signal_1568, signal_861}), .c ({signal_1889, signal_296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_111 ( .a ({1'b0, 1'b0}), .b ({signal_1592, signal_781}), .c ({signal_1890, signal_295}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_112 ( .a ({signal_1891, signal_297}), .b ({signal_1568, signal_861}), .c ({signal_1937, signal_829}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_113 ( .a ({1'b0, 1'b0}), .b ({signal_1584, signal_797}), .c ({signal_1891, signal_297}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_129 ( .a ({signal_1893, signal_307}), .b ({signal_1892, signal_308}), .c ({signal_1947, signal_809}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_130 ( .a ({signal_1578, signal_841}), .b ({signal_1570, signal_857}), .c ({signal_1892, signal_308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_131 ( .a ({1'b0, 1'b0}), .b ({signal_1594, signal_777}), .c ({signal_1893, signal_307}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_132 ( .a ({signal_1894, signal_309}), .b ({signal_1570, signal_857}), .c ({signal_1948, signal_825}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_133 ( .a ({1'b0, 1'b0}), .b ({signal_1586, signal_793}), .c ({signal_1894, signal_309}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_146 ( .a ({signal_2011, signal_317}), .b ({signal_1711, signal_885}), .c ({signal_2044, signal_949}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_147 ( .a ({1'b0, 1'b0}), .b ({signal_1914, signal_821}), .c ({signal_2011, signal_317}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_154 ( .a ({signal_2012, signal_321}), .b ({signal_1310, signal_881}), .c ({signal_2048, signal_945}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_155 ( .a ({1'b0, 1'b0}), .b ({signal_1925, signal_817}), .c ({signal_2012, signal_321}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_162 ( .a ({signal_2013, signal_325}), .b ({signal_1726, signal_877}), .c ({signal_2052, signal_941}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_163 ( .a ({1'b0, 1'b0}), .b ({signal_1936, signal_813}), .c ({signal_2013, signal_325}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_170 ( .a ({signal_2014, signal_329}), .b ({signal_1735, signal_873}), .c ({signal_2056, signal_937}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_171 ( .a ({1'b0, 1'b0}), .b ({signal_1947, signal_809}), .c ({signal_2014, signal_329}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_179 ( .a ({signal_2015, signal_334}), .b ({signal_1896, signal_335}), .c ({signal_2060, signal_957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_181 ( .a ({1'b0, 1'b0}), .b ({signal_1937, signal_829}), .c ({signal_2015, signal_334}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_191 ( .a ({signal_2016, signal_342}), .b ({signal_1900, signal_343}), .c ({signal_2064, signal_953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_193 ( .a ({1'b0, 1'b0}), .b ({signal_1948, signal_825}), .c ({signal_2016, signal_342}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_202 ( .a ({signal_1903, signal_349}), .b ({signal_1597, signal_933}), .c ({signal_1956, signal_997}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_203 ( .a ({1'b0, 1'b0}), .b ({signal_1564, signal_869}), .c ({signal_1903, signal_349}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_210 ( .a ({signal_1904, signal_353}), .b ({signal_1606, signal_929}), .c ({signal_1960, signal_993}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_211 ( .a ({1'b0, 1'b0}), .b ({signal_1566, signal_865}), .c ({signal_1904, signal_353}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_218 ( .a ({signal_1905, signal_357}), .b ({signal_1618, signal_925}), .c ({signal_1964, signal_989}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_219 ( .a ({1'b0, 1'b0}), .b ({signal_1568, signal_861}), .c ({signal_1905, signal_357}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_226 ( .a ({signal_1906, signal_361}), .b ({signal_1630, signal_921}), .c ({signal_1968, signal_985}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_227 ( .a ({1'b0, 1'b0}), .b ({signal_1570, signal_857}), .c ({signal_1906, signal_361}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_234 ( .a ({signal_1907, signal_365}), .b ({signal_1642, signal_917}), .c ({signal_1972, signal_981}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_235 ( .a ({1'b0, 1'b0}), .b ({signal_1572, signal_853}), .c ({signal_1907, signal_365}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_242 ( .a ({signal_1908, signal_369}), .b ({signal_1654, signal_913}), .c ({signal_1976, signal_977}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_243 ( .a ({1'b0, 1'b0}), .b ({signal_1574, signal_849}), .c ({signal_1908, signal_369}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_250 ( .a ({signal_1909, signal_373}), .b ({signal_1292, signal_909}), .c ({signal_1980, signal_973}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_251 ( .a ({1'b0, 1'b0}), .b ({signal_1576, signal_845}), .c ({signal_1909, signal_373}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_258 ( .a ({signal_1910, signal_377}), .b ({signal_1660, signal_905}), .c ({signal_1984, signal_969}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_259 ( .a ({1'b0, 1'b0}), .b ({signal_1578, signal_841}), .c ({signal_1910, signal_377}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_266 ( .a ({signal_2041, signal_381}), .b ({signal_1301, signal_901}), .c ({signal_2068, signal_965}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_267 ( .a ({1'b0, 1'b0}), .b ({signal_1915, signal_837}), .c ({signal_2041, signal_381}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_274 ( .a ({signal_2042, signal_385}), .b ({signal_1678, signal_897}), .c ({signal_2072, signal_961}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_275 ( .a ({1'b0, 1'b0}), .b ({signal_1926, signal_833}), .c ({signal_2042, signal_385}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_931 ( .s ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_1325, signal_1052}), .a ({signal_1324, signal_1051}), .clk (clk), .r (Fresh[112]), .c ({signal_1420, signal_1131}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_932 ( .s ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({1'b0, 1'b0}), .a ({signal_1324, signal_1051}), .clk (clk), .r (Fresh[113]), .c ({signal_1421, signal_1132}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_933 ( .s ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_1327, signal_1054}), .a ({signal_1326, signal_1053}), .clk (clk), .r (Fresh[114]), .c ({signal_1423, signal_773}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_934 ( .s ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({1'b0, 1'b0}), .a ({signal_1328, signal_1055}), .clk (clk), .r (Fresh[115]), .c ({signal_1424, signal_1133}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_935 ( .s ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_1228, signal_1019}), .a ({signal_1326, signal_1053}), .clk (clk), .r (Fresh[116]), .c ({signal_1425, signal_1134}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_936 ( .s ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_1324, signal_1051}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[117]), .c ({signal_1426, signal_1135}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_937 ( .s ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_1324, signal_1051}), .a ({signal_1228, signal_1019}), .clk (clk), .r (Fresh[118]), .c ({signal_1427, signal_1136}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_938 ( .s ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({signal_1331, signal_1057}), .a ({signal_1330, signal_1056}), .clk (clk), .r (Fresh[119]), .c ({signal_1429, signal_1137}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_939 ( .s ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({1'b0, 1'b0}), .a ({signal_1330, signal_1056}), .clk (clk), .r (Fresh[120]), .c ({signal_1430, signal_1138}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_940 ( .s ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_1333, signal_1059}), .a ({signal_1332, signal_1058}), .clk (clk), .r (Fresh[121]), .c ({signal_1432, signal_769}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_941 ( .s ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({1'b0, 1'b0}), .a ({signal_1334, signal_1060}), .clk (clk), .r (Fresh[122]), .c ({signal_1433, signal_1139}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_942 ( .s ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({signal_1231, signal_1021}), .a ({signal_1332, signal_1058}), .clk (clk), .r (Fresh[123]), .c ({signal_1434, signal_1140}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_943 ( .s ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({signal_1330, signal_1056}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[124]), .c ({signal_1435, signal_1141}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_944 ( .s ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({signal_1330, signal_1056}), .a ({signal_1231, signal_1021}), .clk (clk), .r (Fresh[125]), .c ({signal_1436, signal_1142}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_945 ( .s ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({signal_1337, signal_1062}), .a ({signal_1336, signal_1061}), .clk (clk), .r (Fresh[126]), .c ({signal_1438, signal_1143}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_946 ( .s ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({1'b0, 1'b0}), .a ({signal_1336, signal_1061}), .clk (clk), .r (Fresh[127]), .c ({signal_1439, signal_1144}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_947 ( .s ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_1339, signal_1064}), .a ({signal_1338, signal_1063}), .clk (clk), .r (Fresh[128]), .c ({signal_1441, signal_765}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_948 ( .s ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({1'b0, 1'b0}), .a ({signal_1340, signal_1065}), .clk (clk), .r (Fresh[129]), .c ({signal_1442, signal_1145}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_949 ( .s ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({signal_1234, signal_1023}), .a ({signal_1338, signal_1063}), .clk (clk), .r (Fresh[130]), .c ({signal_1443, signal_1146}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_950 ( .s ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({signal_1336, signal_1061}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[131]), .c ({signal_1444, signal_1147}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_951 ( .s ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({signal_1336, signal_1061}), .a ({signal_1234, signal_1023}), .clk (clk), .r (Fresh[132]), .c ({signal_1445, signal_1148}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_952 ( .s ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_1343, signal_1067}), .a ({signal_1342, signal_1066}), .clk (clk), .r (Fresh[133]), .c ({signal_1447, signal_1149}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_953 ( .s ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({1'b0, 1'b0}), .a ({signal_1342, signal_1066}), .clk (clk), .r (Fresh[134]), .c ({signal_1448, signal_1150}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_954 ( .s ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_1345, signal_1069}), .a ({signal_1344, signal_1068}), .clk (clk), .r (Fresh[135]), .c ({signal_1450, signal_761}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_955 ( .s ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({1'b0, 1'b0}), .a ({signal_1346, signal_1070}), .clk (clk), .r (Fresh[136]), .c ({signal_1451, signal_1151}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_956 ( .s ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_1237, signal_1025}), .a ({signal_1344, signal_1068}), .clk (clk), .r (Fresh[137]), .c ({signal_1452, signal_1152}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_957 ( .s ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_1342, signal_1066}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[138]), .c ({signal_1453, signal_1153}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_958 ( .s ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_1342, signal_1066}), .a ({signal_1237, signal_1025}), .clk (clk), .r (Fresh[139]), .c ({signal_1454, signal_1154}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_959 ( .s ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({signal_1349, signal_1072}), .a ({signal_1348, signal_1071}), .clk (clk), .r (Fresh[140]), .c ({signal_1456, signal_1155}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_960 ( .s ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({1'b0, 1'b0}), .a ({signal_1348, signal_1071}), .clk (clk), .r (Fresh[141]), .c ({signal_1457, signal_1156}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_961 ( .s ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_1351, signal_1074}), .a ({signal_1350, signal_1073}), .clk (clk), .r (Fresh[142]), .c ({signal_1459, signal_757}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_962 ( .s ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({1'b0, 1'b0}), .a ({signal_1352, signal_1075}), .clk (clk), .r (Fresh[143]), .c ({signal_1460, signal_1157}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_963 ( .s ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({signal_1240, signal_1027}), .a ({signal_1350, signal_1073}), .clk (clk), .r (Fresh[144]), .c ({signal_1461, signal_1158}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_964 ( .s ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({signal_1348, signal_1071}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[145]), .c ({signal_1462, signal_1159}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_965 ( .s ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({signal_1348, signal_1071}), .a ({signal_1240, signal_1027}), .clk (clk), .r (Fresh[146]), .c ({signal_1463, signal_1160}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_966 ( .s ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({signal_1355, signal_1077}), .a ({signal_1354, signal_1076}), .clk (clk), .r (Fresh[147]), .c ({signal_1465, signal_1161}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_967 ( .s ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({1'b0, 1'b0}), .a ({signal_1354, signal_1076}), .clk (clk), .r (Fresh[148]), .c ({signal_1466, signal_1162}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_968 ( .s ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_1357, signal_1079}), .a ({signal_1356, signal_1078}), .clk (clk), .r (Fresh[149]), .c ({signal_1468, signal_753}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_969 ( .s ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({1'b0, 1'b0}), .a ({signal_1358, signal_1080}), .clk (clk), .r (Fresh[150]), .c ({signal_1469, signal_1163}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_970 ( .s ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({signal_1243, signal_1029}), .a ({signal_1356, signal_1078}), .clk (clk), .r (Fresh[151]), .c ({signal_1470, signal_1164}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_971 ( .s ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({signal_1354, signal_1076}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[152]), .c ({signal_1471, signal_1165}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_972 ( .s ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({signal_1354, signal_1076}), .a ({signal_1243, signal_1029}), .clk (clk), .r (Fresh[153]), .c ({signal_1472, signal_1166}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_973 ( .s ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({signal_1361, signal_1082}), .a ({signal_1360, signal_1081}), .clk (clk), .r (Fresh[154]), .c ({signal_1474, signal_1167}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_974 ( .s ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({1'b0, 1'b0}), .a ({signal_1360, signal_1081}), .clk (clk), .r (Fresh[155]), .c ({signal_1475, signal_1168}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_975 ( .s ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_1363, signal_1084}), .a ({signal_1362, signal_1083}), .clk (clk), .r (Fresh[156]), .c ({signal_1477, signal_749}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_976 ( .s ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({1'b0, 1'b0}), .a ({signal_1364, signal_1085}), .clk (clk), .r (Fresh[157]), .c ({signal_1478, signal_1169}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_977 ( .s ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({signal_1246, signal_1031}), .a ({signal_1362, signal_1083}), .clk (clk), .r (Fresh[158]), .c ({signal_1479, signal_1170}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_978 ( .s ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({signal_1360, signal_1081}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[159]), .c ({signal_1480, signal_1171}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_979 ( .s ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({signal_1360, signal_1081}), .a ({signal_1246, signal_1031}), .clk (clk), .r (Fresh[160]), .c ({signal_1481, signal_1172}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_980 ( .s ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({signal_1367, signal_1087}), .a ({signal_1366, signal_1086}), .clk (clk), .r (Fresh[161]), .c ({signal_1483, signal_1173}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_981 ( .s ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({1'b0, 1'b0}), .a ({signal_1366, signal_1086}), .clk (clk), .r (Fresh[162]), .c ({signal_1484, signal_1174}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_982 ( .s ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_1369, signal_1089}), .a ({signal_1368, signal_1088}), .clk (clk), .r (Fresh[163]), .c ({signal_1486, signal_745}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_983 ( .s ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({1'b0, 1'b0}), .a ({signal_1370, signal_1090}), .clk (clk), .r (Fresh[164]), .c ({signal_1487, signal_1175}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_984 ( .s ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({signal_1249, signal_1033}), .a ({signal_1368, signal_1088}), .clk (clk), .r (Fresh[165]), .c ({signal_1488, signal_1176}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_985 ( .s ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({signal_1366, signal_1086}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[166]), .c ({signal_1489, signal_1177}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_986 ( .s ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({signal_1366, signal_1086}), .a ({signal_1249, signal_1033}), .clk (clk), .r (Fresh[167]), .c ({signal_1490, signal_1178}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_987 ( .s ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({signal_1373, signal_1092}), .a ({signal_1372, signal_1091}), .clk (clk), .r (Fresh[168]), .c ({signal_1492, signal_1179}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_988 ( .s ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({1'b0, 1'b0}), .a ({signal_1372, signal_1091}), .clk (clk), .r (Fresh[169]), .c ({signal_1493, signal_1180}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_989 ( .s ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_1375, signal_1094}), .a ({signal_1374, signal_1093}), .clk (clk), .r (Fresh[170]), .c ({signal_1495, signal_741}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_990 ( .s ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({1'b0, 1'b0}), .a ({signal_1376, signal_1095}), .clk (clk), .r (Fresh[171]), .c ({signal_1496, signal_1181}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_991 ( .s ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({signal_1252, signal_1035}), .a ({signal_1374, signal_1093}), .clk (clk), .r (Fresh[172]), .c ({signal_1497, signal_1182}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_992 ( .s ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({signal_1372, signal_1091}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[173]), .c ({signal_1498, signal_1183}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_993 ( .s ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({signal_1372, signal_1091}), .a ({signal_1252, signal_1035}), .clk (clk), .r (Fresh[174]), .c ({signal_1499, signal_1184}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_994 ( .s ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_1379, signal_1097}), .a ({signal_1378, signal_1096}), .clk (clk), .r (Fresh[175]), .c ({signal_1501, signal_1185}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_995 ( .s ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({1'b0, 1'b0}), .a ({signal_1378, signal_1096}), .clk (clk), .r (Fresh[176]), .c ({signal_1502, signal_1186}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_996 ( .s ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_1381, signal_1099}), .a ({signal_1380, signal_1098}), .clk (clk), .r (Fresh[177]), .c ({signal_1504, signal_737}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_997 ( .s ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({1'b0, 1'b0}), .a ({signal_1382, signal_1100}), .clk (clk), .r (Fresh[178]), .c ({signal_1505, signal_1187}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_998 ( .s ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_1255, signal_1037}), .a ({signal_1380, signal_1098}), .clk (clk), .r (Fresh[179]), .c ({signal_1506, signal_1188}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_999 ( .s ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_1378, signal_1096}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[180]), .c ({signal_1507, signal_1189}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1000 ( .s ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_1378, signal_1096}), .a ({signal_1255, signal_1037}), .clk (clk), .r (Fresh[181]), .c ({signal_1508, signal_1190}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1001 ( .s ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_1385, signal_1102}), .a ({signal_1384, signal_1101}), .clk (clk), .r (Fresh[182]), .c ({signal_1510, signal_1191}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1002 ( .s ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({1'b0, 1'b0}), .a ({signal_1384, signal_1101}), .clk (clk), .r (Fresh[183]), .c ({signal_1511, signal_1192}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1003 ( .s ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_1387, signal_1104}), .a ({signal_1386, signal_1103}), .clk (clk), .r (Fresh[184]), .c ({signal_1513, signal_733}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1004 ( .s ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({1'b0, 1'b0}), .a ({signal_1388, signal_1105}), .clk (clk), .r (Fresh[185]), .c ({signal_1514, signal_1193}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1005 ( .s ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_1258, signal_1039}), .a ({signal_1386, signal_1103}), .clk (clk), .r (Fresh[186]), .c ({signal_1515, signal_1194}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1006 ( .s ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_1384, signal_1101}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[187]), .c ({signal_1516, signal_1195}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1007 ( .s ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_1384, signal_1101}), .a ({signal_1258, signal_1039}), .clk (clk), .r (Fresh[188]), .c ({signal_1517, signal_1196}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1008 ( .s ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({signal_1391, signal_1107}), .a ({signal_1390, signal_1106}), .clk (clk), .r (Fresh[189]), .c ({signal_1519, signal_1197}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1009 ( .s ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({1'b0, 1'b0}), .a ({signal_1390, signal_1106}), .clk (clk), .r (Fresh[190]), .c ({signal_1520, signal_1198}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1010 ( .s ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_1393, signal_1109}), .a ({signal_1392, signal_1108}), .clk (clk), .r (Fresh[191]), .c ({signal_1522, signal_729}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1011 ( .s ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({1'b0, 1'b0}), .a ({signal_1394, signal_1110}), .clk (clk), .r (Fresh[192]), .c ({signal_1523, signal_1199}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1012 ( .s ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({signal_1261, signal_1041}), .a ({signal_1392, signal_1108}), .clk (clk), .r (Fresh[193]), .c ({signal_1524, signal_1200}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1013 ( .s ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({signal_1390, signal_1106}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[194]), .c ({signal_1525, signal_1201}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1014 ( .s ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({signal_1390, signal_1106}), .a ({signal_1261, signal_1041}), .clk (clk), .r (Fresh[195]), .c ({signal_1526, signal_1202}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1015 ( .s ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({signal_1397, signal_1112}), .a ({signal_1396, signal_1111}), .clk (clk), .r (Fresh[196]), .c ({signal_1528, signal_1203}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1016 ( .s ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({1'b0, 1'b0}), .a ({signal_1396, signal_1111}), .clk (clk), .r (Fresh[197]), .c ({signal_1529, signal_1204}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1017 ( .s ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_1399, signal_1114}), .a ({signal_1398, signal_1113}), .clk (clk), .r (Fresh[198]), .c ({signal_1531, signal_725}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1018 ( .s ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({1'b0, 1'b0}), .a ({signal_1400, signal_1115}), .clk (clk), .r (Fresh[199]), .c ({signal_1532, signal_1205}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1019 ( .s ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({signal_1264, signal_1043}), .a ({signal_1398, signal_1113}), .clk (clk), .r (Fresh[200]), .c ({signal_1533, signal_1206}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1020 ( .s ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({signal_1396, signal_1111}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[201]), .c ({signal_1534, signal_1207}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1021 ( .s ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({signal_1396, signal_1111}), .a ({signal_1264, signal_1043}), .clk (clk), .r (Fresh[202]), .c ({signal_1535, signal_1208}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1022 ( .s ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({signal_1403, signal_1117}), .a ({signal_1402, signal_1116}), .clk (clk), .r (Fresh[203]), .c ({signal_1537, signal_1209}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1023 ( .s ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({1'b0, 1'b0}), .a ({signal_1402, signal_1116}), .clk (clk), .r (Fresh[204]), .c ({signal_1538, signal_1210}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1024 ( .s ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_1405, signal_1119}), .a ({signal_1404, signal_1118}), .clk (clk), .r (Fresh[205]), .c ({signal_1540, signal_721}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1025 ( .s ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({1'b0, 1'b0}), .a ({signal_1406, signal_1120}), .clk (clk), .r (Fresh[206]), .c ({signal_1541, signal_1211}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1026 ( .s ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({signal_1267, signal_1045}), .a ({signal_1404, signal_1118}), .clk (clk), .r (Fresh[207]), .c ({signal_1542, signal_1212}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1027 ( .s ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({signal_1402, signal_1116}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[208]), .c ({signal_1543, signal_1213}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1028 ( .s ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({signal_1402, signal_1116}), .a ({signal_1267, signal_1045}), .clk (clk), .r (Fresh[209]), .c ({signal_1544, signal_1214}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1029 ( .s ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({signal_1409, signal_1122}), .a ({signal_1408, signal_1121}), .clk (clk), .r (Fresh[210]), .c ({signal_1546, signal_1215}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1030 ( .s ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({1'b0, 1'b0}), .a ({signal_1408, signal_1121}), .clk (clk), .r (Fresh[211]), .c ({signal_1547, signal_1216}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1031 ( .s ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_1411, signal_1124}), .a ({signal_1410, signal_1123}), .clk (clk), .r (Fresh[212]), .c ({signal_1549, signal_717}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1032 ( .s ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({1'b0, 1'b0}), .a ({signal_1412, signal_1125}), .clk (clk), .r (Fresh[213]), .c ({signal_1550, signal_1217}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1033 ( .s ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({signal_1270, signal_1047}), .a ({signal_1410, signal_1123}), .clk (clk), .r (Fresh[214]), .c ({signal_1551, signal_1218}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1034 ( .s ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({signal_1408, signal_1121}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[215]), .c ({signal_1552, signal_1219}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1035 ( .s ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({signal_1408, signal_1121}), .a ({signal_1270, signal_1047}), .clk (clk), .r (Fresh[216]), .c ({signal_1553, signal_1220}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1036 ( .s ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({signal_1415, signal_1127}), .a ({signal_1414, signal_1126}), .clk (clk), .r (Fresh[217]), .c ({signal_1555, signal_1221}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1037 ( .s ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({1'b0, 1'b0}), .a ({signal_1414, signal_1126}), .clk (clk), .r (Fresh[218]), .c ({signal_1556, signal_1222}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1038 ( .s ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_1417, signal_1129}), .a ({signal_1416, signal_1128}), .clk (clk), .r (Fresh[219]), .c ({signal_1558, signal_713}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1039 ( .s ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({1'b0, 1'b0}), .a ({signal_1418, signal_1130}), .clk (clk), .r (Fresh[220]), .c ({signal_1559, signal_1223}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1040 ( .s ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({signal_1273, signal_1049}), .a ({signal_1416, signal_1128}), .clk (clk), .r (Fresh[221]), .c ({signal_1560, signal_1224}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1041 ( .s ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({signal_1414, signal_1126}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[222]), .c ({signal_1561, signal_1225}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1042 ( .s ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({signal_1414, signal_1126}), .a ({signal_1273, signal_1049}), .clk (clk), .r (Fresh[223]), .c ({signal_1562, signal_1226}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_0 ( .s (rst), .b ({signal_1739, signal_774}), .a ({plaintext_s1[0], plaintext_s0[0]}), .c ({signal_1788, signal_870}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2 ( .s (rst), .b ({signal_1740, signal_772}), .a ({plaintext_s1[2], plaintext_s0[2]}), .c ({signal_1790, signal_868}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3 ( .s (rst), .b ({signal_1741, signal_771}), .a ({plaintext_s1[3], plaintext_s0[3]}), .c ({signal_1792, signal_867}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_4 ( .s (rst), .b ({signal_1742, signal_770}), .a ({plaintext_s1[4], plaintext_s0[4]}), .c ({signal_1794, signal_866}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_6 ( .s (rst), .b ({signal_1743, signal_768}), .a ({plaintext_s1[6], plaintext_s0[6]}), .c ({signal_1796, signal_864}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_7 ( .s (rst), .b ({signal_1744, signal_767}), .a ({plaintext_s1[7], plaintext_s0[7]}), .c ({signal_1798, signal_863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_8 ( .s (rst), .b ({signal_1745, signal_766}), .a ({plaintext_s1[8], plaintext_s0[8]}), .c ({signal_1800, signal_862}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_10 ( .s (rst), .b ({signal_1746, signal_764}), .a ({plaintext_s1[10], plaintext_s0[10]}), .c ({signal_1802, signal_860}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_11 ( .s (rst), .b ({signal_1747, signal_763}), .a ({plaintext_s1[11], plaintext_s0[11]}), .c ({signal_1804, signal_859}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_12 ( .s (rst), .b ({signal_1748, signal_762}), .a ({plaintext_s1[12], plaintext_s0[12]}), .c ({signal_1806, signal_858}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_14 ( .s (rst), .b ({signal_1749, signal_760}), .a ({plaintext_s1[14], plaintext_s0[14]}), .c ({signal_1808, signal_856}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_15 ( .s (rst), .b ({signal_1750, signal_759}), .a ({plaintext_s1[15], plaintext_s0[15]}), .c ({signal_1810, signal_855}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_16 ( .s (rst), .b ({signal_1751, signal_758}), .a ({plaintext_s1[16], plaintext_s0[16]}), .c ({signal_1812, signal_854}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_18 ( .s (rst), .b ({signal_1752, signal_756}), .a ({plaintext_s1[18], plaintext_s0[18]}), .c ({signal_1814, signal_852}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_19 ( .s (rst), .b ({signal_1753, signal_755}), .a ({plaintext_s1[19], plaintext_s0[19]}), .c ({signal_1816, signal_851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_20 ( .s (rst), .b ({signal_1754, signal_754}), .a ({plaintext_s1[20], plaintext_s0[20]}), .c ({signal_1818, signal_850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_22 ( .s (rst), .b ({signal_1755, signal_752}), .a ({plaintext_s1[22], plaintext_s0[22]}), .c ({signal_1820, signal_848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_23 ( .s (rst), .b ({signal_1756, signal_751}), .a ({plaintext_s1[23], plaintext_s0[23]}), .c ({signal_1822, signal_847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_24 ( .s (rst), .b ({signal_1757, signal_750}), .a ({plaintext_s1[24], plaintext_s0[24]}), .c ({signal_1824, signal_846}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_26 ( .s (rst), .b ({signal_1758, signal_748}), .a ({plaintext_s1[26], plaintext_s0[26]}), .c ({signal_1826, signal_844}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_27 ( .s (rst), .b ({signal_1759, signal_747}), .a ({plaintext_s1[27], plaintext_s0[27]}), .c ({signal_1828, signal_843}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_28 ( .s (rst), .b ({signal_1760, signal_746}), .a ({plaintext_s1[28], plaintext_s0[28]}), .c ({signal_1830, signal_842}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_30 ( .s (rst), .b ({signal_1761, signal_744}), .a ({plaintext_s1[30], plaintext_s0[30]}), .c ({signal_1832, signal_840}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_31 ( .s (rst), .b ({signal_1762, signal_743}), .a ({plaintext_s1[31], plaintext_s0[31]}), .c ({signal_1834, signal_839}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_32 ( .s (rst), .b ({signal_1763, signal_742}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({signal_1836, signal_806}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_34 ( .s (rst), .b ({signal_1764, signal_740}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({signal_1838, signal_804}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_35 ( .s (rst), .b ({signal_1765, signal_739}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({signal_1840, signal_803}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_36 ( .s (rst), .b ({signal_1766, signal_738}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({signal_1842, signal_802}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_38 ( .s (rst), .b ({signal_1767, signal_736}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({signal_1844, signal_800}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_39 ( .s (rst), .b ({signal_1768, signal_735}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({signal_1846, signal_799}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_40 ( .s (rst), .b ({signal_1769, signal_734}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({signal_1848, signal_798}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_42 ( .s (rst), .b ({signal_1770, signal_732}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({signal_1850, signal_796}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_43 ( .s (rst), .b ({signal_1771, signal_731}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({signal_1852, signal_795}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_44 ( .s (rst), .b ({signal_1772, signal_730}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({signal_1854, signal_794}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_46 ( .s (rst), .b ({signal_1773, signal_728}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({signal_1856, signal_792}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_47 ( .s (rst), .b ({signal_1774, signal_727}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({signal_1858, signal_791}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_48 ( .s (rst), .b ({signal_1775, signal_726}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({signal_1860, signal_790}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_50 ( .s (rst), .b ({signal_1776, signal_724}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({signal_1862, signal_788}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_51 ( .s (rst), .b ({signal_1777, signal_723}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({signal_1864, signal_787}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_52 ( .s (rst), .b ({signal_1778, signal_722}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({signal_1866, signal_786}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_54 ( .s (rst), .b ({signal_1779, signal_720}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({signal_1868, signal_784}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_55 ( .s (rst), .b ({signal_1780, signal_719}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({signal_1870, signal_783}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_56 ( .s (rst), .b ({signal_1781, signal_718}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({signal_1872, signal_782}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_58 ( .s (rst), .b ({signal_1782, signal_716}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({signal_1874, signal_780}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_59 ( .s (rst), .b ({signal_1783, signal_715}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({signal_1876, signal_779}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_60 ( .s (rst), .b ({signal_1784, signal_714}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({signal_1878, signal_778}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_62 ( .s (rst), .b ({signal_1785, signal_712}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({signal_1880, signal_776}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_63 ( .s (rst), .b ({signal_1786, signal_711}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({signal_1882, signal_775}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_64 ( .a ({signal_1912, signal_268}), .b ({signal_1911, signal_269}), .c ({signal_1987, signal_822}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_65 ( .a ({signal_1812, signal_854}), .b ({signal_1788, signal_870}), .c ({signal_1911, signal_269}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_66 ( .a ({1'b0, 1'b0}), .b ({signal_1860, signal_790}), .c ({signal_1912, signal_268}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_67 ( .a ({signal_1913, signal_270}), .b ({signal_1788, signal_870}), .c ({signal_1988, signal_838}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_68 ( .a ({1'b0, 1'b0}), .b ({signal_1836, signal_806}), .c ({signal_1913, signal_270}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_74 ( .a ({signal_1917, signal_274}), .b ({signal_1916, signal_275}), .c ({signal_1989, signal_820}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_75 ( .a ({signal_1814, signal_852}), .b ({signal_1790, signal_868}), .c ({signal_1916, signal_275}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_76 ( .a ({1'b0, 1'b0}), .b ({signal_1862, signal_788}), .c ({signal_1917, signal_274}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_77 ( .a ({signal_1918, signal_276}), .b ({signal_1790, signal_868}), .c ({signal_1990, signal_836}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_78 ( .a ({1'b0, 1'b0}), .b ({signal_1838, signal_804}), .c ({signal_1918, signal_276}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_79 ( .a ({signal_1920, signal_277}), .b ({signal_1919, signal_278}), .c ({signal_1991, signal_819}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_80 ( .a ({signal_1816, signal_851}), .b ({signal_1792, signal_867}), .c ({signal_1919, signal_278}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_81 ( .a ({1'b0, 1'b0}), .b ({signal_1864, signal_787}), .c ({signal_1920, signal_277}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_82 ( .a ({signal_1921, signal_279}), .b ({signal_1792, signal_867}), .c ({signal_1992, signal_835}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_83 ( .a ({1'b0, 1'b0}), .b ({signal_1840, signal_803}), .c ({signal_1921, signal_279}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_84 ( .a ({signal_1923, signal_280}), .b ({signal_1922, signal_281}), .c ({signal_1993, signal_818}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_85 ( .a ({signal_1818, signal_850}), .b ({signal_1794, signal_866}), .c ({signal_1922, signal_281}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_86 ( .a ({1'b0, 1'b0}), .b ({signal_1866, signal_786}), .c ({signal_1923, signal_280}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_87 ( .a ({signal_1924, signal_282}), .b ({signal_1794, signal_866}), .c ({signal_1994, signal_834}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_88 ( .a ({1'b0, 1'b0}), .b ({signal_1842, signal_802}), .c ({signal_1924, signal_282}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_94 ( .a ({signal_1928, signal_286}), .b ({signal_1927, signal_287}), .c ({signal_1995, signal_816}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_95 ( .a ({signal_1820, signal_848}), .b ({signal_1796, signal_864}), .c ({signal_1927, signal_287}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_96 ( .a ({1'b0, 1'b0}), .b ({signal_1868, signal_784}), .c ({signal_1928, signal_286}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_97 ( .a ({signal_1929, signal_288}), .b ({signal_1796, signal_864}), .c ({signal_1996, signal_832}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_98 ( .a ({1'b0, 1'b0}), .b ({signal_1844, signal_800}), .c ({signal_1929, signal_288}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_99 ( .a ({signal_1931, signal_289}), .b ({signal_1930, signal_290}), .c ({signal_1997, signal_815}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_100 ( .a ({signal_1822, signal_847}), .b ({signal_1798, signal_863}), .c ({signal_1930, signal_290}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_101 ( .a ({1'b0, 1'b0}), .b ({signal_1870, signal_783}), .c ({signal_1931, signal_289}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_102 ( .a ({signal_1932, signal_291}), .b ({signal_1798, signal_863}), .c ({signal_1998, signal_831}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_103 ( .a ({1'b0, 1'b0}), .b ({signal_1846, signal_799}), .c ({signal_1932, signal_291}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_104 ( .a ({signal_1934, signal_292}), .b ({signal_1933, signal_293}), .c ({signal_1999, signal_814}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_105 ( .a ({signal_1824, signal_846}), .b ({signal_1800, signal_862}), .c ({signal_1933, signal_293}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_106 ( .a ({1'b0, 1'b0}), .b ({signal_1872, signal_782}), .c ({signal_1934, signal_292}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_107 ( .a ({signal_1935, signal_294}), .b ({signal_1800, signal_862}), .c ({signal_2000, signal_830}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_108 ( .a ({1'b0, 1'b0}), .b ({signal_1848, signal_798}), .c ({signal_1935, signal_294}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_114 ( .a ({signal_1939, signal_298}), .b ({signal_1938, signal_299}), .c ({signal_2001, signal_812}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_115 ( .a ({signal_1826, signal_844}), .b ({signal_1802, signal_860}), .c ({signal_1938, signal_299}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_116 ( .a ({1'b0, 1'b0}), .b ({signal_1874, signal_780}), .c ({signal_1939, signal_298}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_117 ( .a ({signal_1940, signal_300}), .b ({signal_1802, signal_860}), .c ({signal_2002, signal_828}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_118 ( .a ({1'b0, 1'b0}), .b ({signal_1850, signal_796}), .c ({signal_1940, signal_300}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_119 ( .a ({signal_1942, signal_301}), .b ({signal_1941, signal_302}), .c ({signal_2003, signal_811}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_120 ( .a ({signal_1828, signal_843}), .b ({signal_1804, signal_859}), .c ({signal_1941, signal_302}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_121 ( .a ({1'b0, 1'b0}), .b ({signal_1876, signal_779}), .c ({signal_1942, signal_301}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_122 ( .a ({signal_1943, signal_303}), .b ({signal_1804, signal_859}), .c ({signal_2004, signal_827}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_123 ( .a ({1'b0, 1'b0}), .b ({signal_1852, signal_795}), .c ({signal_1943, signal_303}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_124 ( .a ({signal_1945, signal_304}), .b ({signal_1944, signal_305}), .c ({signal_2005, signal_810}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_125 ( .a ({signal_1830, signal_842}), .b ({signal_1806, signal_858}), .c ({signal_1944, signal_305}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_126 ( .a ({1'b0, 1'b0}), .b ({signal_1878, signal_778}), .c ({signal_1945, signal_304}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_127 ( .a ({signal_1946, signal_306}), .b ({signal_1806, signal_858}), .c ({signal_2006, signal_826}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_128 ( .a ({1'b0, 1'b0}), .b ({signal_1854, signal_794}), .c ({signal_1946, signal_306}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_134 ( .a ({signal_1950, signal_310}), .b ({signal_1949, signal_311}), .c ({signal_2007, signal_808}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_135 ( .a ({signal_1832, signal_840}), .b ({signal_1808, signal_856}), .c ({signal_1949, signal_311}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_136 ( .a ({1'b0, 1'b0}), .b ({signal_1880, signal_776}), .c ({signal_1950, signal_310}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_137 ( .a ({signal_1951, signal_312}), .b ({signal_1808, signal_856}), .c ({signal_2008, signal_824}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_138 ( .a ({1'b0, 1'b0}), .b ({signal_1856, signal_792}), .c ({signal_1951, signal_312}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_139 ( .a ({signal_1953, signal_313}), .b ({signal_1952, signal_314}), .c ({signal_2009, signal_807}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_140 ( .a ({signal_1834, signal_839}), .b ({signal_1810, signal_855}), .c ({signal_1952, signal_314}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_141 ( .a ({1'b0, 1'b0}), .b ({signal_1882, signal_775}), .c ({signal_1953, signal_313}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_142 ( .a ({signal_1954, signal_315}), .b ({signal_1810, signal_855}), .c ({signal_2010, signal_823}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_143 ( .a ({1'b0, 1'b0}), .b ({signal_1858, signal_791}), .c ({signal_1954, signal_315}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_144 ( .a ({signal_2043, signal_316}), .b ({signal_1708, signal_886}), .c ({signal_2075, signal_950}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_145 ( .a ({1'b0, 1'b0}), .b ({signal_1987, signal_822}), .c ({signal_2043, signal_316}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_148 ( .a ({signal_2045, signal_318}), .b ({signal_1714, signal_884}), .c ({signal_2076, signal_948}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_149 ( .a ({1'b0, 1'b0}), .b ({signal_1989, signal_820}), .c ({signal_2045, signal_318}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_150 ( .a ({signal_2046, signal_319}), .b ({signal_1717, signal_883}), .c ({signal_2077, signal_947}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_151 ( .a ({1'b0, 1'b0}), .b ({signal_1991, signal_819}), .c ({signal_2046, signal_319}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_152 ( .a ({signal_2047, signal_320}), .b ({signal_1720, signal_882}), .c ({signal_2078, signal_946}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_153 ( .a ({1'b0, 1'b0}), .b ({signal_1993, signal_818}), .c ({signal_2047, signal_320}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_156 ( .a ({signal_2049, signal_322}), .b ({signal_1313, signal_880}), .c ({signal_2079, signal_944}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_157 ( .a ({1'b0, 1'b0}), .b ({signal_1995, signal_816}), .c ({signal_2049, signal_322}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_158 ( .a ({signal_2050, signal_323}), .b ({signal_1723, signal_879}), .c ({signal_2080, signal_943}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_159 ( .a ({1'b0, 1'b0}), .b ({signal_1997, signal_815}), .c ({signal_2050, signal_323}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_160 ( .a ({signal_2051, signal_324}), .b ({signal_1316, signal_878}), .c ({signal_2081, signal_942}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_161 ( .a ({1'b0, 1'b0}), .b ({signal_1999, signal_814}), .c ({signal_2051, signal_324}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_164 ( .a ({signal_2053, signal_326}), .b ({signal_1729, signal_876}), .c ({signal_2082, signal_940}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_165 ( .a ({1'b0, 1'b0}), .b ({signal_2001, signal_812}), .c ({signal_2053, signal_326}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_166 ( .a ({signal_2054, signal_327}), .b ({signal_1319, signal_875}), .c ({signal_2083, signal_939}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_167 ( .a ({1'b0, 1'b0}), .b ({signal_2003, signal_811}), .c ({signal_2054, signal_327}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_168 ( .a ({signal_2055, signal_328}), .b ({signal_1732, signal_874}), .c ({signal_2084, signal_938}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_169 ( .a ({1'b0, 1'b0}), .b ({signal_2005, signal_810}), .c ({signal_2055, signal_328}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_172 ( .a ({signal_2057, signal_330}), .b ({signal_1322, signal_872}), .c ({signal_2085, signal_936}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_173 ( .a ({1'b0, 1'b0}), .b ({signal_2007, signal_808}), .c ({signal_2057, signal_330}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_174 ( .a ({signal_2058, signal_331}), .b ({signal_1738, signal_871}), .c ({signal_2086, signal_935}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_175 ( .a ({1'b0, 1'b0}), .b ({signal_2009, signal_807}), .c ({signal_2058, signal_331}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_176 ( .a ({signal_2059, signal_332}), .b ({signal_1895, signal_333}), .c ({signal_2087, signal_958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_178 ( .a ({1'b0, 1'b0}), .b ({signal_2000, signal_830}), .c ({signal_2059, signal_332}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_182 ( .a ({signal_2061, signal_336}), .b ({signal_1897, signal_337}), .c ({signal_2088, signal_956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_184 ( .a ({1'b0, 1'b0}), .b ({signal_2002, signal_828}), .c ({signal_2061, signal_336}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_185 ( .a ({signal_2062, signal_338}), .b ({signal_1898, signal_339}), .c ({signal_2089, signal_955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_187 ( .a ({1'b0, 1'b0}), .b ({signal_2004, signal_827}), .c ({signal_2062, signal_338}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_188 ( .a ({signal_2063, signal_340}), .b ({signal_1899, signal_341}), .c ({signal_2090, signal_954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_190 ( .a ({1'b0, 1'b0}), .b ({signal_2006, signal_826}), .c ({signal_2063, signal_340}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_194 ( .a ({signal_2065, signal_344}), .b ({signal_1901, signal_345}), .c ({signal_2091, signal_952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_196 ( .a ({1'b0, 1'b0}), .b ({signal_2008, signal_824}), .c ({signal_2065, signal_344}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_197 ( .a ({signal_2066, signal_346}), .b ({signal_1902, signal_347}), .c ({signal_2092, signal_951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_199 ( .a ({1'b0, 1'b0}), .b ({signal_2010, signal_823}), .c ({signal_2066, signal_346}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_200 ( .a ({signal_1955, signal_348}), .b ({signal_1277, signal_934}), .c ({signal_2017, signal_998}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_201 ( .a ({1'b0, 1'b0}), .b ({signal_1788, signal_870}), .c ({signal_1955, signal_348}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_204 ( .a ({signal_1957, signal_350}), .b ({signal_1280, signal_932}), .c ({signal_2018, signal_996}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_205 ( .a ({1'b0, 1'b0}), .b ({signal_1790, signal_868}), .c ({signal_1957, signal_350}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_206 ( .a ({signal_1958, signal_351}), .b ({signal_1600, signal_931}), .c ({signal_2019, signal_995}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_207 ( .a ({1'b0, 1'b0}), .b ({signal_1792, signal_867}), .c ({signal_1958, signal_351}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_208 ( .a ({signal_1959, signal_352}), .b ({signal_1603, signal_930}), .c ({signal_2020, signal_994}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_209 ( .a ({1'b0, 1'b0}), .b ({signal_1794, signal_866}), .c ({signal_1959, signal_352}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_212 ( .a ({signal_1961, signal_354}), .b ({signal_1609, signal_928}), .c ({signal_2021, signal_992}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_213 ( .a ({1'b0, 1'b0}), .b ({signal_1796, signal_864}), .c ({signal_1961, signal_354}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_214 ( .a ({signal_1962, signal_355}), .b ({signal_1612, signal_927}), .c ({signal_2022, signal_991}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_215 ( .a ({1'b0, 1'b0}), .b ({signal_1798, signal_863}), .c ({signal_1962, signal_355}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_216 ( .a ({signal_1963, signal_356}), .b ({signal_1615, signal_926}), .c ({signal_2023, signal_990}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_217 ( .a ({1'b0, 1'b0}), .b ({signal_1800, signal_862}), .c ({signal_1963, signal_356}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_220 ( .a ({signal_1965, signal_358}), .b ({signal_1621, signal_924}), .c ({signal_2024, signal_988}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_221 ( .a ({1'b0, 1'b0}), .b ({signal_1802, signal_860}), .c ({signal_1965, signal_358}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_222 ( .a ({signal_1966, signal_359}), .b ({signal_1624, signal_923}), .c ({signal_2025, signal_987}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_223 ( .a ({1'b0, 1'b0}), .b ({signal_1804, signal_859}), .c ({signal_1966, signal_359}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_224 ( .a ({signal_1967, signal_360}), .b ({signal_1627, signal_922}), .c ({signal_2026, signal_986}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_225 ( .a ({1'b0, 1'b0}), .b ({signal_1806, signal_858}), .c ({signal_1967, signal_360}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_228 ( .a ({signal_1969, signal_362}), .b ({signal_1633, signal_920}), .c ({signal_2027, signal_984}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_229 ( .a ({1'b0, 1'b0}), .b ({signal_1808, signal_856}), .c ({signal_1969, signal_362}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_230 ( .a ({signal_1970, signal_363}), .b ({signal_1636, signal_919}), .c ({signal_2028, signal_983}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_231 ( .a ({1'b0, 1'b0}), .b ({signal_1810, signal_855}), .c ({signal_1970, signal_363}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_232 ( .a ({signal_1971, signal_364}), .b ({signal_1639, signal_918}), .c ({signal_2029, signal_982}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_233 ( .a ({1'b0, 1'b0}), .b ({signal_1812, signal_854}), .c ({signal_1971, signal_364}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_236 ( .a ({signal_1973, signal_366}), .b ({signal_1645, signal_916}), .c ({signal_2030, signal_980}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_237 ( .a ({1'b0, 1'b0}), .b ({signal_1814, signal_852}), .c ({signal_1973, signal_366}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_238 ( .a ({signal_1974, signal_367}), .b ({signal_1648, signal_915}), .c ({signal_2031, signal_979}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_239 ( .a ({1'b0, 1'b0}), .b ({signal_1816, signal_851}), .c ({signal_1974, signal_367}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_240 ( .a ({signal_1975, signal_368}), .b ({signal_1651, signal_914}), .c ({signal_2032, signal_978}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_241 ( .a ({1'b0, 1'b0}), .b ({signal_1818, signal_850}), .c ({signal_1975, signal_368}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_244 ( .a ({signal_1977, signal_370}), .b ({signal_1283, signal_912}), .c ({signal_2033, signal_976}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_245 ( .a ({1'b0, 1'b0}), .b ({signal_1820, signal_848}), .c ({signal_1977, signal_370}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_246 ( .a ({signal_1978, signal_371}), .b ({signal_1286, signal_911}), .c ({signal_2034, signal_975}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_247 ( .a ({1'b0, 1'b0}), .b ({signal_1822, signal_847}), .c ({signal_1978, signal_371}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_248 ( .a ({signal_1979, signal_372}), .b ({signal_1289, signal_910}), .c ({signal_2035, signal_974}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_249 ( .a ({1'b0, 1'b0}), .b ({signal_1824, signal_846}), .c ({signal_1979, signal_372}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_252 ( .a ({signal_1981, signal_374}), .b ({signal_1295, signal_908}), .c ({signal_2036, signal_972}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_253 ( .a ({1'b0, 1'b0}), .b ({signal_1826, signal_844}), .c ({signal_1981, signal_374}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_254 ( .a ({signal_1982, signal_375}), .b ({signal_1298, signal_907}), .c ({signal_2037, signal_971}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_255 ( .a ({1'b0, 1'b0}), .b ({signal_1828, signal_843}), .c ({signal_1982, signal_375}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_256 ( .a ({signal_1983, signal_376}), .b ({signal_1657, signal_906}), .c ({signal_2038, signal_970}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_257 ( .a ({1'b0, 1'b0}), .b ({signal_1830, signal_842}), .c ({signal_1983, signal_376}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_260 ( .a ({signal_1985, signal_378}), .b ({signal_1663, signal_904}), .c ({signal_2039, signal_968}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_261 ( .a ({1'b0, 1'b0}), .b ({signal_1832, signal_840}), .c ({signal_1985, signal_378}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_262 ( .a ({signal_1986, signal_379}), .b ({signal_1666, signal_903}), .c ({signal_2040, signal_967}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_263 ( .a ({1'b0, 1'b0}), .b ({signal_1834, signal_839}), .c ({signal_1986, signal_379}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_264 ( .a ({signal_2067, signal_380}), .b ({signal_1669, signal_902}), .c ({signal_2093, signal_966}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_265 ( .a ({1'b0, 1'b0}), .b ({signal_1988, signal_838}), .c ({signal_2067, signal_380}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_268 ( .a ({signal_2069, signal_382}), .b ({signal_1672, signal_900}), .c ({signal_2094, signal_964}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_269 ( .a ({1'b0, 1'b0}), .b ({signal_1990, signal_836}), .c ({signal_2069, signal_382}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_270 ( .a ({signal_2070, signal_383}), .b ({signal_1675, signal_899}), .c ({signal_2095, signal_963}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_271 ( .a ({1'b0, 1'b0}), .b ({signal_1992, signal_835}), .c ({signal_2070, signal_383}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_272 ( .a ({signal_2071, signal_384}), .b ({signal_1304, signal_898}), .c ({signal_2096, signal_962}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_273 ( .a ({1'b0, 1'b0}), .b ({signal_1994, signal_834}), .c ({signal_2071, signal_384}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_276 ( .a ({signal_2073, signal_386}), .b ({signal_1681, signal_896}), .c ({signal_2097, signal_960}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_277 ( .a ({1'b0, 1'b0}), .b ({signal_1996, signal_832}), .c ({signal_2073, signal_386}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_278 ( .a ({signal_2074, signal_387}), .b ({signal_1307, signal_895}), .c ({signal_2098, signal_959}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_279 ( .a ({1'b0, 1'b0}), .b ({signal_1998, signal_831}), .c ({signal_2074, signal_387}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1043 ( .s ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_1421, signal_1132}), .a ({signal_1420, signal_1131}), .clk (clk), .r (Fresh[224]), .c ({signal_1739, signal_774}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1044 ( .s ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_1425, signal_1134}), .a ({signal_1424, signal_1133}), .clk (clk), .r (Fresh[225]), .c ({signal_1740, signal_772}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1045 ( .s ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_1427, signal_1136}), .a ({signal_1426, signal_1135}), .clk (clk), .r (Fresh[226]), .c ({signal_1741, signal_771}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1046 ( .s ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_1430, signal_1138}), .a ({signal_1429, signal_1137}), .clk (clk), .r (Fresh[227]), .c ({signal_1742, signal_770}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1047 ( .s ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_1434, signal_1140}), .a ({signal_1433, signal_1139}), .clk (clk), .r (Fresh[228]), .c ({signal_1743, signal_768}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1048 ( .s ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_1436, signal_1142}), .a ({signal_1435, signal_1141}), .clk (clk), .r (Fresh[229]), .c ({signal_1744, signal_767}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1049 ( .s ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_1439, signal_1144}), .a ({signal_1438, signal_1143}), .clk (clk), .r (Fresh[230]), .c ({signal_1745, signal_766}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1050 ( .s ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_1443, signal_1146}), .a ({signal_1442, signal_1145}), .clk (clk), .r (Fresh[231]), .c ({signal_1746, signal_764}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1051 ( .s ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_1445, signal_1148}), .a ({signal_1444, signal_1147}), .clk (clk), .r (Fresh[232]), .c ({signal_1747, signal_763}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1052 ( .s ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_1448, signal_1150}), .a ({signal_1447, signal_1149}), .clk (clk), .r (Fresh[233]), .c ({signal_1748, signal_762}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1053 ( .s ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_1452, signal_1152}), .a ({signal_1451, signal_1151}), .clk (clk), .r (Fresh[234]), .c ({signal_1749, signal_760}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1054 ( .s ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_1454, signal_1154}), .a ({signal_1453, signal_1153}), .clk (clk), .r (Fresh[235]), .c ({signal_1750, signal_759}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1055 ( .s ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_1457, signal_1156}), .a ({signal_1456, signal_1155}), .clk (clk), .r (Fresh[236]), .c ({signal_1751, signal_758}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1056 ( .s ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_1461, signal_1158}), .a ({signal_1460, signal_1157}), .clk (clk), .r (Fresh[237]), .c ({signal_1752, signal_756}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1057 ( .s ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_1463, signal_1160}), .a ({signal_1462, signal_1159}), .clk (clk), .r (Fresh[238]), .c ({signal_1753, signal_755}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1058 ( .s ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_1466, signal_1162}), .a ({signal_1465, signal_1161}), .clk (clk), .r (Fresh[239]), .c ({signal_1754, signal_754}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1059 ( .s ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_1470, signal_1164}), .a ({signal_1469, signal_1163}), .clk (clk), .r (Fresh[240]), .c ({signal_1755, signal_752}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1060 ( .s ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_1472, signal_1166}), .a ({signal_1471, signal_1165}), .clk (clk), .r (Fresh[241]), .c ({signal_1756, signal_751}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1061 ( .s ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_1475, signal_1168}), .a ({signal_1474, signal_1167}), .clk (clk), .r (Fresh[242]), .c ({signal_1757, signal_750}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1062 ( .s ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_1479, signal_1170}), .a ({signal_1478, signal_1169}), .clk (clk), .r (Fresh[243]), .c ({signal_1758, signal_748}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1063 ( .s ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_1481, signal_1172}), .a ({signal_1480, signal_1171}), .clk (clk), .r (Fresh[244]), .c ({signal_1759, signal_747}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1064 ( .s ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_1484, signal_1174}), .a ({signal_1483, signal_1173}), .clk (clk), .r (Fresh[245]), .c ({signal_1760, signal_746}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1065 ( .s ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_1488, signal_1176}), .a ({signal_1487, signal_1175}), .clk (clk), .r (Fresh[246]), .c ({signal_1761, signal_744}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1066 ( .s ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_1490, signal_1178}), .a ({signal_1489, signal_1177}), .clk (clk), .r (Fresh[247]), .c ({signal_1762, signal_743}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1067 ( .s ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_1493, signal_1180}), .a ({signal_1492, signal_1179}), .clk (clk), .r (Fresh[248]), .c ({signal_1763, signal_742}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1068 ( .s ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_1497, signal_1182}), .a ({signal_1496, signal_1181}), .clk (clk), .r (Fresh[249]), .c ({signal_1764, signal_740}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1069 ( .s ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_1499, signal_1184}), .a ({signal_1498, signal_1183}), .clk (clk), .r (Fresh[250]), .c ({signal_1765, signal_739}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1070 ( .s ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_1502, signal_1186}), .a ({signal_1501, signal_1185}), .clk (clk), .r (Fresh[251]), .c ({signal_1766, signal_738}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1071 ( .s ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_1506, signal_1188}), .a ({signal_1505, signal_1187}), .clk (clk), .r (Fresh[252]), .c ({signal_1767, signal_736}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1072 ( .s ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_1508, signal_1190}), .a ({signal_1507, signal_1189}), .clk (clk), .r (Fresh[253]), .c ({signal_1768, signal_735}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1073 ( .s ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_1511, signal_1192}), .a ({signal_1510, signal_1191}), .clk (clk), .r (Fresh[254]), .c ({signal_1769, signal_734}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1074 ( .s ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_1515, signal_1194}), .a ({signal_1514, signal_1193}), .clk (clk), .r (Fresh[255]), .c ({signal_1770, signal_732}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1075 ( .s ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_1517, signal_1196}), .a ({signal_1516, signal_1195}), .clk (clk), .r (Fresh[256]), .c ({signal_1771, signal_731}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1076 ( .s ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_1520, signal_1198}), .a ({signal_1519, signal_1197}), .clk (clk), .r (Fresh[257]), .c ({signal_1772, signal_730}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1077 ( .s ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_1524, signal_1200}), .a ({signal_1523, signal_1199}), .clk (clk), .r (Fresh[258]), .c ({signal_1773, signal_728}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1078 ( .s ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_1526, signal_1202}), .a ({signal_1525, signal_1201}), .clk (clk), .r (Fresh[259]), .c ({signal_1774, signal_727}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1079 ( .s ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_1529, signal_1204}), .a ({signal_1528, signal_1203}), .clk (clk), .r (Fresh[260]), .c ({signal_1775, signal_726}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1080 ( .s ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_1533, signal_1206}), .a ({signal_1532, signal_1205}), .clk (clk), .r (Fresh[261]), .c ({signal_1776, signal_724}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1081 ( .s ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_1535, signal_1208}), .a ({signal_1534, signal_1207}), .clk (clk), .r (Fresh[262]), .c ({signal_1777, signal_723}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1082 ( .s ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_1538, signal_1210}), .a ({signal_1537, signal_1209}), .clk (clk), .r (Fresh[263]), .c ({signal_1778, signal_722}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1083 ( .s ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_1542, signal_1212}), .a ({signal_1541, signal_1211}), .clk (clk), .r (Fresh[264]), .c ({signal_1779, signal_720}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1084 ( .s ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_1544, signal_1214}), .a ({signal_1543, signal_1213}), .clk (clk), .r (Fresh[265]), .c ({signal_1780, signal_719}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1085 ( .s ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_1547, signal_1216}), .a ({signal_1546, signal_1215}), .clk (clk), .r (Fresh[266]), .c ({signal_1781, signal_718}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1086 ( .s ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_1551, signal_1218}), .a ({signal_1550, signal_1217}), .clk (clk), .r (Fresh[267]), .c ({signal_1782, signal_716}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1087 ( .s ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_1553, signal_1220}), .a ({signal_1552, signal_1219}), .clk (clk), .r (Fresh[268]), .c ({signal_1783, signal_715}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1088 ( .s ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_1556, signal_1222}), .a ({signal_1555, signal_1221}), .clk (clk), .r (Fresh[269]), .c ({signal_1784, signal_714}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1089 ( .s ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_1560, signal_1224}), .a ({signal_1559, signal_1223}), .clk (clk), .r (Fresh[270]), .c ({signal_1785, signal_712}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1090 ( .s ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_1562, signal_1226}), .a ({signal_1561, signal_1225}), .clk (clk), .r (Fresh[271]), .c ({signal_1786, signal_711}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) cell_281 ( .clk (signal_2371), .D ({signal_2086, signal_935}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_283 ( .clk (signal_2371), .D ({signal_2085, signal_936}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_285 ( .clk (signal_2371), .D ({signal_2056, signal_937}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_287 ( .clk (signal_2371), .D ({signal_2084, signal_938}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_289 ( .clk (signal_2371), .D ({signal_2083, signal_939}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_291 ( .clk (signal_2371), .D ({signal_2082, signal_940}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_293 ( .clk (signal_2371), .D ({signal_2052, signal_941}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_295 ( .clk (signal_2371), .D ({signal_2081, signal_942}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_297 ( .clk (signal_2371), .D ({signal_2080, signal_943}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_299 ( .clk (signal_2371), .D ({signal_2079, signal_944}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_301 ( .clk (signal_2371), .D ({signal_2048, signal_945}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_303 ( .clk (signal_2371), .D ({signal_2078, signal_946}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_305 ( .clk (signal_2371), .D ({signal_2077, signal_947}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_307 ( .clk (signal_2371), .D ({signal_2076, signal_948}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_309 ( .clk (signal_2371), .D ({signal_2044, signal_949}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_311 ( .clk (signal_2371), .D ({signal_2075, signal_950}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_313 ( .clk (signal_2371), .D ({signal_2092, signal_951}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_315 ( .clk (signal_2371), .D ({signal_2091, signal_952}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_317 ( .clk (signal_2371), .D ({signal_2064, signal_953}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_319 ( .clk (signal_2371), .D ({signal_2090, signal_954}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_321 ( .clk (signal_2371), .D ({signal_2089, signal_955}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_323 ( .clk (signal_2371), .D ({signal_2088, signal_956}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_325 ( .clk (signal_2371), .D ({signal_2060, signal_957}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_327 ( .clk (signal_2371), .D ({signal_2087, signal_958}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_329 ( .clk (signal_2371), .D ({signal_2098, signal_959}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_331 ( .clk (signal_2371), .D ({signal_2097, signal_960}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_333 ( .clk (signal_2371), .D ({signal_2072, signal_961}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_335 ( .clk (signal_2371), .D ({signal_2096, signal_962}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_337 ( .clk (signal_2371), .D ({signal_2095, signal_963}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_339 ( .clk (signal_2371), .D ({signal_2094, signal_964}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_341 ( .clk (signal_2371), .D ({signal_2068, signal_965}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_343 ( .clk (signal_2371), .D ({signal_2093, signal_966}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_345 ( .clk (signal_2371), .D ({signal_2040, signal_967}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_347 ( .clk (signal_2371), .D ({signal_2039, signal_968}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_349 ( .clk (signal_2371), .D ({signal_1984, signal_969}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_351 ( .clk (signal_2371), .D ({signal_2038, signal_970}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_353 ( .clk (signal_2371), .D ({signal_2037, signal_971}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_355 ( .clk (signal_2371), .D ({signal_2036, signal_972}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_357 ( .clk (signal_2371), .D ({signal_1980, signal_973}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_359 ( .clk (signal_2371), .D ({signal_2035, signal_974}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_361 ( .clk (signal_2371), .D ({signal_2034, signal_975}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_363 ( .clk (signal_2371), .D ({signal_2033, signal_976}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_365 ( .clk (signal_2371), .D ({signal_1976, signal_977}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_367 ( .clk (signal_2371), .D ({signal_2032, signal_978}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_369 ( .clk (signal_2371), .D ({signal_2031, signal_979}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_371 ( .clk (signal_2371), .D ({signal_2030, signal_980}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_373 ( .clk (signal_2371), .D ({signal_1972, signal_981}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_375 ( .clk (signal_2371), .D ({signal_2029, signal_982}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_377 ( .clk (signal_2371), .D ({signal_2028, signal_983}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_379 ( .clk (signal_2371), .D ({signal_2027, signal_984}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_381 ( .clk (signal_2371), .D ({signal_1968, signal_985}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_383 ( .clk (signal_2371), .D ({signal_2026, signal_986}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_385 ( .clk (signal_2371), .D ({signal_2025, signal_987}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_387 ( .clk (signal_2371), .D ({signal_2024, signal_988}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_389 ( .clk (signal_2371), .D ({signal_1964, signal_989}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_391 ( .clk (signal_2371), .D ({signal_2023, signal_990}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_393 ( .clk (signal_2371), .D ({signal_2022, signal_991}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_395 ( .clk (signal_2371), .D ({signal_2021, signal_992}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_397 ( .clk (signal_2371), .D ({signal_1960, signal_993}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_399 ( .clk (signal_2371), .D ({signal_2020, signal_994}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_401 ( .clk (signal_2371), .D ({signal_2019, signal_995}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_403 ( .clk (signal_2371), .D ({signal_2018, signal_996}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_405 ( .clk (signal_2371), .D ({signal_1956, signal_997}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_407 ( .clk (signal_2371), .D ({signal_2017, signal_998}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    DFF_X1 cell_789 ( .CK (signal_2371), .D (signal_1008), .Q (signal_1001), .QN () ) ;
    DFF_X1 cell_791 ( .CK (signal_2371), .D (signal_1009), .Q (signal_1002), .QN () ) ;
    DFF_X1 cell_793 ( .CK (signal_2371), .D (signal_1010), .Q (signal_1003), .QN () ) ;
    DFF_X1 cell_795 ( .CK (signal_2371), .D (signal_1011), .Q (signal_1004), .QN () ) ;
    DFF_X1 cell_797 ( .CK (signal_2371), .D (signal_1012), .Q (signal_1005), .QN () ) ;
    DFF_X1 cell_799 ( .CK (signal_2371), .D (signal_1013), .Q (signal_1006), .QN () ) ;
    DFF_X1 cell_801 ( .CK (signal_2371), .D (signal_1014), .Q (signal_1007), .QN () ) ;
    DFF_X1 cell_814 ( .CK (signal_2371), .D (signal_1017), .Q (signal_1015), .QN () ) ;
    DFF_X1 cell_816 ( .CK (signal_2371), .D (signal_1018), .Q (signal_1016), .QN () ) ;
    DFF_X1 cell_818 ( .CK (signal_2371), .D (signal_267), .Q (done), .QN () ) ;
endmodule
