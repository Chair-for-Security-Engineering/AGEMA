/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d1 (X_s0, clk, X_s1, Fresh, Y_s0, Y_s1);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [33:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_277 ;
    wire signal_279 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_284 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_136 ( .a ({X_s1[7], X_s0[7]}), .b ({X_s1[4], X_s0[4]}), .c ({signal_277, signal_151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_137 ( .a ({X_s1[7], X_s0[7]}), .b ({X_s1[2], X_s0[2]}), .c ({signal_279, signal_152}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_138 ( .a ({X_s1[7], X_s0[7]}), .b ({X_s1[1], X_s0[1]}), .c ({signal_281, signal_153}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_139 ( .a ({X_s1[4], X_s0[4]}), .b ({X_s1[2], X_s0[2]}), .c ({signal_282, signal_154}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_140 ( .a ({X_s1[3], X_s0[3]}), .b ({X_s1[1], X_s0[1]}), .c ({signal_284, signal_155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_141 ( .a ({X_s1[6], X_s0[6]}), .b ({X_s1[5], X_s0[5]}), .c ({signal_287, signal_156}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_142 ( .a ({X_s1[6], X_s0[6]}), .b ({X_s1[2], X_s0[2]}), .c ({signal_288, signal_157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_143 ( .a ({X_s1[5], X_s0[5]}), .b ({X_s1[2], X_s0[2]}), .c ({signal_289, signal_158}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_144 ( .a ({X_s1[4], X_s0[4]}), .b ({X_s1[0], X_s0[0]}), .c ({signal_291, signal_159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_145 ( .a ({X_s1[1], X_s0[1]}), .b ({X_s1[0], X_s0[0]}), .c ({signal_292, signal_160}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_146 ( .a ({signal_277, signal_151}), .b ({signal_284, signal_155}), .c ({signal_293, signal_161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_147 ( .a ({X_s1[0], X_s0[0]}), .b ({signal_287, signal_156}), .c ({signal_294, signal_162}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_148 ( .a ({signal_281, signal_153}), .b ({signal_282, signal_154}), .c ({signal_295, signal_163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_149 ( .a ({signal_284, signal_155}), .b ({signal_288, signal_157}), .c ({signal_296, signal_164}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_150 ( .a ({signal_284, signal_155}), .b ({signal_289, signal_158}), .c ({signal_297, signal_165}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_151 ( .a ({signal_287, signal_156}), .b ({signal_291, signal_159}), .c ({signal_298, signal_166}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_152 ( .a ({signal_287, signal_156}), .b ({signal_292, signal_160}), .c ({signal_299, signal_167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_153 ( .a ({signal_277, signal_151}), .b ({signal_289, signal_158}), .c ({signal_300, signal_168}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_160 ( .a ({X_s1[0], X_s0[0]}), .b ({signal_293, signal_161}), .c ({signal_307, signal_175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_161 ( .a ({signal_287, signal_156}), .b ({signal_293, signal_161}), .c ({signal_308, signal_176}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_162 ( .a ({signal_288, signal_157}), .b ({signal_293, signal_161}), .c ({signal_309, signal_177}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_163 ( .a ({signal_294, signal_162}), .b ({signal_297, signal_165}), .c ({signal_310, signal_178}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_164 ( .a ({signal_277, signal_151}), .b ({signal_298, signal_166}), .c ({signal_311, signal_179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_165 ( .a ({signal_279, signal_152}), .b ({signal_299, signal_167}), .c ({signal_312, signal_180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_166 ( .a ({signal_281, signal_153}), .b ({signal_297, signal_165}), .c ({signal_313, signal_181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_170 ( .a ({signal_279, signal_152}), .b ({signal_308, signal_176}), .c ({signal_317, signal_185}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_171 ( .a ({signal_310, signal_178}), .b ({signal_311, signal_179}), .c ({signal_318, signal_186}) ) ;

    /* cells in depth 1 */
    buf_clk cell_268 ( .C (clk), .D (signal_177), .Q (signal_457) ) ;
    buf_clk cell_270 ( .C (clk), .D (signal_309), .Q (signal_459) ) ;
    buf_clk cell_272 ( .C (clk), .D (signal_181), .Q (signal_461) ) ;
    buf_clk cell_274 ( .C (clk), .D (signal_313), .Q (signal_463) ) ;
    buf_clk cell_276 ( .C (clk), .D (signal_185), .Q (signal_465) ) ;
    buf_clk cell_278 ( .C (clk), .D (signal_317), .Q (signal_467) ) ;
    buf_clk cell_280 ( .C (clk), .D (signal_186), .Q (signal_469) ) ;
    buf_clk cell_282 ( .C (clk), .D (signal_318), .Q (signal_471) ) ;
    buf_clk cell_316 ( .C (clk), .D (signal_175), .Q (signal_505) ) ;
    buf_clk cell_322 ( .C (clk), .D (signal_307), .Q (signal_511) ) ;
    buf_clk cell_328 ( .C (clk), .D (X_s0[0]), .Q (signal_517) ) ;
    buf_clk cell_334 ( .C (clk), .D (X_s1[0]), .Q (signal_523) ) ;
    buf_clk cell_340 ( .C (clk), .D (signal_162), .Q (signal_529) ) ;
    buf_clk cell_346 ( .C (clk), .D (signal_294), .Q (signal_535) ) ;
    buf_clk cell_352 ( .C (clk), .D (signal_178), .Q (signal_541) ) ;
    buf_clk cell_358 ( .C (clk), .D (signal_310), .Q (signal_547) ) ;
    buf_clk cell_364 ( .C (clk), .D (signal_180), .Q (signal_553) ) ;
    buf_clk cell_370 ( .C (clk), .D (signal_312), .Q (signal_559) ) ;
    buf_clk cell_376 ( .C (clk), .D (signal_166), .Q (signal_565) ) ;
    buf_clk cell_382 ( .C (clk), .D (signal_298), .Q (signal_571) ) ;
    buf_clk cell_388 ( .C (clk), .D (signal_167), .Q (signal_577) ) ;
    buf_clk cell_394 ( .C (clk), .D (signal_299), .Q (signal_583) ) ;
    buf_clk cell_400 ( .C (clk), .D (signal_179), .Q (signal_589) ) ;
    buf_clk cell_406 ( .C (clk), .D (signal_311), .Q (signal_595) ) ;
    buf_clk cell_412 ( .C (clk), .D (signal_161), .Q (signal_601) ) ;
    buf_clk cell_418 ( .C (clk), .D (signal_293), .Q (signal_607) ) ;
    buf_clk cell_424 ( .C (clk), .D (signal_165), .Q (signal_613) ) ;
    buf_clk cell_430 ( .C (clk), .D (signal_297), .Q (signal_619) ) ;
    buf_clk cell_436 ( .C (clk), .D (signal_164), .Q (signal_625) ) ;
    buf_clk cell_442 ( .C (clk), .D (signal_296), .Q (signal_631) ) ;
    buf_clk cell_448 ( .C (clk), .D (signal_176), .Q (signal_637) ) ;
    buf_clk cell_454 ( .C (clk), .D (signal_308), .Q (signal_643) ) ;
    buf_clk cell_460 ( .C (clk), .D (signal_163), .Q (signal_649) ) ;
    buf_clk cell_466 ( .C (clk), .D (signal_295), .Q (signal_655) ) ;
    buf_clk cell_472 ( .C (clk), .D (signal_153), .Q (signal_661) ) ;
    buf_clk cell_478 ( .C (clk), .D (signal_281), .Q (signal_667) ) ;
    buf_clk cell_484 ( .C (clk), .D (signal_151), .Q (signal_673) ) ;
    buf_clk cell_490 ( .C (clk), .D (signal_277), .Q (signal_679) ) ;
    buf_clk cell_496 ( .C (clk), .D (signal_152), .Q (signal_685) ) ;
    buf_clk cell_502 ( .C (clk), .D (signal_279), .Q (signal_691) ) ;
    buf_clk cell_508 ( .C (clk), .D (signal_168), .Q (signal_697) ) ;
    buf_clk cell_514 ( .C (clk), .D (signal_300), .Q (signal_703) ) ;
    buf_clk cell_520 ( .C (clk), .D (signal_154), .Q (signal_709) ) ;
    buf_clk cell_526 ( .C (clk), .D (signal_282), .Q (signal_715) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_154 ( .a ({signal_293, signal_161}), .b ({signal_295, signal_163}), .clk (clk), .r (Fresh[0]), .c ({signal_301, signal_169}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_155 ( .a ({X_s1[0], X_s0[0]}), .b ({signal_298, signal_166}), .clk (clk), .r (Fresh[1]), .c ({signal_302, signal_170}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_156 ( .a ({signal_281, signal_153}), .b ({signal_297, signal_165}), .clk (clk), .r (Fresh[2]), .c ({signal_303, signal_171}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_157 ( .a ({signal_294, signal_162}), .b ({signal_299, signal_167}), .clk (clk), .r (Fresh[3]), .c ({signal_304, signal_172}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_158 ( .a ({signal_277, signal_151}), .b ({signal_296, signal_164}), .clk (clk), .r (Fresh[4]), .c ({signal_305, signal_173}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_159 ( .a ({signal_282, signal_154}), .b ({signal_300, signal_168}), .clk (clk), .r (Fresh[5]), .c ({signal_306, signal_174}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_167 ( .a ({signal_307, signal_175}), .b ({signal_312, signal_180}), .clk (clk), .r (Fresh[6]), .c ({signal_314, signal_182}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_168 ( .a ({signal_310, signal_178}), .b ({signal_311, signal_179}), .clk (clk), .r (Fresh[7]), .c ({signal_315, signal_183}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_169 ( .a ({signal_279, signal_152}), .b ({signal_308, signal_176}), .clk (clk), .r (Fresh[8]), .c ({signal_316, signal_184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_172 ( .a ({signal_460, signal_458}), .b ({signal_301, signal_169}), .c ({signal_319, signal_187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_173 ( .a ({signal_301, signal_169}), .b ({signal_302, signal_170}), .c ({signal_320, signal_188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_174 ( .a ({signal_464, signal_462}), .b ({signal_303, signal_171}), .c ({signal_321, signal_189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_175 ( .a ({signal_305, signal_173}), .b ({signal_306, signal_174}), .c ({signal_322, signal_190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_176 ( .a ({signal_303, signal_171}), .b ({signal_315, signal_183}), .c ({signal_323, signal_191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_177 ( .a ({signal_305, signal_173}), .b ({signal_316, signal_184}), .c ({signal_324, signal_192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_178 ( .a ({signal_314, signal_182}), .b ({signal_319, signal_187}), .c ({signal_325, signal_193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_179 ( .a ({signal_468, signal_466}), .b ({signal_320, signal_188}), .c ({signal_326, signal_194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_180 ( .a ({signal_304, signal_172}), .b ({signal_321, signal_189}), .c ({signal_327, signal_195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_181 ( .a ({signal_323, signal_191}), .b ({signal_324, signal_192}), .c ({signal_328, signal_196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_182 ( .a ({signal_322, signal_190}), .b ({signal_325, signal_193}), .c ({signal_329, signal_197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_183 ( .a ({signal_324, signal_192}), .b ({signal_326, signal_194}), .c ({signal_330, signal_198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_184 ( .a ({signal_322, signal_190}), .b ({signal_327, signal_195}), .c ({signal_331, signal_199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_187 ( .a ({signal_472, signal_470}), .b ({signal_328, signal_196}), .c ({signal_334, signal_202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_188 ( .a ({signal_329, signal_197}), .b ({signal_330, signal_198}), .c ({signal_335, signal_203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_190 ( .a ({signal_331, signal_199}), .b ({signal_334, signal_202}), .c ({signal_337, signal_205}) ) ;
    buf_clk cell_269 ( .C (clk), .D (signal_457), .Q (signal_458) ) ;
    buf_clk cell_271 ( .C (clk), .D (signal_459), .Q (signal_460) ) ;
    buf_clk cell_273 ( .C (clk), .D (signal_461), .Q (signal_462) ) ;
    buf_clk cell_275 ( .C (clk), .D (signal_463), .Q (signal_464) ) ;
    buf_clk cell_277 ( .C (clk), .D (signal_465), .Q (signal_466) ) ;
    buf_clk cell_279 ( .C (clk), .D (signal_467), .Q (signal_468) ) ;
    buf_clk cell_281 ( .C (clk), .D (signal_469), .Q (signal_470) ) ;
    buf_clk cell_283 ( .C (clk), .D (signal_471), .Q (signal_472) ) ;
    buf_clk cell_317 ( .C (clk), .D (signal_505), .Q (signal_506) ) ;
    buf_clk cell_323 ( .C (clk), .D (signal_511), .Q (signal_512) ) ;
    buf_clk cell_329 ( .C (clk), .D (signal_517), .Q (signal_518) ) ;
    buf_clk cell_335 ( .C (clk), .D (signal_523), .Q (signal_524) ) ;
    buf_clk cell_341 ( .C (clk), .D (signal_529), .Q (signal_530) ) ;
    buf_clk cell_347 ( .C (clk), .D (signal_535), .Q (signal_536) ) ;
    buf_clk cell_353 ( .C (clk), .D (signal_541), .Q (signal_542) ) ;
    buf_clk cell_359 ( .C (clk), .D (signal_547), .Q (signal_548) ) ;
    buf_clk cell_365 ( .C (clk), .D (signal_553), .Q (signal_554) ) ;
    buf_clk cell_371 ( .C (clk), .D (signal_559), .Q (signal_560) ) ;
    buf_clk cell_377 ( .C (clk), .D (signal_565), .Q (signal_566) ) ;
    buf_clk cell_383 ( .C (clk), .D (signal_571), .Q (signal_572) ) ;
    buf_clk cell_389 ( .C (clk), .D (signal_577), .Q (signal_578) ) ;
    buf_clk cell_395 ( .C (clk), .D (signal_583), .Q (signal_584) ) ;
    buf_clk cell_401 ( .C (clk), .D (signal_589), .Q (signal_590) ) ;
    buf_clk cell_407 ( .C (clk), .D (signal_595), .Q (signal_596) ) ;
    buf_clk cell_413 ( .C (clk), .D (signal_601), .Q (signal_602) ) ;
    buf_clk cell_419 ( .C (clk), .D (signal_607), .Q (signal_608) ) ;
    buf_clk cell_425 ( .C (clk), .D (signal_613), .Q (signal_614) ) ;
    buf_clk cell_431 ( .C (clk), .D (signal_619), .Q (signal_620) ) ;
    buf_clk cell_437 ( .C (clk), .D (signal_625), .Q (signal_626) ) ;
    buf_clk cell_443 ( .C (clk), .D (signal_631), .Q (signal_632) ) ;
    buf_clk cell_449 ( .C (clk), .D (signal_637), .Q (signal_638) ) ;
    buf_clk cell_455 ( .C (clk), .D (signal_643), .Q (signal_644) ) ;
    buf_clk cell_461 ( .C (clk), .D (signal_649), .Q (signal_650) ) ;
    buf_clk cell_467 ( .C (clk), .D (signal_655), .Q (signal_656) ) ;
    buf_clk cell_473 ( .C (clk), .D (signal_661), .Q (signal_662) ) ;
    buf_clk cell_479 ( .C (clk), .D (signal_667), .Q (signal_668) ) ;
    buf_clk cell_485 ( .C (clk), .D (signal_673), .Q (signal_674) ) ;
    buf_clk cell_491 ( .C (clk), .D (signal_679), .Q (signal_680) ) ;
    buf_clk cell_497 ( .C (clk), .D (signal_685), .Q (signal_686) ) ;
    buf_clk cell_503 ( .C (clk), .D (signal_691), .Q (signal_692) ) ;
    buf_clk cell_509 ( .C (clk), .D (signal_697), .Q (signal_698) ) ;
    buf_clk cell_515 ( .C (clk), .D (signal_703), .Q (signal_704) ) ;
    buf_clk cell_521 ( .C (clk), .D (signal_709), .Q (signal_710) ) ;
    buf_clk cell_527 ( .C (clk), .D (signal_715), .Q (signal_716) ) ;

    /* cells in depth 3 */
    buf_clk cell_284 ( .C (clk), .D (signal_198), .Q (signal_473) ) ;
    buf_clk cell_286 ( .C (clk), .D (signal_330), .Q (signal_475) ) ;
    buf_clk cell_288 ( .C (clk), .D (signal_202), .Q (signal_477) ) ;
    buf_clk cell_290 ( .C (clk), .D (signal_334), .Q (signal_479) ) ;
    buf_clk cell_292 ( .C (clk), .D (signal_203), .Q (signal_481) ) ;
    buf_clk cell_294 ( .C (clk), .D (signal_335), .Q (signal_483) ) ;
    buf_clk cell_296 ( .C (clk), .D (signal_205), .Q (signal_485) ) ;
    buf_clk cell_298 ( .C (clk), .D (signal_337), .Q (signal_487) ) ;
    buf_clk cell_318 ( .C (clk), .D (signal_506), .Q (signal_507) ) ;
    buf_clk cell_324 ( .C (clk), .D (signal_512), .Q (signal_513) ) ;
    buf_clk cell_330 ( .C (clk), .D (signal_518), .Q (signal_519) ) ;
    buf_clk cell_336 ( .C (clk), .D (signal_524), .Q (signal_525) ) ;
    buf_clk cell_342 ( .C (clk), .D (signal_530), .Q (signal_531) ) ;
    buf_clk cell_348 ( .C (clk), .D (signal_536), .Q (signal_537) ) ;
    buf_clk cell_354 ( .C (clk), .D (signal_542), .Q (signal_543) ) ;
    buf_clk cell_360 ( .C (clk), .D (signal_548), .Q (signal_549) ) ;
    buf_clk cell_366 ( .C (clk), .D (signal_554), .Q (signal_555) ) ;
    buf_clk cell_372 ( .C (clk), .D (signal_560), .Q (signal_561) ) ;
    buf_clk cell_378 ( .C (clk), .D (signal_566), .Q (signal_567) ) ;
    buf_clk cell_384 ( .C (clk), .D (signal_572), .Q (signal_573) ) ;
    buf_clk cell_390 ( .C (clk), .D (signal_578), .Q (signal_579) ) ;
    buf_clk cell_396 ( .C (clk), .D (signal_584), .Q (signal_585) ) ;
    buf_clk cell_402 ( .C (clk), .D (signal_590), .Q (signal_591) ) ;
    buf_clk cell_408 ( .C (clk), .D (signal_596), .Q (signal_597) ) ;
    buf_clk cell_414 ( .C (clk), .D (signal_602), .Q (signal_603) ) ;
    buf_clk cell_420 ( .C (clk), .D (signal_608), .Q (signal_609) ) ;
    buf_clk cell_426 ( .C (clk), .D (signal_614), .Q (signal_615) ) ;
    buf_clk cell_432 ( .C (clk), .D (signal_620), .Q (signal_621) ) ;
    buf_clk cell_438 ( .C (clk), .D (signal_626), .Q (signal_627) ) ;
    buf_clk cell_444 ( .C (clk), .D (signal_632), .Q (signal_633) ) ;
    buf_clk cell_450 ( .C (clk), .D (signal_638), .Q (signal_639) ) ;
    buf_clk cell_456 ( .C (clk), .D (signal_644), .Q (signal_645) ) ;
    buf_clk cell_462 ( .C (clk), .D (signal_650), .Q (signal_651) ) ;
    buf_clk cell_468 ( .C (clk), .D (signal_656), .Q (signal_657) ) ;
    buf_clk cell_474 ( .C (clk), .D (signal_662), .Q (signal_663) ) ;
    buf_clk cell_480 ( .C (clk), .D (signal_668), .Q (signal_669) ) ;
    buf_clk cell_486 ( .C (clk), .D (signal_674), .Q (signal_675) ) ;
    buf_clk cell_492 ( .C (clk), .D (signal_680), .Q (signal_681) ) ;
    buf_clk cell_498 ( .C (clk), .D (signal_686), .Q (signal_687) ) ;
    buf_clk cell_504 ( .C (clk), .D (signal_692), .Q (signal_693) ) ;
    buf_clk cell_510 ( .C (clk), .D (signal_698), .Q (signal_699) ) ;
    buf_clk cell_516 ( .C (clk), .D (signal_704), .Q (signal_705) ) ;
    buf_clk cell_522 ( .C (clk), .D (signal_710), .Q (signal_711) ) ;
    buf_clk cell_528 ( .C (clk), .D (signal_716), .Q (signal_717) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_185 ( .a ({signal_329, signal_197}), .b ({signal_331, signal_199}), .clk (clk), .r (Fresh[9]), .c ({signal_332, signal_200}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_186 ( .a ({signal_330, signal_198}), .b ({signal_331, signal_199}), .clk (clk), .r (Fresh[10]), .c ({signal_333, signal_201}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_189 ( .a ({signal_329, signal_197}), .b ({signal_334, signal_202}), .clk (clk), .r (Fresh[11]), .c ({signal_336, signal_204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_191 ( .a ({signal_476, signal_474}), .b ({signal_332, signal_200}), .c ({signal_338, signal_206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_192 ( .a ({signal_480, signal_478}), .b ({signal_332, signal_200}), .c ({signal_339, signal_207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_193 ( .a ({signal_332, signal_200}), .b ({signal_484, signal_482}), .c ({signal_340, signal_208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_198 ( .a ({signal_332, signal_200}), .b ({signal_488, signal_486}), .c ({signal_345, signal_213}) ) ;
    buf_clk cell_285 ( .C (clk), .D (signal_473), .Q (signal_474) ) ;
    buf_clk cell_287 ( .C (clk), .D (signal_475), .Q (signal_476) ) ;
    buf_clk cell_289 ( .C (clk), .D (signal_477), .Q (signal_478) ) ;
    buf_clk cell_291 ( .C (clk), .D (signal_479), .Q (signal_480) ) ;
    buf_clk cell_293 ( .C (clk), .D (signal_481), .Q (signal_482) ) ;
    buf_clk cell_295 ( .C (clk), .D (signal_483), .Q (signal_484) ) ;
    buf_clk cell_297 ( .C (clk), .D (signal_485), .Q (signal_486) ) ;
    buf_clk cell_299 ( .C (clk), .D (signal_487), .Q (signal_488) ) ;
    buf_clk cell_319 ( .C (clk), .D (signal_507), .Q (signal_508) ) ;
    buf_clk cell_325 ( .C (clk), .D (signal_513), .Q (signal_514) ) ;
    buf_clk cell_331 ( .C (clk), .D (signal_519), .Q (signal_520) ) ;
    buf_clk cell_337 ( .C (clk), .D (signal_525), .Q (signal_526) ) ;
    buf_clk cell_343 ( .C (clk), .D (signal_531), .Q (signal_532) ) ;
    buf_clk cell_349 ( .C (clk), .D (signal_537), .Q (signal_538) ) ;
    buf_clk cell_355 ( .C (clk), .D (signal_543), .Q (signal_544) ) ;
    buf_clk cell_361 ( .C (clk), .D (signal_549), .Q (signal_550) ) ;
    buf_clk cell_367 ( .C (clk), .D (signal_555), .Q (signal_556) ) ;
    buf_clk cell_373 ( .C (clk), .D (signal_561), .Q (signal_562) ) ;
    buf_clk cell_379 ( .C (clk), .D (signal_567), .Q (signal_568) ) ;
    buf_clk cell_385 ( .C (clk), .D (signal_573), .Q (signal_574) ) ;
    buf_clk cell_391 ( .C (clk), .D (signal_579), .Q (signal_580) ) ;
    buf_clk cell_397 ( .C (clk), .D (signal_585), .Q (signal_586) ) ;
    buf_clk cell_403 ( .C (clk), .D (signal_591), .Q (signal_592) ) ;
    buf_clk cell_409 ( .C (clk), .D (signal_597), .Q (signal_598) ) ;
    buf_clk cell_415 ( .C (clk), .D (signal_603), .Q (signal_604) ) ;
    buf_clk cell_421 ( .C (clk), .D (signal_609), .Q (signal_610) ) ;
    buf_clk cell_427 ( .C (clk), .D (signal_615), .Q (signal_616) ) ;
    buf_clk cell_433 ( .C (clk), .D (signal_621), .Q (signal_622) ) ;
    buf_clk cell_439 ( .C (clk), .D (signal_627), .Q (signal_628) ) ;
    buf_clk cell_445 ( .C (clk), .D (signal_633), .Q (signal_634) ) ;
    buf_clk cell_451 ( .C (clk), .D (signal_639), .Q (signal_640) ) ;
    buf_clk cell_457 ( .C (clk), .D (signal_645), .Q (signal_646) ) ;
    buf_clk cell_463 ( .C (clk), .D (signal_651), .Q (signal_652) ) ;
    buf_clk cell_469 ( .C (clk), .D (signal_657), .Q (signal_658) ) ;
    buf_clk cell_475 ( .C (clk), .D (signal_663), .Q (signal_664) ) ;
    buf_clk cell_481 ( .C (clk), .D (signal_669), .Q (signal_670) ) ;
    buf_clk cell_487 ( .C (clk), .D (signal_675), .Q (signal_676) ) ;
    buf_clk cell_493 ( .C (clk), .D (signal_681), .Q (signal_682) ) ;
    buf_clk cell_499 ( .C (clk), .D (signal_687), .Q (signal_688) ) ;
    buf_clk cell_505 ( .C (clk), .D (signal_693), .Q (signal_694) ) ;
    buf_clk cell_511 ( .C (clk), .D (signal_699), .Q (signal_700) ) ;
    buf_clk cell_517 ( .C (clk), .D (signal_705), .Q (signal_706) ) ;
    buf_clk cell_523 ( .C (clk), .D (signal_711), .Q (signal_712) ) ;
    buf_clk cell_529 ( .C (clk), .D (signal_717), .Q (signal_718) ) ;

    /* cells in depth 5 */
    buf_clk cell_300 ( .C (clk), .D (signal_474), .Q (signal_489) ) ;
    buf_clk cell_302 ( .C (clk), .D (signal_476), .Q (signal_491) ) ;
    buf_clk cell_304 ( .C (clk), .D (signal_208), .Q (signal_493) ) ;
    buf_clk cell_306 ( .C (clk), .D (signal_340), .Q (signal_495) ) ;
    buf_clk cell_308 ( .C (clk), .D (signal_478), .Q (signal_497) ) ;
    buf_clk cell_310 ( .C (clk), .D (signal_480), .Q (signal_499) ) ;
    buf_clk cell_312 ( .C (clk), .D (signal_213), .Q (signal_501) ) ;
    buf_clk cell_314 ( .C (clk), .D (signal_345), .Q (signal_503) ) ;
    buf_clk cell_320 ( .C (clk), .D (signal_508), .Q (signal_509) ) ;
    buf_clk cell_326 ( .C (clk), .D (signal_514), .Q (signal_515) ) ;
    buf_clk cell_332 ( .C (clk), .D (signal_520), .Q (signal_521) ) ;
    buf_clk cell_338 ( .C (clk), .D (signal_526), .Q (signal_527) ) ;
    buf_clk cell_344 ( .C (clk), .D (signal_532), .Q (signal_533) ) ;
    buf_clk cell_350 ( .C (clk), .D (signal_538), .Q (signal_539) ) ;
    buf_clk cell_356 ( .C (clk), .D (signal_544), .Q (signal_545) ) ;
    buf_clk cell_362 ( .C (clk), .D (signal_550), .Q (signal_551) ) ;
    buf_clk cell_368 ( .C (clk), .D (signal_556), .Q (signal_557) ) ;
    buf_clk cell_374 ( .C (clk), .D (signal_562), .Q (signal_563) ) ;
    buf_clk cell_380 ( .C (clk), .D (signal_568), .Q (signal_569) ) ;
    buf_clk cell_386 ( .C (clk), .D (signal_574), .Q (signal_575) ) ;
    buf_clk cell_392 ( .C (clk), .D (signal_580), .Q (signal_581) ) ;
    buf_clk cell_398 ( .C (clk), .D (signal_586), .Q (signal_587) ) ;
    buf_clk cell_404 ( .C (clk), .D (signal_592), .Q (signal_593) ) ;
    buf_clk cell_410 ( .C (clk), .D (signal_598), .Q (signal_599) ) ;
    buf_clk cell_416 ( .C (clk), .D (signal_604), .Q (signal_605) ) ;
    buf_clk cell_422 ( .C (clk), .D (signal_610), .Q (signal_611) ) ;
    buf_clk cell_428 ( .C (clk), .D (signal_616), .Q (signal_617) ) ;
    buf_clk cell_434 ( .C (clk), .D (signal_622), .Q (signal_623) ) ;
    buf_clk cell_440 ( .C (clk), .D (signal_628), .Q (signal_629) ) ;
    buf_clk cell_446 ( .C (clk), .D (signal_634), .Q (signal_635) ) ;
    buf_clk cell_452 ( .C (clk), .D (signal_640), .Q (signal_641) ) ;
    buf_clk cell_458 ( .C (clk), .D (signal_646), .Q (signal_647) ) ;
    buf_clk cell_464 ( .C (clk), .D (signal_652), .Q (signal_653) ) ;
    buf_clk cell_470 ( .C (clk), .D (signal_658), .Q (signal_659) ) ;
    buf_clk cell_476 ( .C (clk), .D (signal_664), .Q (signal_665) ) ;
    buf_clk cell_482 ( .C (clk), .D (signal_670), .Q (signal_671) ) ;
    buf_clk cell_488 ( .C (clk), .D (signal_676), .Q (signal_677) ) ;
    buf_clk cell_494 ( .C (clk), .D (signal_682), .Q (signal_683) ) ;
    buf_clk cell_500 ( .C (clk), .D (signal_688), .Q (signal_689) ) ;
    buf_clk cell_506 ( .C (clk), .D (signal_694), .Q (signal_695) ) ;
    buf_clk cell_512 ( .C (clk), .D (signal_700), .Q (signal_701) ) ;
    buf_clk cell_518 ( .C (clk), .D (signal_706), .Q (signal_707) ) ;
    buf_clk cell_524 ( .C (clk), .D (signal_712), .Q (signal_713) ) ;
    buf_clk cell_530 ( .C (clk), .D (signal_718), .Q (signal_719) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_194 ( .a ({signal_484, signal_482}), .b ({signal_339, signal_207}), .clk (clk), .r (Fresh[12]), .c ({signal_341, signal_209}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_195 ( .a ({signal_488, signal_486}), .b ({signal_338, signal_206}), .clk (clk), .r (Fresh[13]), .c ({signal_342, signal_210}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_196 ( .a ({signal_484, signal_482}), .b ({signal_336, signal_204}), .clk (clk), .r (Fresh[14]), .c ({signal_343, signal_211}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_197 ( .a ({signal_333, signal_201}), .b ({signal_488, signal_486}), .clk (clk), .r (Fresh[15]), .c ({signal_344, signal_212}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_199 ( .a ({signal_492, signal_490}), .b ({signal_341, signal_209}), .c ({signal_346, signal_214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_200 ( .a ({signal_496, signal_494}), .b ({signal_343, signal_211}), .c ({signal_347, signal_215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_201 ( .a ({signal_500, signal_498}), .b ({signal_342, signal_210}), .c ({signal_348, signal_216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_202 ( .a ({signal_344, signal_212}), .b ({signal_504, signal_502}), .c ({signal_349, signal_217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_211 ( .a ({signal_347, signal_215}), .b ({signal_349, signal_217}), .c ({signal_358, signal_226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_212 ( .a ({signal_346, signal_214}), .b ({signal_348, signal_216}), .c ({signal_359, signal_227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_213 ( .a ({signal_346, signal_214}), .b ({signal_347, signal_215}), .c ({signal_360, signal_228}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_214 ( .a ({signal_348, signal_216}), .b ({signal_349, signal_217}), .c ({signal_361, signal_229}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_223 ( .a ({signal_358, signal_226}), .b ({signal_359, signal_227}), .c ({signal_370, signal_238}) ) ;
    buf_clk cell_301 ( .C (clk), .D (signal_489), .Q (signal_490) ) ;
    buf_clk cell_303 ( .C (clk), .D (signal_491), .Q (signal_492) ) ;
    buf_clk cell_305 ( .C (clk), .D (signal_493), .Q (signal_494) ) ;
    buf_clk cell_307 ( .C (clk), .D (signal_495), .Q (signal_496) ) ;
    buf_clk cell_309 ( .C (clk), .D (signal_497), .Q (signal_498) ) ;
    buf_clk cell_311 ( .C (clk), .D (signal_499), .Q (signal_500) ) ;
    buf_clk cell_313 ( .C (clk), .D (signal_501), .Q (signal_502) ) ;
    buf_clk cell_315 ( .C (clk), .D (signal_503), .Q (signal_504) ) ;
    buf_clk cell_321 ( .C (clk), .D (signal_509), .Q (signal_510) ) ;
    buf_clk cell_327 ( .C (clk), .D (signal_515), .Q (signal_516) ) ;
    buf_clk cell_333 ( .C (clk), .D (signal_521), .Q (signal_522) ) ;
    buf_clk cell_339 ( .C (clk), .D (signal_527), .Q (signal_528) ) ;
    buf_clk cell_345 ( .C (clk), .D (signal_533), .Q (signal_534) ) ;
    buf_clk cell_351 ( .C (clk), .D (signal_539), .Q (signal_540) ) ;
    buf_clk cell_357 ( .C (clk), .D (signal_545), .Q (signal_546) ) ;
    buf_clk cell_363 ( .C (clk), .D (signal_551), .Q (signal_552) ) ;
    buf_clk cell_369 ( .C (clk), .D (signal_557), .Q (signal_558) ) ;
    buf_clk cell_375 ( .C (clk), .D (signal_563), .Q (signal_564) ) ;
    buf_clk cell_381 ( .C (clk), .D (signal_569), .Q (signal_570) ) ;
    buf_clk cell_387 ( .C (clk), .D (signal_575), .Q (signal_576) ) ;
    buf_clk cell_393 ( .C (clk), .D (signal_581), .Q (signal_582) ) ;
    buf_clk cell_399 ( .C (clk), .D (signal_587), .Q (signal_588) ) ;
    buf_clk cell_405 ( .C (clk), .D (signal_593), .Q (signal_594) ) ;
    buf_clk cell_411 ( .C (clk), .D (signal_599), .Q (signal_600) ) ;
    buf_clk cell_417 ( .C (clk), .D (signal_605), .Q (signal_606) ) ;
    buf_clk cell_423 ( .C (clk), .D (signal_611), .Q (signal_612) ) ;
    buf_clk cell_429 ( .C (clk), .D (signal_617), .Q (signal_618) ) ;
    buf_clk cell_435 ( .C (clk), .D (signal_623), .Q (signal_624) ) ;
    buf_clk cell_441 ( .C (clk), .D (signal_629), .Q (signal_630) ) ;
    buf_clk cell_447 ( .C (clk), .D (signal_635), .Q (signal_636) ) ;
    buf_clk cell_453 ( .C (clk), .D (signal_641), .Q (signal_642) ) ;
    buf_clk cell_459 ( .C (clk), .D (signal_647), .Q (signal_648) ) ;
    buf_clk cell_465 ( .C (clk), .D (signal_653), .Q (signal_654) ) ;
    buf_clk cell_471 ( .C (clk), .D (signal_659), .Q (signal_660) ) ;
    buf_clk cell_477 ( .C (clk), .D (signal_665), .Q (signal_666) ) ;
    buf_clk cell_483 ( .C (clk), .D (signal_671), .Q (signal_672) ) ;
    buf_clk cell_489 ( .C (clk), .D (signal_677), .Q (signal_678) ) ;
    buf_clk cell_495 ( .C (clk), .D (signal_683), .Q (signal_684) ) ;
    buf_clk cell_501 ( .C (clk), .D (signal_689), .Q (signal_690) ) ;
    buf_clk cell_507 ( .C (clk), .D (signal_695), .Q (signal_696) ) ;
    buf_clk cell_513 ( .C (clk), .D (signal_701), .Q (signal_702) ) ;
    buf_clk cell_519 ( .C (clk), .D (signal_707), .Q (signal_708) ) ;
    buf_clk cell_525 ( .C (clk), .D (signal_713), .Q (signal_714) ) ;
    buf_clk cell_531 ( .C (clk), .D (signal_719), .Q (signal_720) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_203 ( .a ({signal_516, signal_510}), .b ({signal_349, signal_217}), .clk (clk), .r (Fresh[16]), .c ({signal_350, signal_218}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_204 ( .a ({signal_528, signal_522}), .b ({signal_348, signal_216}), .clk (clk), .r (Fresh[17]), .c ({signal_351, signal_219}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_205 ( .a ({signal_540, signal_534}), .b ({signal_347, signal_215}), .clk (clk), .r (Fresh[18]), .c ({signal_352, signal_220}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_206 ( .a ({signal_552, signal_546}), .b ({signal_346, signal_214}), .clk (clk), .r (Fresh[19]), .c ({signal_353, signal_221}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_207 ( .a ({signal_564, signal_558}), .b ({signal_349, signal_217}), .clk (clk), .r (Fresh[20]), .c ({signal_354, signal_222}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_208 ( .a ({signal_576, signal_570}), .b ({signal_348, signal_216}), .clk (clk), .r (Fresh[21]), .c ({signal_355, signal_223}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_209 ( .a ({signal_588, signal_582}), .b ({signal_347, signal_215}), .clk (clk), .r (Fresh[22]), .c ({signal_356, signal_224}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_210 ( .a ({signal_600, signal_594}), .b ({signal_346, signal_214}), .clk (clk), .r (Fresh[23]), .c ({signal_357, signal_225}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_215 ( .a ({signal_612, signal_606}), .b ({signal_361, signal_229}), .clk (clk), .r (Fresh[24]), .c ({signal_362, signal_230}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_216 ( .a ({signal_624, signal_618}), .b ({signal_360, signal_228}), .clk (clk), .r (Fresh[25]), .c ({signal_363, signal_231}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_217 ( .a ({signal_636, signal_630}), .b ({signal_359, signal_227}), .clk (clk), .r (Fresh[26]), .c ({signal_364, signal_232}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_218 ( .a ({signal_648, signal_642}), .b ({signal_358, signal_226}), .clk (clk), .r (Fresh[27]), .c ({signal_365, signal_233}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_219 ( .a ({signal_660, signal_654}), .b ({signal_361, signal_229}), .clk (clk), .r (Fresh[28]), .c ({signal_366, signal_234}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_220 ( .a ({signal_672, signal_666}), .b ({signal_360, signal_228}), .clk (clk), .r (Fresh[29]), .c ({signal_367, signal_235}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_221 ( .a ({signal_684, signal_678}), .b ({signal_359, signal_227}), .clk (clk), .r (Fresh[30]), .c ({signal_368, signal_236}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_222 ( .a ({signal_696, signal_690}), .b ({signal_358, signal_226}), .clk (clk), .r (Fresh[31]), .c ({signal_369, signal_237}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_224 ( .a ({signal_352, signal_220}), .b ({signal_354, signal_222}), .c ({signal_371, signal_239}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_225 ( .a ({signal_353, signal_221}), .b ({signal_356, signal_224}), .c ({signal_372, signal_240}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_226 ( .a ({signal_351, signal_219}), .b ({signal_353, signal_221}), .c ({signal_373, signal_241}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_227 ( .a ({signal_708, signal_702}), .b ({signal_370, signal_238}), .clk (clk), .r (Fresh[32]), .c ({signal_374, signal_242}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_228 ( .a ({signal_720, signal_714}), .b ({signal_370, signal_238}), .clk (clk), .r (Fresh[33]), .c ({signal_375, signal_243}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_229 ( .a ({signal_351, signal_219}), .b ({signal_362, signal_230}), .c ({signal_376, signal_244}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_230 ( .a ({signal_350, signal_218}), .b ({signal_366, signal_234}), .c ({signal_377, signal_245}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_231 ( .a ({signal_365, signal_233}), .b ({signal_367, signal_235}), .c ({signal_378, signal_246}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_232 ( .a ({signal_363, signal_231}), .b ({signal_368, signal_236}), .c ({signal_379, signal_247}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_233 ( .a ({signal_364, signal_232}), .b ({signal_368, signal_236}), .c ({signal_380, signal_248}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_234 ( .a ({signal_366, signal_234}), .b ({signal_371, signal_239}), .c ({signal_381, signal_249}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_235 ( .a ({signal_355, signal_223}), .b ({signal_371, signal_239}), .c ({signal_382, signal_250}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_236 ( .a ({signal_367, signal_235}), .b ({signal_372, signal_240}), .c ({signal_383, signal_251}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_237 ( .a ({signal_368, signal_236}), .b ({signal_375, signal_243}), .c ({signal_384, signal_252}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_238 ( .a ({signal_375, signal_243}), .b ({signal_379, signal_247}), .c ({signal_385, signal_253}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_239 ( .a ({signal_362, signal_230}), .b ({signal_377, signal_245}), .c ({signal_386, signal_254}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_240 ( .a ({signal_364, signal_232}), .b ({signal_374, signal_242}), .c ({signal_387, signal_255}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_241 ( .a ({signal_374, signal_242}), .b ({signal_378, signal_246}), .c ({signal_388, signal_256}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_242 ( .a ({signal_357, signal_225}), .b ({signal_376, signal_244}), .c ({signal_389, signal_257}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_243 ( .a ({signal_369, signal_237}), .b ({signal_378, signal_246}), .c ({signal_390, signal_258}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_244 ( .a ({signal_373, signal_241}), .b ({signal_377, signal_245}), .c ({signal_391, signal_259}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_245 ( .a ({signal_376, signal_244}), .b ({signal_383, signal_251}), .c ({signal_392, signal_260}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_246 ( .a ({signal_352, signal_220}), .b ({signal_384, signal_252}), .c ({signal_393, signal_261}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_247 ( .a ({signal_354, signal_222}), .b ({signal_384, signal_252}), .c ({signal_394, signal_262}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_248 ( .a ({signal_371, signal_239}), .b ({signal_384, signal_252}), .c ({signal_395, signal_263}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_249 ( .a ({signal_371, signal_239}), .b ({signal_386, signal_254}), .c ({signal_396, signal_264}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_250 ( .a ({signal_381, signal_249}), .b ({signal_387, signal_255}), .c ({signal_397, signal_265}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_251 ( .a ({signal_385, signal_253}), .b ({signal_388, signal_256}), .c ({signal_398, signal_266}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_252 ( .a ({signal_386, signal_254}), .b ({signal_387, signal_255}), .c ({signal_399, signal_267}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_253 ( .a ({signal_372, signal_240}), .b ({signal_388, signal_256}), .c ({signal_400, signal_268}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_254 ( .a ({signal_380, signal_248}), .b ({signal_389, signal_257}), .c ({signal_401, signal_269}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_255 ( .a ({signal_382, signal_250}), .b ({signal_389, signal_257}), .c ({signal_402, signal_270}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_256 ( .a ({signal_385, signal_253}), .b ({signal_392, signal_260}), .c ({signal_403, signal_271}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_257 ( .a ({signal_403, signal_271}), .b ({signal_404, signal_150}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_258 ( .a ({signal_385, signal_253}), .b ({signal_397, signal_265}), .c ({signal_405, signal_143}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_259 ( .a ({signal_394, signal_262}), .b ({signal_399, signal_267}), .c ({signal_406, signal_272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_260 ( .a ({signal_390, signal_258}), .b ({signal_401, signal_269}), .c ({signal_407, signal_273}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_261 ( .a ({signal_385, signal_253}), .b ({signal_396, signal_264}), .c ({signal_408, signal_146}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_262 ( .a ({signal_391, signal_259}), .b ({signal_395, signal_263}), .c ({signal_409, signal_147}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_263 ( .a ({signal_398, signal_266}), .b ({signal_402, signal_270}), .c ({signal_410, signal_148}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_264 ( .a ({signal_393, signal_261}), .b ({signal_400, signal_268}), .c ({signal_411, signal_274}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_265 ( .a ({signal_406, signal_272}), .b ({signal_412, signal_144}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_266 ( .a ({signal_407, signal_273}), .b ({signal_413, signal_145}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_267 ( .a ({signal_411, signal_274}), .b ({signal_414, signal_149}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_405, signal_143}), .Q ({Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_412, signal_144}), .Q ({Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_413, signal_145}), .Q ({Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_408, signal_146}), .Q ({Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_4 ( .clk (clk), .D ({signal_409, signal_147}), .Q ({Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_5 ( .clk (clk), .D ({signal_410, signal_148}), .Q ({Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_6 ( .clk (clk), .D ({signal_414, signal_149}), .Q ({Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_7 ( .clk (clk), .D ({signal_404, signal_150}), .Q ({Y_s1[0], Y_s0[0]}) ) ;
endmodule
