module Reg1(x, y);
 input [75:0] x;
 output [74:0] y;

  register_stage #(.WIDTH(75)) inst_0(.clk(x[0]), .D({x[75],x[5],x[6],x[7],x[8],x[9],x[10],x[1],x[2],x[3],x[4],x[11],x[22],x[33],x[44],x[55],x[66],x[71],x[72],x[73],x[74],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[67],x[68],x[69],x[70]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74]}));
endmodule

module Reg2(x, y);
 input [150:0] x;
 output [149:0] y;

  register_stage #(.WIDTH(150)) inst_0(.clk(x[0]), .D({x[149],x[150],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[21],x[22],x[43],x[44],x[65],x[66],x[87],x[88],x[109],x[110],x[131],x[132],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx1(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx2(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx3(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx6(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx7(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx8(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx11(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx12(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx13(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx16(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx17(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx18(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx21(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx22(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx23(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx26(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx27(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx33(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [224:0] x;
 output [149:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx1 Fx1_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx2 Fx2_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx3 Fx3_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx4 Fx4_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx5 Fx5_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx6 Fx6_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx7 Fx7_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx8 Fx8_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx9 Fx9_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx10 Fx10_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx11 Fx11_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx12 Fx12_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx13 Fx13_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx14 Fx14_inst(.x({x[22], x[21]}), .y(y[14]));
  Fx15 Fx15_inst(.x({x[23], x[21]}), .y(y[15]));
  Fx16 Fx16_inst(.x({x[25], x[24]}), .y(y[16]));
  Fx17 Fx17_inst(.x({x[26], x[24]}), .y(y[17]));
  Fx18 Fx18_inst(.x({x[28], x[27]}), .y(y[18]));
  Fx19 Fx19_inst(.x({x[29], x[27]}), .y(y[19]));
  Fx20 Fx20_inst(.x({x[31], x[30]}), .y(y[20]));
  Fx21 Fx21_inst(.x({x[32], x[30]}), .y(y[21]));
  Fx22 Fx22_inst(.x({x[34], x[33]}), .y(y[22]));
  Fx23 Fx23_inst(.x({x[35], x[33]}), .y(y[23]));
  Fx24 Fx24_inst(.x({x[37], x[36]}), .y(y[24]));
  Fx25 Fx25_inst(.x({x[38], x[36]}), .y(y[25]));
  Fx26 Fx26_inst(.x({x[40], x[39]}), .y(y[26]));
  Fx27 Fx27_inst(.x({x[41], x[39]}), .y(y[27]));
  Fx28 Fx28_inst(.x({x[43], x[42]}), .y(y[28]));
  Fx29 Fx29_inst(.x({x[44], x[42]}), .y(y[29]));
  Fx30 Fx30_inst(.x({x[46], x[45]}), .y(y[30]));
  Fx31 Fx31_inst(.x({x[47], x[45]}), .y(y[31]));
  Fx32 Fx32_inst(.x({x[49], x[48]}), .y(y[32]));
  Fx33 Fx33_inst(.x({x[50], x[48]}), .y(y[33]));
  Fx34 Fx34_inst(.x({x[52], x[51]}), .y(y[34]));
  Fx35 Fx35_inst(.x({x[53], x[51]}), .y(y[35]));
  Fx36 Fx36_inst(.x({x[55], x[54]}), .y(y[36]));
  Fx37 Fx37_inst(.x({x[56], x[54]}), .y(y[37]));
  Fx38 Fx38_inst(.x({x[58], x[57]}), .y(y[38]));
  Fx39 Fx39_inst(.x({x[59], x[57]}), .y(y[39]));
  Fx40 Fx40_inst(.x({x[61], x[60]}), .y(y[40]));
  Fx41 Fx41_inst(.x({x[62], x[60]}), .y(y[41]));
  Fx42 Fx42_inst(.x({x[64], x[63]}), .y(y[42]));
  Fx43 Fx43_inst(.x({x[65], x[63]}), .y(y[43]));
  Fx44 Fx44_inst(.x({x[67], x[66]}), .y(y[44]));
  Fx45 Fx45_inst(.x({x[68], x[66]}), .y(y[45]));
  Fx46 Fx46_inst(.x({x[70], x[69]}), .y(y[46]));
  Fx47 Fx47_inst(.x({x[71], x[69]}), .y(y[47]));
  Fx48 Fx48_inst(.x({x[73], x[72]}), .y(y[48]));
  Fx49 Fx49_inst(.x({x[74], x[72]}), .y(y[49]));
  Fx50 Fx50_inst(.x({x[76], x[75]}), .y(y[50]));
  Fx51 Fx51_inst(.x({x[77], x[75]}), .y(y[51]));
  Fx52 Fx52_inst(.x({x[79], x[78]}), .y(y[52]));
  Fx53 Fx53_inst(.x({x[80], x[78]}), .y(y[53]));
  Fx54 Fx54_inst(.x({x[82], x[81]}), .y(y[54]));
  Fx55 Fx55_inst(.x({x[83], x[81]}), .y(y[55]));
  Fx56 Fx56_inst(.x({x[85], x[84]}), .y(y[56]));
  Fx57 Fx57_inst(.x({x[86], x[84]}), .y(y[57]));
  Fx58 Fx58_inst(.x({x[88], x[87]}), .y(y[58]));
  Fx59 Fx59_inst(.x({x[89], x[87]}), .y(y[59]));
  Fx60 Fx60_inst(.x({x[91], x[90]}), .y(y[60]));
  Fx61 Fx61_inst(.x({x[92], x[90]}), .y(y[61]));
  Fx62 Fx62_inst(.x({x[94], x[93]}), .y(y[62]));
  Fx63 Fx63_inst(.x({x[95], x[93]}), .y(y[63]));
  Fx64 Fx64_inst(.x({x[97], x[96]}), .y(y[64]));
  Fx65 Fx65_inst(.x({x[98], x[96]}), .y(y[65]));
  Fx66 Fx66_inst(.x({x[100], x[99]}), .y(y[66]));
  Fx67 Fx67_inst(.x({x[101], x[99]}), .y(y[67]));
  Fx68 Fx68_inst(.x({x[103], x[102]}), .y(y[68]));
  Fx69 Fx69_inst(.x({x[104], x[102]}), .y(y[69]));
  Fx70 Fx70_inst(.x({x[106], x[105]}), .y(y[70]));
  Fx71 Fx71_inst(.x({x[107], x[105]}), .y(y[71]));
  Fx72 Fx72_inst(.x({x[109], x[108]}), .y(y[72]));
  Fx73 Fx73_inst(.x({x[110], x[108]}), .y(y[73]));
  Fx74 Fx74_inst(.x({x[112], x[111]}), .y(y[74]));
  Fx75 Fx75_inst(.x({x[113], x[111]}), .y(y[75]));
  Fx76 Fx76_inst(.x({x[115], x[114]}), .y(y[76]));
  Fx77 Fx77_inst(.x({x[116], x[114]}), .y(y[77]));
  Fx78 Fx78_inst(.x({x[118], x[117]}), .y(y[78]));
  Fx79 Fx79_inst(.x({x[119], x[117]}), .y(y[79]));
  Fx80 Fx80_inst(.x({x[121], x[120]}), .y(y[80]));
  Fx81 Fx81_inst(.x({x[122], x[120]}), .y(y[81]));
  Fx82 Fx82_inst(.x({x[124], x[123]}), .y(y[82]));
  Fx83 Fx83_inst(.x({x[125], x[123]}), .y(y[83]));
  Fx84 Fx84_inst(.x({x[127], x[126]}), .y(y[84]));
  Fx85 Fx85_inst(.x({x[128], x[126]}), .y(y[85]));
  Fx86 Fx86_inst(.x({x[130], x[129]}), .y(y[86]));
  Fx87 Fx87_inst(.x({x[131], x[129]}), .y(y[87]));
  Fx88 Fx88_inst(.x({x[133], x[132]}), .y(y[88]));
  Fx89 Fx89_inst(.x({x[134], x[132]}), .y(y[89]));
  Fx90 Fx90_inst(.x({x[136], x[135]}), .y(y[90]));
  Fx91 Fx91_inst(.x({x[137], x[135]}), .y(y[91]));
  Fx92 Fx92_inst(.x({x[139], x[138]}), .y(y[92]));
  Fx93 Fx93_inst(.x({x[140], x[138]}), .y(y[93]));
  Fx94 Fx94_inst(.x({x[142], x[141]}), .y(y[94]));
  Fx95 Fx95_inst(.x({x[143], x[141]}), .y(y[95]));
  Fx96 Fx96_inst(.x({x[145], x[144]}), .y(y[96]));
  Fx97 Fx97_inst(.x({x[146], x[144]}), .y(y[97]));
  Fx98 Fx98_inst(.x({x[148], x[147]}), .y(y[98]));
  Fx99 Fx99_inst(.x({x[149], x[147]}), .y(y[99]));
  Fx100 Fx100_inst(.x({x[151], x[150]}), .y(y[100]));
  Fx101 Fx101_inst(.x({x[152], x[150]}), .y(y[101]));
  Fx102 Fx102_inst(.x({x[154], x[153]}), .y(y[102]));
  Fx103 Fx103_inst(.x({x[155], x[153]}), .y(y[103]));
  Fx104 Fx104_inst(.x({x[157], x[156]}), .y(y[104]));
  Fx105 Fx105_inst(.x({x[158], x[156]}), .y(y[105]));
  Fx106 Fx106_inst(.x({x[160], x[159]}), .y(y[106]));
  Fx107 Fx107_inst(.x({x[161], x[159]}), .y(y[107]));
  Fx108 Fx108_inst(.x({x[163], x[162]}), .y(y[108]));
  Fx109 Fx109_inst(.x({x[164], x[162]}), .y(y[109]));
  Fx110 Fx110_inst(.x({x[166], x[165]}), .y(y[110]));
  Fx111 Fx111_inst(.x({x[167], x[165]}), .y(y[111]));
  Fx112 Fx112_inst(.x({x[169], x[168]}), .y(y[112]));
  Fx113 Fx113_inst(.x({x[170], x[168]}), .y(y[113]));
  Fx114 Fx114_inst(.x({x[172], x[171]}), .y(y[114]));
  Fx115 Fx115_inst(.x({x[173], x[171]}), .y(y[115]));
  Fx116 Fx116_inst(.x({x[175], x[174]}), .y(y[116]));
  Fx117 Fx117_inst(.x({x[176], x[174]}), .y(y[117]));
  Fx118 Fx118_inst(.x({x[178], x[177]}), .y(y[118]));
  Fx119 Fx119_inst(.x({x[179], x[177]}), .y(y[119]));
  Fx120 Fx120_inst(.x({x[181], x[180]}), .y(y[120]));
  Fx121 Fx121_inst(.x({x[182], x[180]}), .y(y[121]));
  Fx122 Fx122_inst(.x({x[184], x[183]}), .y(y[122]));
  Fx123 Fx123_inst(.x({x[185], x[183]}), .y(y[123]));
  Fx124 Fx124_inst(.x({x[187], x[186]}), .y(y[124]));
  Fx125 Fx125_inst(.x({x[188], x[186]}), .y(y[125]));
  Fx126 Fx126_inst(.x({x[190], x[189]}), .y(y[126]));
  Fx127 Fx127_inst(.x({x[191], x[189]}), .y(y[127]));
  Fx128 Fx128_inst(.x({x[193], x[192]}), .y(y[128]));
  Fx129 Fx129_inst(.x({x[194], x[192]}), .y(y[129]));
  Fx130 Fx130_inst(.x({x[196], x[195]}), .y(y[130]));
  Fx131 Fx131_inst(.x({x[197], x[195]}), .y(y[131]));
  Fx132 Fx132_inst(.x({x[199], x[198]}), .y(y[132]));
  Fx133 Fx133_inst(.x({x[200], x[198]}), .y(y[133]));
  Fx134 Fx134_inst(.x({x[202], x[201]}), .y(y[134]));
  Fx135 Fx135_inst(.x({x[203], x[201]}), .y(y[135]));
  Fx136 Fx136_inst(.x({x[205], x[204]}), .y(y[136]));
  Fx137 Fx137_inst(.x({x[206], x[204]}), .y(y[137]));
  Fx138 Fx138_inst(.x({x[208], x[207]}), .y(y[138]));
  Fx139 Fx139_inst(.x({x[209], x[207]}), .y(y[139]));
  Fx140 Fx140_inst(.x({x[211], x[210]}), .y(y[140]));
  Fx141 Fx141_inst(.x({x[212], x[210]}), .y(y[141]));
  Fx142 Fx142_inst(.x({x[214], x[213]}), .y(y[142]));
  Fx143 Fx143_inst(.x({x[215], x[213]}), .y(y[143]));
  Fx144 Fx144_inst(.x({x[217], x[216]}), .y(y[144]));
  Fx145 Fx145_inst(.x({x[218], x[216]}), .y(y[145]));
  Fx146 Fx146_inst(.x({x[220], x[219]}), .y(y[146]));
  Fx147 Fx147_inst(.x({x[221], x[219]}), .y(y[147]));
  Fx148 Fx148_inst(.x({x[223], x[222]}), .y(y[148]));
  Fx149 Fx149_inst(.x({x[224], x[222]}), .y(y[149]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [21:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~(t[6] | t[1]);
  assign t[10] = t[17] ^ x[15];
  assign t[11] = t[18] ^ x[18];
  assign t[12] = t[19] ^ x[21];
  assign t[13] = (x[1] & x[2]);
  assign t[14] = (x[4] & x[5]);
  assign t[15] = (x[7] & x[8]);
  assign t[16] = (x[10] & x[11]);
  assign t[17] = (x[13] & x[14]);
  assign t[18] = (x[16] & x[17]);
  assign t[19] = (x[19] & x[20]);
  assign t[1] = ~(t[7] | t[2]);
  assign t[2] = ~(t[8] & t[3]);
  assign t[3] = ~(t[9] | t[4]);
  assign t[4] = ~(t[10] & t[5]);
  assign t[5] = ~(t[11] | t[12]);
  assign t[6] = t[13] ^ x[3];
  assign t[7] = t[14] ^ x[6];
  assign t[8] = t[15] ^ x[9];
  assign t[9] = t[16] ^ x[12];
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind66(x, y);
 input [116:0] x;
 output y;

 wire [262:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[27] ? x[50] : x[49];
  assign t[101] = t[27] ? x[52] : x[51];
  assign t[102] = t[219] ^ t[142];
  assign t[103] = ~(t[143] & t[144]);
  assign t[104] = t[145] ^ t[224];
  assign t[105] = ~(t[220]);
  assign t[106] = t[146] & t[145];
  assign t[107] = t[86] ^ t[126];
  assign t[108] = t[147] & t[148];
  assign t[109] = t[131] ? t[149] : t[225];
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = t[111] ^ t[61];
  assign t[111] = t[150] ^ t[151];
  assign t[112] = t[152] & t[153];
  assign t[113] = t[26] ? t[154] : t[226];
  assign t[114] = t[155] ^ t[58];
  assign t[115] = t[126] ^ t[77];
  assign t[116] = t[114] ^ t[156];
  assign t[117] = t[157] ^ t[128];
  assign t[118] = t[158] & t[159];
  assign t[119] = t[62] ^ t[160];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[140] ^ t[97];
  assign t[121] = t[157] ^ t[123];
  assign t[122] = t[161] & t[162];
  assign t[123] = t[217] ^ t[163];
  assign t[124] = t[129] ^ t[118];
  assign t[125] = t[26] ? t[164] : t[227];
  assign t[126] = t[165];
  assign t[127] = t[26] ? t[166] : t[228];
  assign t[128] = t[210] ^ t[167];
  assign t[129] = t[168] ^ t[122];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[169] & t[170];
  assign t[131] = ~(t[14]);
  assign t[132] = t[222] ^ t[171];
  assign t[133] = t[223] ^ t[172];
  assign t[134] = t[131] ? t[173] : t[229];
  assign t[135] = t[27] ? x[72] : x[71];
  assign t[136] = ~(t[141]);
  assign t[137] = ~(t[41]);
  assign t[138] = ~(t[42]);
  assign t[139] = t[39] ^ t[41];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[41] ^ t[62];
  assign t[141] = t[67] ^ t[42];
  assign t[142] = t[27] ? x[74] : x[73];
  assign t[143] = ~(t[146] | t[145]);
  assign t[144] = ~(t[174] | t[105]);
  assign t[145] = ~(t[230]);
  assign t[146] = ~(t[224]);
  assign t[147] = ~(t[107] ^ t[114]);
  assign t[148] = t[115] ^ t[88];
  assign t[149] = t[225] ^ t[175];
  assign t[14] = ~(t[26]);
  assign t[150] = t[176] & t[177];
  assign t[151] = t[178] & t[134];
  assign t[152] = ~(t[150] ^ t[179]);
  assign t[153] = t[180] ^ t[181];
  assign t[154] = t[226] ^ t[182];
  assign t[155] = t[183] & t[184];
  assign t[156] = t[185] & t[186];
  assign t[157] = t[7] ? t[187] : t[231];
  assign t[158] = ~(t[117] ^ t[129]);
  assign t[159] = t[89] ^ t[162];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[63] ^ t[25];
  assign t[161] = ~(t[128]);
  assign t[162] = t[211] ^ t[188];
  assign t[163] = t[7] ? t[189] : t[232];
  assign t[164] = t[227] ^ t[190];
  assign t[165] = t[26] ? t[191] : t[233];
  assign t[166] = t[228] ^ t[192];
  assign t[167] = t[26] ? t[193] : t[234];
  assign t[168] = t[194] & t[195];
  assign t[169] = ~(t[168] ^ t[196]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[121] ^ t[197];
  assign t[171] = t[198] ? x[91] : x[90];
  assign t[172] = t[198] ? x[93] : x[92];
  assign t[173] = t[229] ^ t[199];
  assign t[174] = ~(t[215]);
  assign t[175] = t[198] ? x[95] : x[94];
  assign t[176] = ~(t[181]);
  assign t[177] = ~(t[91]);
  assign t[178] = ~(t[92]);
  assign t[179] = t[75] ^ t[91];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[91] ^ t[109];
  assign t[181] = t[134] ^ t[92];
  assign t[182] = t[71] ? x[97] : x[96];
  assign t[183] = ~(t[200]);
  assign t[184] = ~(t[86]);
  assign t[185] = ~(t[155] ^ t[201]);
  assign t[186] = t[57] ^ t[200];
  assign t[187] = t[231] ^ t[202];
  assign t[188] = t[7] ? t[203] : t[235];
  assign t[189] = t[232] ^ t[204];
  assign t[18] = ~(t[23] ^ t[32]);
  assign t[190] = t[71] ? x[102] : x[101];
  assign t[191] = t[233] ^ t[205];
  assign t[192] = t[27] ? x[104] : x[103];
  assign t[193] = t[234] ^ t[206];
  assign t[194] = ~(t[197]);
  assign t[195] = ~(t[157]);
  assign t[196] = t[89] ^ t[157];
  assign t[197] = t[162] ^ t[128];
  assign t[198] = ~(t[47]);
  assign t[199] = t[198] ? x[106] : x[105];
  assign t[19] = ~(t[33] ^ t[34]);
  assign t[1] = ~(t[4]);
  assign t[200] = t[88] ^ t[126];
  assign t[201] = t[115] ^ t[86];
  assign t[202] = t[71] ? x[108] : x[107];
  assign t[203] = t[235] ^ t[207];
  assign t[204] = t[71] ? x[110] : x[109];
  assign t[205] = t[208] ? x[112] : x[111];
  assign t[206] = t[208] ? x[114] : x[113];
  assign t[207] = t[208] ? x[116] : x[115];
  assign t[208] = ~(t[47]);
  assign t[209] = t[236] ^ x[4];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[237] ^ x[9];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[37] ^ t[13]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[55];
  assign t[225] = t[252] ^ x[58];
  assign t[226] = t[253] ^ x[61];
  assign t[227] = t[254] ^ x[64];
  assign t[228] = t[255] ^ x[67];
  assign t[229] = t[256] ^ x[70];
  assign t[22] = ~(t[37] ^ t[38]);
  assign t[230] = t[257] ^ x[77];
  assign t[231] = t[258] ^ x[80];
  assign t[232] = t[259] ^ x[83];
  assign t[233] = t[260] ^ x[86];
  assign t[234] = t[261] ^ x[89];
  assign t[235] = t[262] ^ x[100];
  assign t[236] = (x[2] & x[3]);
  assign t[237] = (x[7] & x[8]);
  assign t[238] = (x[10] & x[11]);
  assign t[239] = (x[13] & x[14]);
  assign t[23] = t[39] ^ t[40];
  assign t[240] = (x[16] & x[17]);
  assign t[241] = (x[19] & x[20]);
  assign t[242] = (x[22] & x[23]);
  assign t[243] = (x[25] & x[26]);
  assign t[244] = (x[28] & x[29]);
  assign t[245] = (x[31] & x[32]);
  assign t[246] = (x[34] & x[35]);
  assign t[247] = (x[37] & x[38]);
  assign t[248] = (x[40] & x[41]);
  assign t[249] = (x[43] & x[44]);
  assign t[24] = t[41] ^ t[42];
  assign t[250] = (x[46] & x[47]);
  assign t[251] = (x[53] & x[54]);
  assign t[252] = (x[56] & x[57]);
  assign t[253] = (x[59] & x[60]);
  assign t[254] = (x[62] & x[63]);
  assign t[255] = (x[65] & x[66]);
  assign t[256] = (x[68] & x[69]);
  assign t[257] = (x[75] & x[76]);
  assign t[258] = (x[78] & x[79]);
  assign t[259] = (x[81] & x[82]);
  assign t[25] = t[43] & t[44];
  assign t[260] = (x[84] & x[85]);
  assign t[261] = (x[87] & x[88]);
  assign t[262] = (x[98] & x[99]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[210]);
  assign t[29] = ~(t[211]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[212]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = ~(t[50] ^ t[51]);
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[34] = t[12] ^ t[54];
  assign t[35] = ~(t[55] ^ t[56]);
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ t[52];
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[42] ^ t[62];
  assign t[3] = t[7] ? t[8] : t[209];
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[7] ? t[65] : t[213];
  assign t[42] = t[7] ? t[66] : t[214];
  assign t[43] = ~(t[24] ^ t[63]);
  assign t[44] = t[39] ^ t[67];
  assign t[45] = ~(t[68] & t[69]);
  assign t[46] = t[215] | t[70];
  assign t[47] = ~(t[71]);
  assign t[48] = ~(t[216]);
  assign t[49] = ~(t[72] & t[217]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[73] ^ t[74]);
  assign t[51] = t[75] ^ t[76];
  assign t[52] = t[77] ^ t[78];
  assign t[53] = t[79] ^ t[80];
  assign t[54] = ~(t[81] ^ t[82]);
  assign t[55] = t[83] ^ t[32];
  assign t[56] = ~(t[84] ^ t[85]);
  assign t[57] = t[86] ^ t[77];
  assign t[58] = t[87] & t[88];
  assign t[59] = t[89] ^ t[90];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[91] ^ t[92];
  assign t[61] = t[93] & t[94];
  assign t[62] = t[7] ? t[95] : t[218];
  assign t[63] = t[96] ^ t[97];
  assign t[64] = t[98] & t[99];
  assign t[65] = t[213] ^ t[100];
  assign t[66] = t[214] ^ t[101];
  assign t[67] = t[7] ? t[102] : t[219];
  assign t[68] = ~(t[70] & t[103]);
  assign t[69] = ~(t[220] ^ t[104]);
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[105] & t[106]);
  assign t[71] = ~(t[46]);
  assign t[72] = ~(t[221]);
  assign t[73] = t[107] ^ t[108];
  assign t[74] = t[109] ^ t[110];
  assign t[75] = t[92] ^ t[109];
  assign t[76] = t[111] ^ t[112];
  assign t[77] = ~t[113];
  assign t[78] = t[114] ^ t[108];
  assign t[79] = t[115] ^ t[116];
  assign t[7] = ~(t[14]);
  assign t[80] = t[117] ^ t[118];
  assign t[81] = t[51] ^ t[36];
  assign t[82] = ~(t[119] ^ t[85]);
  assign t[83] = t[119] ^ t[120];
  assign t[84] = t[121] ^ t[122];
  assign t[85] = t[123] ^ t[124];
  assign t[86] = ~t[125];
  assign t[87] = ~(t[126]);
  assign t[88] = t[127];
  assign t[89] = t[128] ^ t[123];
  assign t[8] = t[209] ^ t[15];
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[131] ? t[132] : t[222];
  assign t[92] = t[131] ? t[133] : t[223];
  assign t[93] = ~(t[60] ^ t[111]);
  assign t[94] = t[75] ^ t[134];
  assign t[95] = t[218] ^ t[135];
  assign t[96] = t[136] & t[137];
  assign t[97] = t[138] & t[67];
  assign t[98] = ~(t[96] ^ t[139]);
  assign t[99] = t[140] ^ t[141];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind67(x, y);
 input [116:0] x;
 output y;

 wire [264:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[212] ^ t[139];
  assign t[101] = t[140] ^ t[105];
  assign t[102] = t[141] & t[142];
  assign t[103] = t[7] ? t[143] : t[226];
  assign t[104] = t[122] ^ t[66];
  assign t[105] = t[144] & t[145];
  assign t[106] = t[7] ? t[146] : t[227];
  assign t[107] = t[118] ^ t[53];
  assign t[108] = t[147] ^ t[120];
  assign t[109] = ~(t[148] & t[149]);
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = t[150] ^ t[228];
  assign t[111] = ~(t[219]);
  assign t[112] = t[151] & t[150];
  assign t[113] = t[221] ^ t[152];
  assign t[114] = t[87] ? t[153] : t[229];
  assign t[115] = t[222] ^ t[154];
  assign t[116] = t[223] ^ t[155];
  assign t[117] = t[224] ^ t[156];
  assign t[118] = t[157] ^ t[158];
  assign t[119] = t[7] ? t[159] : t[230];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[160];
  assign t[121] = t[161] & t[162];
  assign t[122] = t[7] ? t[163] : t[231];
  assign t[123] = ~(t[85] ^ t[101]);
  assign t[124] = t[64] ^ t[145];
  assign t[125] = t[164] ? x[68] : x[67];
  assign t[126] = t[165] & t[166];
  assign t[127] = ~(t[134] ^ t[89]);
  assign t[128] = t[136] ^ t[78];
  assign t[129] = t[225] ^ t[167];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[168] & t[169];
  assign t[131] = t[170] & t[171];
  assign t[132] = ~(t[108] ^ t[92]);
  assign t[133] = t[83] ^ t[171];
  assign t[134] = t[76] ^ t[114];
  assign t[135] = t[172] & t[173];
  assign t[136] = t[114] ^ t[56];
  assign t[137] = t[89] ^ t[174];
  assign t[138] = t[147] ^ t[58];
  assign t[139] = t[26] ? t[175] : t[232];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[176] & t[177];
  assign t[141] = ~(t[140] ^ t[178]);
  assign t[142] = t[104] ^ t[179];
  assign t[143] = t[226] ^ t[180];
  assign t[144] = ~(t[100]);
  assign t[145] = t[213] ^ t[181];
  assign t[146] = t[227] ^ t[182];
  assign t[147] = ~t[183];
  assign t[148] = ~(t[151] | t[150]);
  assign t[149] = ~(t[184] | t[111]);
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[233]);
  assign t[151] = ~(t[228]);
  assign t[152] = t[164] ? x[76] : x[75];
  assign t[153] = t[229] ^ t[185];
  assign t[154] = t[164] ? x[78] : x[77];
  assign t[155] = t[27] ? x[80] : x[79];
  assign t[156] = t[27] ? x[82] : x[81];
  assign t[157] = t[186] & t[187];
  assign t[158] = t[188] & t[119];
  assign t[159] = t[230] ^ t[189];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[26] ? t[190] : t[234];
  assign t[161] = ~(t[130] ^ t[191]);
  assign t[162] = t[138] ^ t[192];
  assign t[163] = t[231] ^ t[193];
  assign t[164] = ~(t[47]);
  assign t[165] = ~(t[194]);
  assign t[166] = ~(t[76]);
  assign t[167] = t[74] ? x[87] : x[86];
  assign t[168] = ~(t[192]);
  assign t[169] = ~(t[147]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = ~(t[120]);
  assign t[171] = t[195];
  assign t[172] = ~(t[157] ^ t[196]);
  assign t[173] = t[197] ^ t[198];
  assign t[174] = t[199] & t[200];
  assign t[175] = t[232] ^ t[201];
  assign t[176] = ~(t[179]);
  assign t[177] = ~(t[122]);
  assign t[178] = t[64] ^ t[122];
  assign t[179] = t[145] ^ t[100];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[74] ? x[89] : x[88];
  assign t[181] = t[7] ? t[202] : t[235];
  assign t[182] = t[27] ? x[94] : x[93];
  assign t[183] = t[26] ? t[203] : t[236];
  assign t[184] = ~(t[215]);
  assign t[185] = t[164] ? x[99] : x[98];
  assign t[186] = ~(t[198]);
  assign t[187] = ~(t[79]);
  assign t[188] = ~(t[80]);
  assign t[189] = t[27] ? x[101] : x[100];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[234] ^ t[204];
  assign t[191] = t[83] ^ t[147];
  assign t[192] = t[171] ^ t[120];
  assign t[193] = t[74] ? x[103] : x[102];
  assign t[194] = t[78] ^ t[114];
  assign t[195] = t[26] ? t[205] : t[237];
  assign t[196] = t[96] ^ t[79];
  assign t[197] = t[79] ^ t[106];
  assign t[198] = t[119] ^ t[80];
  assign t[199] = ~(t[126] ^ t[206]);
  assign t[19] = ~(t[34] ^ t[35]);
  assign t[1] = ~(t[4]);
  assign t[200] = t[50] ^ t[194];
  assign t[201] = t[207] ? x[108] : x[107];
  assign t[202] = t[235] ^ t[208];
  assign t[203] = t[236] ^ t[209];
  assign t[204] = t[207] ? x[110] : x[109];
  assign t[205] = t[237] ^ t[210];
  assign t[206] = t[136] ^ t[76];
  assign t[207] = ~(t[47]);
  assign t[208] = t[207] ? x[112] : x[111];
  assign t[209] = t[74] ? x[114] : x[113];
  assign t[20] = ~(t[36] ^ t[34]);
  assign t[210] = t[27] ? x[116] : x[115];
  assign t[211] = t[238] ^ x[4];
  assign t[212] = t[239] ^ x[9];
  assign t[213] = t[240] ^ x[12];
  assign t[214] = t[241] ^ x[15];
  assign t[215] = t[242] ^ x[18];
  assign t[216] = t[243] ^ x[21];
  assign t[217] = t[244] ^ x[24];
  assign t[218] = t[245] ^ x[27];
  assign t[219] = t[246] ^ x[30];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[33];
  assign t[221] = t[248] ^ x[36];
  assign t[222] = t[249] ^ x[39];
  assign t[223] = t[250] ^ x[42];
  assign t[224] = t[251] ^ x[45];
  assign t[225] = t[252] ^ x[48];
  assign t[226] = t[253] ^ x[51];
  assign t[227] = t[254] ^ x[54];
  assign t[228] = t[255] ^ x[57];
  assign t[229] = t[256] ^ x[60];
  assign t[22] = t[21] ^ t[33];
  assign t[230] = t[257] ^ x[63];
  assign t[231] = t[258] ^ x[66];
  assign t[232] = t[259] ^ x[71];
  assign t[233] = t[260] ^ x[74];
  assign t[234] = t[261] ^ x[85];
  assign t[235] = t[262] ^ x[92];
  assign t[236] = t[263] ^ x[97];
  assign t[237] = t[264] ^ x[106];
  assign t[238] = (x[2] & x[3]);
  assign t[239] = (x[7] & x[8]);
  assign t[23] = ~(t[39] ^ t[40]);
  assign t[240] = (x[10] & x[11]);
  assign t[241] = (x[13] & x[14]);
  assign t[242] = (x[16] & x[17]);
  assign t[243] = (x[19] & x[20]);
  assign t[244] = (x[22] & x[23]);
  assign t[245] = (x[25] & x[26]);
  assign t[246] = (x[28] & x[29]);
  assign t[247] = (x[31] & x[32]);
  assign t[248] = (x[34] & x[35]);
  assign t[249] = (x[37] & x[38]);
  assign t[24] = ~(t[41] ^ t[42]);
  assign t[250] = (x[40] & x[41]);
  assign t[251] = (x[43] & x[44]);
  assign t[252] = (x[46] & x[47]);
  assign t[253] = (x[49] & x[50]);
  assign t[254] = (x[52] & x[53]);
  assign t[255] = (x[55] & x[56]);
  assign t[256] = (x[58] & x[59]);
  assign t[257] = (x[61] & x[62]);
  assign t[258] = (x[64] & x[65]);
  assign t[259] = (x[69] & x[70]);
  assign t[25] = ~(t[43] ^ t[44]);
  assign t[260] = (x[72] & x[73]);
  assign t[261] = (x[83] & x[84]);
  assign t[262] = (x[90] & x[91]);
  assign t[263] = (x[95] & x[96]);
  assign t[264] = (x[104] & x[105]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[212]);
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[214]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = t[50] ^ t[51];
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] ^ t[57];
  assign t[36] = t[58] ^ t[59];
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[38] = ~(t[62] ^ t[63]);
  assign t[39] = t[64] ^ t[65];
  assign t[3] = t[7] ? t[8] : t[211];
  assign t[40] = t[66] ^ t[67];
  assign t[41] = t[68] ^ t[54];
  assign t[42] = ~(t[37] ^ t[69]);
  assign t[43] = t[10] ^ t[70];
  assign t[44] = ~(t[61] ^ t[40]);
  assign t[45] = ~(t[71] & t[72]);
  assign t[46] = t[215] | t[73];
  assign t[47] = ~(t[74]);
  assign t[48] = ~(t[216]);
  assign t[49] = ~(t[75] & t[217]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[76] ^ t[56];
  assign t[51] = t[77] & t[78];
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] & t[82];
  assign t[54] = t[83] ^ t[84];
  assign t[55] = t[85] ^ t[86];
  assign t[56] = t[87] ? t[88] : t[218];
  assign t[57] = t[89] ^ t[90];
  assign t[58] = ~t[91];
  assign t[59] = t[92] ^ t[93];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = ~(t[94] ^ t[95]);
  assign t[61] = t[96] ^ t[97];
  assign t[62] = t[98] ^ t[99];
  assign t[63] = ~(t[69] ^ t[40]);
  assign t[64] = t[100] ^ t[66];
  assign t[65] = t[101] ^ t[102];
  assign t[66] = t[217] ^ t[103];
  assign t[67] = t[101] ^ t[86];
  assign t[68] = t[104] ^ t[105];
  assign t[69] = t[106] ^ t[107];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[108] ^ t[93];
  assign t[71] = ~(t[73] & t[109]);
  assign t[72] = ~(t[219] ^ t[110]);
  assign t[73] = ~(t[111] & t[112]);
  assign t[74] = ~(t[46]);
  assign t[75] = ~(t[220]);
  assign t[76] = t[87] ? t[113] : t[221];
  assign t[77] = ~(t[114]);
  assign t[78] = t[87] ? t[115] : t[222];
  assign t[79] = t[7] ? t[116] : t[223];
  assign t[7] = ~(t[14]);
  assign t[80] = t[7] ? t[117] : t[224];
  assign t[81] = ~(t[52] ^ t[118]);
  assign t[82] = t[96] ^ t[119];
  assign t[83] = t[120] ^ t[58];
  assign t[84] = t[92] ^ t[121];
  assign t[85] = t[122] ^ t[100];
  assign t[86] = t[123] & t[124];
  assign t[87] = ~(t[14]);
  assign t[88] = t[218] ^ t[125];
  assign t[89] = t[126] ^ t[51];
  assign t[8] = t[211] ^ t[15];
  assign t[90] = t[127] & t[128];
  assign t[91] = t[26] ? t[129] : t[225];
  assign t[92] = t[130] ^ t[131];
  assign t[93] = t[132] & t[133];
  assign t[94] = t[39] ^ t[36];
  assign t[95] = t[134] ^ t[90];
  assign t[96] = t[80] ^ t[106];
  assign t[97] = t[118] ^ t[135];
  assign t[98] = t[136] ^ t[137];
  assign t[99] = t[138] ^ t[131];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind68(x, y);
 input [116:0] x;
 output y;

 wire [273:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[140] ^ t[141];
  assign t[101] = t[142] ^ t[143];
  assign t[102] = t[128] ^ t[59];
  assign t[103] = t[41] ^ t[85];
  assign t[104] = t[144] ^ t[145];
  assign t[105] = ~t[146];
  assign t[106] = ~(t[69] ^ t[97]);
  assign t[107] = t[64] ^ t[147];
  assign t[108] = t[7] ? t[148] : t[232];
  assign t[109] = t[149] ^ t[63];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[150] & t[151];
  assign t[111] = ~(t[152] & t[153]);
  assign t[112] = t[154] ^ t[233];
  assign t[113] = ~(t[228]);
  assign t[114] = t[155] & t[154];
  assign t[115] = t[7] ? t[156] : t[234];
  assign t[116] = ~(t[82]);
  assign t[117] = t[7] ? t[157] : t[235];
  assign t[118] = t[221] ^ t[158];
  assign t[119] = t[159] & t[160];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[230] ^ t[161];
  assign t[121] = ~(t[87] ^ t[162]);
  assign t[122] = t[78] ^ t[163];
  assign t[123] = t[21] ^ t[164];
  assign t[124] = ~(t[99] ^ t[102]);
  assign t[125] = t[92] ^ t[118];
  assign t[126] = ~(t[163]);
  assign t[127] = ~(t[115]);
  assign t[128] = t[115] ^ t[82];
  assign t[129] = t[165] ^ t[144];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[166] ^ t[167];
  assign t[131] = t[231] ^ t[168];
  assign t[132] = t[7] ? t[169] : t[236];
  assign t[133] = t[26] ? t[170] : t[237];
  assign t[134] = t[26] ? t[171] : t[238];
  assign t[135] = t[172] & t[173];
  assign t[136] = t[174] & t[147];
  assign t[137] = ~(t[135] ^ t[175]);
  assign t[138] = t[176] ^ t[177];
  assign t[139] = t[96] ^ t[178];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[179] ^ t[165];
  assign t[141] = t[180] & t[181];
  assign t[142] = t[179] ^ t[144];
  assign t[143] = t[182] & t[183];
  assign t[144] = t[184] ? t[185] : t[239];
  assign t[145] = t[166] ^ t[141];
  assign t[146] = t[26] ? t[186] : t[240];
  assign t[147] = t[187];
  assign t[148] = t[232] ^ t[188];
  assign t[149] = t[189] & t[190];
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[125] ^ t[109]);
  assign t[151] = t[80] ^ t[94];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[191] | t[113]);
  assign t[154] = ~(t[241]);
  assign t[155] = ~(t[233]);
  assign t[156] = t[234] ^ t[192];
  assign t[157] = t[235] ^ t[193];
  assign t[158] = t[26] ? t[194] : t[242];
  assign t[159] = ~(t[149] ^ t[195]);
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[62] ^ t[196];
  assign t[161] = t[27] ? x[76] : x[75];
  assign t[162] = t[53] ^ t[115];
  assign t[163] = t[117] ^ t[82];
  assign t[164] = t[176] ^ t[136];
  assign t[165] = t[184] ? t[197] : t[243];
  assign t[166] = t[198] ^ t[143];
  assign t[167] = t[199] & t[200];
  assign t[168] = t[76] ? x[81] : x[80];
  assign t[169] = t[236] ^ t[201];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[237] ^ t[202];
  assign t[171] = t[238] ^ t[203];
  assign t[172] = ~(t[177]);
  assign t[173] = ~(t[105]);
  assign t[174] = ~(t[95]);
  assign t[175] = t[64] ^ t[105];
  assign t[176] = t[105] ^ t[96];
  assign t[177] = t[147] ^ t[95];
  assign t[178] = t[97] ^ t[70];
  assign t[179] = t[184] ? t[204] : t[244];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = ~(t[140] ^ t[166]);
  assign t[181] = t[129] ^ t[183];
  assign t[182] = ~(t[165]);
  assign t[183] = t[184] ? t[205] : t[245];
  assign t[184] = ~(t[14]);
  assign t[185] = t[239] ^ t[206];
  assign t[186] = t[240] ^ t[207];
  assign t[187] = t[26] ? t[208] : t[246];
  assign t[188] = t[76] ? x[92] : x[91];
  assign t[189] = ~(t[196]);
  assign t[18] = ~(t[32] ^ t[33]);
  assign t[190] = ~(t[92]);
  assign t[191] = ~(t[225]);
  assign t[192] = t[27] ? x[94] : x[93];
  assign t[193] = t[27] ? x[96] : x[95];
  assign t[194] = t[242] ^ t[209];
  assign t[195] = t[80] ^ t[92];
  assign t[196] = t[94] ^ t[118];
  assign t[197] = t[243] ^ t[210];
  assign t[198] = t[211] & t[212];
  assign t[199] = ~(t[198] ^ t[213]);
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[142] ^ t[214];
  assign t[201] = t[215] ? x[98] : x[97];
  assign t[202] = t[215] ? x[100] : x[99];
  assign t[203] = t[76] ? x[102] : x[101];
  assign t[204] = t[244] ^ t[216];
  assign t[205] = t[245] ^ t[217];
  assign t[206] = t[218] ? x[104] : x[103];
  assign t[207] = t[76] ? x[106] : x[105];
  assign t[208] = t[246] ^ t[219];
  assign t[209] = t[215] ? x[108] : x[107];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[218] ? x[110] : x[109];
  assign t[211] = ~(t[214]);
  assign t[212] = ~(t[179]);
  assign t[213] = t[129] ^ t[179];
  assign t[214] = t[183] ^ t[165];
  assign t[215] = ~(t[48]);
  assign t[216] = t[218] ? x[112] : x[111];
  assign t[217] = t[218] ? x[114] : x[113];
  assign t[218] = ~(t[48]);
  assign t[219] = t[27] ? x[116] : x[115];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[4];
  assign t[221] = t[248] ^ x[9];
  assign t[222] = t[249] ^ x[12];
  assign t[223] = t[250] ^ x[15];
  assign t[224] = t[251] ^ x[18];
  assign t[225] = t[252] ^ x[21];
  assign t[226] = t[253] ^ x[24];
  assign t[227] = t[254] ^ x[27];
  assign t[228] = t[255] ^ x[30];
  assign t[229] = t[256] ^ x[33];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[36];
  assign t[231] = t[258] ^ x[41];
  assign t[232] = t[259] ^ x[44];
  assign t[233] = t[260] ^ x[47];
  assign t[234] = t[261] ^ x[50];
  assign t[235] = t[262] ^ x[53];
  assign t[236] = t[263] ^ x[56];
  assign t[237] = t[264] ^ x[59];
  assign t[238] = t[265] ^ x[62];
  assign t[239] = t[266] ^ x[65];
  assign t[23] = ~(t[42] ^ t[20]);
  assign t[240] = t[267] ^ x[68];
  assign t[241] = t[268] ^ x[71];
  assign t[242] = t[269] ^ x[74];
  assign t[243] = t[270] ^ x[79];
  assign t[244] = t[271] ^ x[84];
  assign t[245] = t[272] ^ x[87];
  assign t[246] = t[273] ^ x[90];
  assign t[247] = (x[2] & x[3]);
  assign t[248] = (x[7] & x[8]);
  assign t[249] = (x[10] & x[11]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (x[13] & x[14]);
  assign t[251] = (x[16] & x[17]);
  assign t[252] = (x[19] & x[20]);
  assign t[253] = (x[22] & x[23]);
  assign t[254] = (x[25] & x[26]);
  assign t[255] = (x[28] & x[29]);
  assign t[256] = (x[31] & x[32]);
  assign t[257] = (x[34] & x[35]);
  assign t[258] = (x[39] & x[40]);
  assign t[259] = (x[42] & x[43]);
  assign t[25] = ~(t[34] ^ t[45]);
  assign t[260] = (x[45] & x[46]);
  assign t[261] = (x[48] & x[49]);
  assign t[262] = (x[51] & x[52]);
  assign t[263] = (x[54] & x[55]);
  assign t[264] = (x[57] & x[58]);
  assign t[265] = (x[60] & x[61]);
  assign t[266] = (x[63] & x[64]);
  assign t[267] = (x[66] & x[67]);
  assign t[268] = (x[69] & x[70]);
  assign t[269] = (x[72] & x[73]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[270] = (x[77] & x[78]);
  assign t[271] = (x[82] & x[83]);
  assign t[272] = (x[85] & x[86]);
  assign t[273] = (x[88] & x[89]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[221]);
  assign t[29] = ~(t[222]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[223]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[51] ^ t[13];
  assign t[33] = ~(t[52] ^ t[42]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] ^ t[56]);
  assign t[36] = t[7] ? t[57] : t[224];
  assign t[37] = t[58] ^ t[59];
  assign t[38] = t[60] ^ t[61];
  assign t[39] = ~(t[40] ^ t[45]);
  assign t[3] = t[7] ? t[8] : t[220];
  assign t[40] = t[62] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = ~(t[66] ^ t[34]);
  assign t[43] = ~(t[67] ^ t[68]);
  assign t[44] = t[69] ^ t[70];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = ~(t[73] & t[74]);
  assign t[47] = t[225] | t[75];
  assign t[48] = ~(t[76]);
  assign t[49] = ~(t[226]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[77] & t[227]);
  assign t[51] = t[78] ^ t[79];
  assign t[52] = t[80] ^ t[81];
  assign t[53] = t[82] ^ t[36];
  assign t[54] = t[58] ^ t[83];
  assign t[55] = t[84] ^ t[43];
  assign t[56] = ~(t[20] ^ t[85]);
  assign t[57] = t[224] ^ t[86];
  assign t[58] = t[87] ^ t[79];
  assign t[59] = t[88] & t[89];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[20] ^ t[51];
  assign t[61] = ~(t[90] ^ t[91]);
  assign t[62] = t[92] ^ t[71];
  assign t[63] = t[93] & t[94];
  assign t[64] = t[95] ^ t[96];
  assign t[65] = t[97] ^ t[98];
  assign t[66] = ~(t[99] ^ t[100]);
  assign t[67] = t[101] ^ t[102];
  assign t[68] = ~(t[103] ^ t[104]);
  assign t[69] = t[105] ^ t[95];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[106] & t[107];
  assign t[71] = t[227] ^ t[108];
  assign t[72] = t[109] ^ t[110];
  assign t[73] = ~(t[75] & t[111]);
  assign t[74] = ~(t[228] ^ t[112]);
  assign t[75] = ~(t[113] & t[114]);
  assign t[76] = ~(t[47]);
  assign t[77] = ~(t[229]);
  assign t[78] = t[115] ^ t[36];
  assign t[79] = t[116] & t[117];
  assign t[7] = ~(t[14]);
  assign t[80] = t[118] ^ t[71];
  assign t[81] = t[109] ^ t[119];
  assign t[82] = t[7] ? t[120] : t[230];
  assign t[83] = t[121] & t[122];
  assign t[84] = ~(t[123] ^ t[124]);
  assign t[85] = t[125] ^ t[110];
  assign t[86] = t[27] ? x[38] : x[37];
  assign t[87] = t[126] & t[127];
  assign t[88] = ~(t[128] ^ t[58]);
  assign t[89] = t[53] ^ t[117];
  assign t[8] = t[220] ^ t[15];
  assign t[90] = ~(t[44] ^ t[104]);
  assign t[91] = t[129] ^ t[130];
  assign t[92] = t[7] ? t[131] : t[231];
  assign t[93] = ~(t[118]);
  assign t[94] = t[222] ^ t[132];
  assign t[95] = t[133];
  assign t[96] = ~t[134];
  assign t[97] = t[135] ^ t[136];
  assign t[98] = t[137] & t[138];
  assign t[99] = t[52] ^ t[139];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind69(x, y);
 input [116:0] x;
 output y;

 wire [264:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[26] ? t[142] : t[225];
  assign t[101] = t[26] ? t[143] : t[226];
  assign t[102] = t[26] ? t[144] : t[227];
  assign t[103] = t[27] ? x[56] : x[55];
  assign t[104] = ~(t[116] ^ t[56]);
  assign t[105] = t[34] ^ t[126];
  assign t[106] = t[222] ^ t[145];
  assign t[107] = t[146] & t[147];
  assign t[108] = t[148] & t[149];
  assign t[109] = ~(t[92] ^ t[71]);
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = t[150] ^ t[149];
  assign t[111] = ~(t[151] & t[152]);
  assign t[112] = t[153] ^ t[228];
  assign t[113] = ~(t[223]);
  assign t[114] = t[154] & t[153];
  assign t[115] = t[155] ^ t[61];
  assign t[116] = t[156] ^ t[55];
  assign t[117] = t[121] ^ t[157];
  assign t[118] = t[62] ^ t[158];
  assign t[119] = t[26] ? t[159] : t[229];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[160] ^ t[41];
  assign t[121] = t[82] ^ t[65];
  assign t[122] = t[27] ? x[64] : x[63];
  assign t[123] = ~(t[129]);
  assign t[124] = ~(t[156]);
  assign t[125] = ~(t[55]);
  assign t[126] = t[7] ? t[161] : t[230];
  assign t[127] = t[34] ^ t[156];
  assign t[128] = t[156] ^ t[42];
  assign t[129] = t[126] ^ t[55];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = ~(t[162] ^ t[163]);
  assign t[131] = t[164] ^ t[165];
  assign t[132] = t[7] ? t[166] : t[231];
  assign t[133] = t[212] ^ t[167];
  assign t[134] = t[168] ? x[72] : x[71];
  assign t[135] = t[168] ? x[74] : x[73];
  assign t[136] = ~(t[141]);
  assign t[137] = ~(t[155]);
  assign t[138] = ~(t[60]);
  assign t[139] = t[93] ? t[169] : t[232];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[38] ^ t[155];
  assign t[141] = t[139] ^ t[60];
  assign t[142] = t[225] ^ t[170];
  assign t[143] = t[226] ^ t[171];
  assign t[144] = t[227] ^ t[172];
  assign t[145] = t[76] ? x[79] : x[78];
  assign t[146] = ~(t[173]);
  assign t[147] = ~(t[132]);
  assign t[148] = ~(t[133]);
  assign t[149] = t[213] ^ t[174];
  assign t[14] = ~(t[26]);
  assign t[150] = t[133] ^ t[44];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[175] | t[113]);
  assign t[153] = ~(t[233]);
  assign t[154] = ~(t[228]);
  assign t[155] = t[93] ? t[176] : t[234];
  assign t[156] = t[7] ? t[177] : t[235];
  assign t[157] = t[120] ^ t[178];
  assign t[158] = t[179] & t[180];
  assign t[159] = t[229] ^ t[181];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[182] & t[183];
  assign t[161] = t[230] ^ t[184];
  assign t[162] = t[185] ^ t[186];
  assign t[163] = ~(t[187] ^ t[25]);
  assign t[164] = t[150] ^ t[188];
  assign t[165] = t[65] ^ t[189];
  assign t[166] = t[231] ^ t[190];
  assign t[167] = t[26] ? t[191] : t[236];
  assign t[168] = ~(t[48]);
  assign t[169] = t[232] ^ t[192];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[76] ? x[93] : x[92];
  assign t[171] = t[76] ? x[95] : x[94];
  assign t[172] = t[27] ? x[97] : x[96];
  assign t[173] = t[149] ^ t[133];
  assign t[174] = t[7] ? t[193] : t[237];
  assign t[175] = ~(t[217]);
  assign t[176] = t[234] ^ t[194];
  assign t[177] = t[235] ^ t[195];
  assign t[178] = t[196] & t[197];
  assign t[179] = ~(t[198] ^ t[62]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[38] ^ t[139];
  assign t[181] = t[199] ? x[102] : x[101];
  assign t[182] = ~(t[200]);
  assign t[183] = ~(t[64]);
  assign t[184] = t[27] ? x[104] : x[103];
  assign t[185] = t[24] ^ t[201];
  assign t[186] = ~(t[202] ^ t[22]);
  assign t[187] = t[203] ^ t[108];
  assign t[188] = t[71] ^ t[204];
  assign t[189] = t[120] ^ t[54];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[76] ? x[106] : x[105];
  assign t[191] = t[236] ^ t[205];
  assign t[192] = t[168] ? x[108] : x[107];
  assign t[193] = t[237] ^ t[206];
  assign t[194] = t[168] ? x[110] : x[109];
  assign t[195] = t[27] ? x[112] : x[111];
  assign t[196] = ~(t[160] ^ t[207]);
  assign t[197] = t[40] ^ t[200];
  assign t[198] = t[155] ^ t[60];
  assign t[199] = ~(t[48]);
  assign t[19] = ~(t[20] ^ t[25]);
  assign t[1] = ~(t[4]);
  assign t[200] = t[67] ^ t[82];
  assign t[201] = t[128] ^ t[87];
  assign t[202] = ~(t[33] ^ t[81]);
  assign t[203] = t[132] ^ t[44];
  assign t[204] = t[208] & t[209];
  assign t[205] = t[199] ? x[114] : x[113];
  assign t[206] = t[199] ? x[116] : x[115];
  assign t[207] = t[121] ^ t[64];
  assign t[208] = ~(t[107] ^ t[210]);
  assign t[209] = t[203] ^ t[173];
  assign t[20] = t[34] ^ t[35];
  assign t[210] = t[150] ^ t[132];
  assign t[211] = t[238] ^ x[4];
  assign t[212] = t[239] ^ x[9];
  assign t[213] = t[240] ^ x[12];
  assign t[214] = t[241] ^ x[15];
  assign t[215] = t[242] ^ x[18];
  assign t[216] = t[243] ^ x[21];
  assign t[217] = t[244] ^ x[24];
  assign t[218] = t[245] ^ x[27];
  assign t[219] = t[246] ^ x[30];
  assign t[21] = ~(t[36] ^ t[37]);
  assign t[220] = t[247] ^ x[33];
  assign t[221] = t[248] ^ x[36];
  assign t[222] = t[249] ^ x[39];
  assign t[223] = t[250] ^ x[42];
  assign t[224] = t[251] ^ x[45];
  assign t[225] = t[252] ^ x[48];
  assign t[226] = t[253] ^ x[51];
  assign t[227] = t[254] ^ x[54];
  assign t[228] = t[255] ^ x[59];
  assign t[229] = t[256] ^ x[62];
  assign t[22] = t[38] ^ t[39];
  assign t[230] = t[257] ^ x[67];
  assign t[231] = t[258] ^ x[70];
  assign t[232] = t[259] ^ x[77];
  assign t[233] = t[260] ^ x[82];
  assign t[234] = t[261] ^ x[85];
  assign t[235] = t[262] ^ x[88];
  assign t[236] = t[263] ^ x[91];
  assign t[237] = t[264] ^ x[100];
  assign t[238] = (x[2] & x[3]);
  assign t[239] = (x[7] & x[8]);
  assign t[23] = t[40] ^ t[41];
  assign t[240] = (x[10] & x[11]);
  assign t[241] = (x[13] & x[14]);
  assign t[242] = (x[16] & x[17]);
  assign t[243] = (x[19] & x[20]);
  assign t[244] = (x[22] & x[23]);
  assign t[245] = (x[25] & x[26]);
  assign t[246] = (x[28] & x[29]);
  assign t[247] = (x[31] & x[32]);
  assign t[248] = (x[34] & x[35]);
  assign t[249] = (x[37] & x[38]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (x[40] & x[41]);
  assign t[251] = (x[43] & x[44]);
  assign t[252] = (x[46] & x[47]);
  assign t[253] = (x[49] & x[50]);
  assign t[254] = (x[52] & x[53]);
  assign t[255] = (x[57] & x[58]);
  assign t[256] = (x[60] & x[61]);
  assign t[257] = (x[65] & x[66]);
  assign t[258] = (x[68] & x[69]);
  assign t[259] = (x[75] & x[76]);
  assign t[25] = t[44] ^ t[45];
  assign t[260] = (x[80] & x[81]);
  assign t[261] = (x[83] & x[84]);
  assign t[262] = (x[86] & x[87]);
  assign t[263] = (x[89] & x[90]);
  assign t[264] = (x[98] & x[99]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[212]);
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[214]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = ~(t[51] ^ t[52]);
  assign t[33] = t[53] ^ t[54];
  assign t[34] = t[55] ^ t[42];
  assign t[35] = t[56] ^ t[57];
  assign t[36] = t[58] ^ t[32];
  assign t[37] = ~(t[24] ^ t[59]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[62] ^ t[63];
  assign t[3] = t[7] ? t[8] : t[211];
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[66] & t[67];
  assign t[42] = t[7] ? t[68] : t[215];
  assign t[43] = t[56] ^ t[69];
  assign t[44] = t[216] ^ t[70];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = ~(t[73] & t[74]);
  assign t[47] = t[217] | t[75];
  assign t[48] = ~(t[76]);
  assign t[49] = ~(t[218]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[77] & t[216]);
  assign t[51] = t[78] ^ t[79];
  assign t[52] = ~(t[80] ^ t[81]);
  assign t[53] = t[64] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[7] ? t[85] : t[219];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] & t[89];
  assign t[58] = ~(t[90] ^ t[91]);
  assign t[59] = t[92] ^ t[72];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[93] ? t[94] : t[220];
  assign t[61] = t[93] ? t[95] : t[221];
  assign t[62] = t[96] ^ t[97];
  assign t[63] = t[98] & t[99];
  assign t[64] = ~t[100];
  assign t[65] = ~t[101];
  assign t[66] = ~(t[82]);
  assign t[67] = t[102];
  assign t[68] = t[215] ^ t[103];
  assign t[69] = t[104] & t[105];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[7] ? t[106] : t[222];
  assign t[71] = t[107] ^ t[108];
  assign t[72] = t[109] & t[110];
  assign t[73] = ~(t[75] & t[111]);
  assign t[74] = ~(t[223] ^ t[112]);
  assign t[75] = ~(t[113] & t[114]);
  assign t[76] = ~(t[47]);
  assign t[77] = ~(t[224]);
  assign t[78] = t[115] ^ t[97];
  assign t[79] = t[116] ^ t[69];
  assign t[7] = ~(t[14]);
  assign t[80] = t[117] ^ t[59];
  assign t[81] = t[61] ^ t[118];
  assign t[82] = t[119];
  assign t[83] = ~(t[53] ^ t[120]);
  assign t[84] = t[121] ^ t[67];
  assign t[85] = t[219] ^ t[122];
  assign t[86] = t[123] & t[124];
  assign t[87] = t[125] & t[126];
  assign t[88] = ~(t[86] ^ t[127]);
  assign t[89] = t[128] ^ t[129];
  assign t[8] = t[211] ^ t[15];
  assign t[90] = t[130] ^ t[23];
  assign t[91] = ~(t[131] ^ t[79]);
  assign t[92] = t[132] ^ t[133];
  assign t[93] = ~(t[14]);
  assign t[94] = t[220] ^ t[134];
  assign t[95] = t[221] ^ t[135];
  assign t[96] = t[136] & t[137];
  assign t[97] = t[138] & t[139];
  assign t[98] = ~(t[96] ^ t[140]);
  assign t[99] = t[115] ^ t[141];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind70(x, y);
 input [116:0] x;
 output y;

 wire [262:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[27] ? x[56] : x[55];
  assign t[101] = t[217] ^ t[142];
  assign t[102] = t[7] ? t[143] : t[226];
  assign t[103] = ~(t[144] & t[145]);
  assign t[104] = t[146] ^ t[227];
  assign t[105] = ~(t[219]);
  assign t[106] = t[147] & t[146];
  assign t[107] = t[86] ^ t[126];
  assign t[108] = t[148] & t[149];
  assign t[109] = t[131] ? t[150] : t[228];
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = t[111] ^ t[61];
  assign t[111] = t[151] ^ t[152];
  assign t[112] = t[153] & t[154];
  assign t[113] = t[220] ^ t[155];
  assign t[114] = t[156] ^ t[58];
  assign t[115] = t[126] ^ t[77];
  assign t[116] = t[114] ^ t[157];
  assign t[117] = t[158] ^ t[128];
  assign t[118] = t[159] & t[160];
  assign t[119] = t[62] ^ t[161];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[140] ^ t[97];
  assign t[121] = t[158] ^ t[123];
  assign t[122] = t[162] & t[163];
  assign t[123] = t[164];
  assign t[124] = t[129] ^ t[118];
  assign t[125] = t[221] ^ t[165];
  assign t[126] = t[7] ? t[166] : t[229];
  assign t[127] = t[222] ^ t[167];
  assign t[128] = ~t[168];
  assign t[129] = t[169] ^ t[122];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[170] & t[171];
  assign t[131] = ~(t[14]);
  assign t[132] = t[223] ^ t[172];
  assign t[133] = t[224] ^ t[173];
  assign t[134] = t[131] ? t[174] : t[230];
  assign t[135] = t[225] ^ t[175];
  assign t[136] = ~(t[141]);
  assign t[137] = ~(t[41]);
  assign t[138] = ~(t[42]);
  assign t[139] = t[39] ^ t[41];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[41] ^ t[62];
  assign t[141] = t[67] ^ t[42];
  assign t[142] = t[27] ? x[73] : x[72];
  assign t[143] = t[226] ^ t[176];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[177] | t[105]);
  assign t[146] = ~(t[231]);
  assign t[147] = ~(t[227]);
  assign t[148] = ~(t[107] ^ t[114]);
  assign t[149] = t[115] ^ t[88];
  assign t[14] = ~(t[26]);
  assign t[150] = t[228] ^ t[178];
  assign t[151] = t[179] & t[180];
  assign t[152] = t[181] & t[134];
  assign t[153] = ~(t[151] ^ t[182]);
  assign t[154] = t[183] ^ t[184];
  assign t[155] = t[71] ? x[78] : x[77];
  assign t[156] = t[185] & t[186];
  assign t[157] = t[187] & t[188];
  assign t[158] = t[189];
  assign t[159] = ~(t[117] ^ t[129]);
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[89] ^ t[163];
  assign t[161] = t[63] ^ t[25];
  assign t[162] = ~(t[128]);
  assign t[163] = t[190];
  assign t[164] = t[7] ? t[191] : t[232];
  assign t[165] = t[192] ? x[83] : x[82];
  assign t[166] = t[229] ^ t[193];
  assign t[167] = t[192] ? x[85] : x[84];
  assign t[168] = t[7] ? t[194] : t[233];
  assign t[169] = t[195] & t[196];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = ~(t[169] ^ t[197]);
  assign t[171] = t[121] ^ t[198];
  assign t[172] = t[199] ? x[90] : x[89];
  assign t[173] = t[199] ? x[92] : x[91];
  assign t[174] = t[230] ^ t[200];
  assign t[175] = t[27] ? x[94] : x[93];
  assign t[176] = t[27] ? x[96] : x[95];
  assign t[177] = ~(t[214]);
  assign t[178] = t[199] ? x[98] : x[97];
  assign t[179] = ~(t[184]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = ~(t[91]);
  assign t[181] = ~(t[92]);
  assign t[182] = t[75] ^ t[91];
  assign t[183] = t[91] ^ t[109];
  assign t[184] = t[134] ^ t[92];
  assign t[185] = ~(t[201]);
  assign t[186] = ~(t[86]);
  assign t[187] = ~(t[156] ^ t[202]);
  assign t[188] = t[57] ^ t[201];
  assign t[189] = t[7] ? t[203] : t[234];
  assign t[18] = ~(t[23] ^ t[32]);
  assign t[190] = t[7] ? t[204] : t[235];
  assign t[191] = t[232] ^ t[205];
  assign t[192] = ~(t[47]);
  assign t[193] = t[192] ? x[106] : x[105];
  assign t[194] = t[233] ^ t[206];
  assign t[195] = ~(t[198]);
  assign t[196] = ~(t[158]);
  assign t[197] = t[89] ^ t[158];
  assign t[198] = t[163] ^ t[128];
  assign t[199] = ~(t[47]);
  assign t[19] = ~(t[33] ^ t[34]);
  assign t[1] = ~(t[4]);
  assign t[200] = t[199] ? x[108] : x[107];
  assign t[201] = t[88] ^ t[126];
  assign t[202] = t[115] ^ t[86];
  assign t[203] = t[234] ^ t[207];
  assign t[204] = t[235] ^ t[208];
  assign t[205] = t[71] ? x[110] : x[109];
  assign t[206] = t[27] ? x[112] : x[111];
  assign t[207] = t[71] ? x[114] : x[113];
  assign t[208] = t[71] ? x[116] : x[115];
  assign t[209] = t[236] ^ x[4];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[237] ^ x[9];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[37] ^ t[13]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[59];
  assign t[227] = t[254] ^ x[62];
  assign t[228] = t[255] ^ x[65];
  assign t[229] = t[256] ^ x[68];
  assign t[22] = ~(t[37] ^ t[38]);
  assign t[230] = t[257] ^ x[71];
  assign t[231] = t[258] ^ x[76];
  assign t[232] = t[259] ^ x[81];
  assign t[233] = t[260] ^ x[88];
  assign t[234] = t[261] ^ x[101];
  assign t[235] = t[262] ^ x[104];
  assign t[236] = (x[2] & x[3]);
  assign t[237] = (x[7] & x[8]);
  assign t[238] = (x[10] & x[11]);
  assign t[239] = (x[13] & x[14]);
  assign t[23] = t[39] ^ t[40];
  assign t[240] = (x[16] & x[17]);
  assign t[241] = (x[19] & x[20]);
  assign t[242] = (x[22] & x[23]);
  assign t[243] = (x[25] & x[26]);
  assign t[244] = (x[28] & x[29]);
  assign t[245] = (x[31] & x[32]);
  assign t[246] = (x[34] & x[35]);
  assign t[247] = (x[37] & x[38]);
  assign t[248] = (x[40] & x[41]);
  assign t[249] = (x[43] & x[44]);
  assign t[24] = t[41] ^ t[42];
  assign t[250] = (x[46] & x[47]);
  assign t[251] = (x[49] & x[50]);
  assign t[252] = (x[52] & x[53]);
  assign t[253] = (x[57] & x[58]);
  assign t[254] = (x[60] & x[61]);
  assign t[255] = (x[63] & x[64]);
  assign t[256] = (x[66] & x[67]);
  assign t[257] = (x[69] & x[70]);
  assign t[258] = (x[74] & x[75]);
  assign t[259] = (x[79] & x[80]);
  assign t[25] = t[43] & t[44];
  assign t[260] = (x[86] & x[87]);
  assign t[261] = (x[99] & x[100]);
  assign t[262] = (x[102] & x[103]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[210]);
  assign t[29] = ~(t[211]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[212]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = ~(t[50] ^ t[51]);
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[34] = t[12] ^ t[54];
  assign t[35] = ~(t[55] ^ t[56]);
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ t[52];
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[42] ^ t[62];
  assign t[3] = t[7] ? t[8] : t[209];
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[7] ? t[65] : t[213];
  assign t[42] = t[212] ^ t[66];
  assign t[43] = ~(t[24] ^ t[63]);
  assign t[44] = t[39] ^ t[67];
  assign t[45] = ~(t[68] & t[69]);
  assign t[46] = t[214] | t[70];
  assign t[47] = ~(t[71]);
  assign t[48] = ~(t[215]);
  assign t[49] = ~(t[72] & t[216]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[73] ^ t[74]);
  assign t[51] = t[75] ^ t[76];
  assign t[52] = t[77] ^ t[78];
  assign t[53] = t[79] ^ t[80];
  assign t[54] = ~(t[81] ^ t[82]);
  assign t[55] = t[83] ^ t[32];
  assign t[56] = ~(t[84] ^ t[85]);
  assign t[57] = t[86] ^ t[77];
  assign t[58] = t[87] & t[88];
  assign t[59] = t[89] ^ t[90];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[91] ^ t[92];
  assign t[61] = t[93] & t[94];
  assign t[62] = t[215] ^ t[95];
  assign t[63] = t[96] ^ t[97];
  assign t[64] = t[98] & t[99];
  assign t[65] = t[213] ^ t[100];
  assign t[66] = t[7] ? t[101] : t[217];
  assign t[67] = t[218] ^ t[102];
  assign t[68] = ~(t[70] & t[103]);
  assign t[69] = ~(t[219] ^ t[104]);
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[105] & t[106]);
  assign t[71] = ~(t[46]);
  assign t[72] = ~(t[218]);
  assign t[73] = t[107] ^ t[108];
  assign t[74] = t[109] ^ t[110];
  assign t[75] = t[92] ^ t[109];
  assign t[76] = t[111] ^ t[112];
  assign t[77] = t[7] ? t[113] : t[220];
  assign t[78] = t[114] ^ t[108];
  assign t[79] = t[115] ^ t[116];
  assign t[7] = ~(t[14]);
  assign t[80] = t[117] ^ t[118];
  assign t[81] = t[51] ^ t[36];
  assign t[82] = ~(t[119] ^ t[85]);
  assign t[83] = t[119] ^ t[120];
  assign t[84] = t[121] ^ t[122];
  assign t[85] = t[123] ^ t[124];
  assign t[86] = t[7] ? t[125] : t[221];
  assign t[87] = ~(t[126]);
  assign t[88] = t[7] ? t[127] : t[222];
  assign t[89] = t[128] ^ t[123];
  assign t[8] = t[209] ^ t[15];
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[131] ? t[132] : t[223];
  assign t[92] = t[131] ? t[133] : t[224];
  assign t[93] = ~(t[60] ^ t[111]);
  assign t[94] = t[75] ^ t[134];
  assign t[95] = t[7] ? t[135] : t[225];
  assign t[96] = t[136] & t[137];
  assign t[97] = t[138] & t[67];
  assign t[98] = ~(t[96] ^ t[139]);
  assign t[99] = t[140] ^ t[141];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind71(x, y);
 input [116:0] x;
 output y;

 wire [264:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~t[139];
  assign t[101] = t[140] ^ t[105];
  assign t[102] = t[141] & t[142];
  assign t[103] = t[7] ? t[143] : t[225];
  assign t[104] = t[122] ^ t[66];
  assign t[105] = t[144] & t[145];
  assign t[106] = t[216] ^ t[146];
  assign t[107] = t[118] ^ t[53];
  assign t[108] = t[147] ^ t[120];
  assign t[109] = ~(t[148] & t[149]);
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = t[150] ^ t[226];
  assign t[111] = ~(t[220]);
  assign t[112] = t[151] & t[150];
  assign t[113] = t[222] ^ t[152];
  assign t[114] = t[87] ? t[153] : t[227];
  assign t[115] = t[223] ^ t[154];
  assign t[116] = t[224] ^ t[155];
  assign t[117] = t[7] ? t[156] : t[228];
  assign t[118] = t[157] ^ t[158];
  assign t[119] = t[221] ^ t[159];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[7] ? t[160] : t[229];
  assign t[121] = t[161] & t[162];
  assign t[122] = t[163];
  assign t[123] = ~(t[85] ^ t[101]);
  assign t[124] = t[64] ^ t[145];
  assign t[125] = t[164] ? x[62] : x[61];
  assign t[126] = t[165] & t[166];
  assign t[127] = ~(t[134] ^ t[89]);
  assign t[128] = t[136] ^ t[78];
  assign t[129] = t[74] ? x[64] : x[63];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[167] & t[168];
  assign t[131] = t[169] & t[170];
  assign t[132] = ~(t[108] ^ t[92]);
  assign t[133] = t[83] ^ t[170];
  assign t[134] = t[76] ^ t[114];
  assign t[135] = t[171] & t[172];
  assign t[136] = t[114] ^ t[56];
  assign t[137] = t[89] ^ t[173];
  assign t[138] = t[147] ^ t[58];
  assign t[139] = t[7] ? t[174] : t[230];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[175] & t[176];
  assign t[141] = ~(t[140] ^ t[177]);
  assign t[142] = t[104] ^ t[178];
  assign t[143] = t[225] ^ t[179];
  assign t[144] = ~(t[100]);
  assign t[145] = t[180];
  assign t[146] = t[7] ? t[181] : t[231];
  assign t[147] = t[7] ? t[182] : t[232];
  assign t[148] = ~(t[151] | t[150]);
  assign t[149] = ~(t[183] | t[111]);
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[233]);
  assign t[151] = ~(t[226]);
  assign t[152] = t[164] ? x[78] : x[77];
  assign t[153] = t[227] ^ t[184];
  assign t[154] = t[164] ? x[80] : x[79];
  assign t[155] = t[27] ? x[82] : x[81];
  assign t[156] = t[228] ^ t[185];
  assign t[157] = t[186] & t[187];
  assign t[158] = t[188] & t[119];
  assign t[159] = t[7] ? t[189] : t[234];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[229] ^ t[190];
  assign t[161] = ~(t[130] ^ t[191]);
  assign t[162] = t[138] ^ t[192];
  assign t[163] = t[7] ? t[193] : t[235];
  assign t[164] = ~(t[47]);
  assign t[165] = ~(t[194]);
  assign t[166] = ~(t[76]);
  assign t[167] = ~(t[192]);
  assign t[168] = ~(t[147]);
  assign t[169] = ~(t[120]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[7] ? t[195] : t[236];
  assign t[171] = ~(t[157] ^ t[196]);
  assign t[172] = t[197] ^ t[198];
  assign t[173] = t[199] & t[200];
  assign t[174] = t[230] ^ t[201];
  assign t[175] = ~(t[178]);
  assign t[176] = ~(t[122]);
  assign t[177] = t[64] ^ t[122];
  assign t[178] = t[145] ^ t[100];
  assign t[179] = t[74] ? x[93] : x[92];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[7] ? t[202] : t[237];
  assign t[181] = t[231] ^ t[203];
  assign t[182] = t[232] ^ t[204];
  assign t[183] = ~(t[215]);
  assign t[184] = t[164] ? x[98] : x[97];
  assign t[185] = t[27] ? x[100] : x[99];
  assign t[186] = ~(t[198]);
  assign t[187] = ~(t[79]);
  assign t[188] = ~(t[80]);
  assign t[189] = t[234] ^ t[205];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[206] ? x[102] : x[101];
  assign t[191] = t[83] ^ t[147];
  assign t[192] = t[170] ^ t[120];
  assign t[193] = t[235] ^ t[207];
  assign t[194] = t[78] ^ t[114];
  assign t[195] = t[236] ^ t[208];
  assign t[196] = t[96] ^ t[79];
  assign t[197] = t[79] ^ t[106];
  assign t[198] = t[119] ^ t[80];
  assign t[199] = ~(t[126] ^ t[209]);
  assign t[19] = ~(t[34] ^ t[35]);
  assign t[1] = ~(t[4]);
  assign t[200] = t[50] ^ t[194];
  assign t[201] = t[27] ? x[104] : x[103];
  assign t[202] = t[237] ^ t[210];
  assign t[203] = t[27] ? x[106] : x[105];
  assign t[204] = t[206] ? x[108] : x[107];
  assign t[205] = t[27] ? x[110] : x[109];
  assign t[206] = ~(t[47]);
  assign t[207] = t[74] ? x[112] : x[111];
  assign t[208] = t[206] ? x[114] : x[113];
  assign t[209] = t[136] ^ t[76];
  assign t[20] = ~(t[36] ^ t[34]);
  assign t[210] = t[74] ? x[116] : x[115];
  assign t[211] = t[238] ^ x[4];
  assign t[212] = t[239] ^ x[9];
  assign t[213] = t[240] ^ x[12];
  assign t[214] = t[241] ^ x[15];
  assign t[215] = t[242] ^ x[18];
  assign t[216] = t[243] ^ x[21];
  assign t[217] = t[244] ^ x[24];
  assign t[218] = t[245] ^ x[27];
  assign t[219] = t[246] ^ x[30];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[33];
  assign t[221] = t[248] ^ x[36];
  assign t[222] = t[249] ^ x[39];
  assign t[223] = t[250] ^ x[42];
  assign t[224] = t[251] ^ x[45];
  assign t[225] = t[252] ^ x[48];
  assign t[226] = t[253] ^ x[51];
  assign t[227] = t[254] ^ x[54];
  assign t[228] = t[255] ^ x[57];
  assign t[229] = t[256] ^ x[60];
  assign t[22] = t[21] ^ t[33];
  assign t[230] = t[257] ^ x[67];
  assign t[231] = t[258] ^ x[70];
  assign t[232] = t[259] ^ x[73];
  assign t[233] = t[260] ^ x[76];
  assign t[234] = t[261] ^ x[85];
  assign t[235] = t[262] ^ x[88];
  assign t[236] = t[263] ^ x[91];
  assign t[237] = t[264] ^ x[96];
  assign t[238] = (x[2] & x[3]);
  assign t[239] = (x[7] & x[8]);
  assign t[23] = ~(t[39] ^ t[40]);
  assign t[240] = (x[10] & x[11]);
  assign t[241] = (x[13] & x[14]);
  assign t[242] = (x[16] & x[17]);
  assign t[243] = (x[19] & x[20]);
  assign t[244] = (x[22] & x[23]);
  assign t[245] = (x[25] & x[26]);
  assign t[246] = (x[28] & x[29]);
  assign t[247] = (x[31] & x[32]);
  assign t[248] = (x[34] & x[35]);
  assign t[249] = (x[37] & x[38]);
  assign t[24] = ~(t[41] ^ t[42]);
  assign t[250] = (x[40] & x[41]);
  assign t[251] = (x[43] & x[44]);
  assign t[252] = (x[46] & x[47]);
  assign t[253] = (x[49] & x[50]);
  assign t[254] = (x[52] & x[53]);
  assign t[255] = (x[55] & x[56]);
  assign t[256] = (x[58] & x[59]);
  assign t[257] = (x[65] & x[66]);
  assign t[258] = (x[68] & x[69]);
  assign t[259] = (x[71] & x[72]);
  assign t[25] = ~(t[43] ^ t[44]);
  assign t[260] = (x[74] & x[75]);
  assign t[261] = (x[83] & x[84]);
  assign t[262] = (x[86] & x[87]);
  assign t[263] = (x[89] & x[90]);
  assign t[264] = (x[94] & x[95]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[212]);
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[214]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = t[50] ^ t[51];
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] ^ t[57];
  assign t[36] = t[58] ^ t[59];
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[38] = ~(t[62] ^ t[63]);
  assign t[39] = t[64] ^ t[65];
  assign t[3] = t[7] ? t[8] : t[211];
  assign t[40] = t[66] ^ t[67];
  assign t[41] = t[68] ^ t[54];
  assign t[42] = ~(t[37] ^ t[69]);
  assign t[43] = t[10] ^ t[70];
  assign t[44] = ~(t[61] ^ t[40]);
  assign t[45] = ~(t[71] & t[72]);
  assign t[46] = t[215] | t[73];
  assign t[47] = ~(t[74]);
  assign t[48] = ~(t[216]);
  assign t[49] = ~(t[75] & t[217]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[76] ^ t[56];
  assign t[51] = t[77] & t[78];
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] & t[82];
  assign t[54] = t[83] ^ t[84];
  assign t[55] = t[85] ^ t[86];
  assign t[56] = t[87] ? t[88] : t[218];
  assign t[57] = t[89] ^ t[90];
  assign t[58] = t[7] ? t[91] : t[219];
  assign t[59] = t[92] ^ t[93];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = ~(t[94] ^ t[95]);
  assign t[61] = t[96] ^ t[97];
  assign t[62] = t[98] ^ t[99];
  assign t[63] = ~(t[69] ^ t[40]);
  assign t[64] = t[100] ^ t[66];
  assign t[65] = t[101] ^ t[102];
  assign t[66] = t[103];
  assign t[67] = t[101] ^ t[86];
  assign t[68] = t[104] ^ t[105];
  assign t[69] = t[106] ^ t[107];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[108] ^ t[93];
  assign t[71] = ~(t[73] & t[109]);
  assign t[72] = ~(t[220] ^ t[110]);
  assign t[73] = ~(t[111] & t[112]);
  assign t[74] = ~(t[46]);
  assign t[75] = ~(t[221]);
  assign t[76] = t[87] ? t[113] : t[222];
  assign t[77] = ~(t[114]);
  assign t[78] = t[87] ? t[115] : t[223];
  assign t[79] = t[7] ? t[116] : t[224];
  assign t[7] = ~(t[14]);
  assign t[80] = t[214] ^ t[117];
  assign t[81] = ~(t[52] ^ t[118]);
  assign t[82] = t[96] ^ t[119];
  assign t[83] = t[120] ^ t[58];
  assign t[84] = t[92] ^ t[121];
  assign t[85] = t[122] ^ t[100];
  assign t[86] = t[123] & t[124];
  assign t[87] = ~(t[14]);
  assign t[88] = t[218] ^ t[125];
  assign t[89] = t[126] ^ t[51];
  assign t[8] = t[211] ^ t[15];
  assign t[90] = t[127] & t[128];
  assign t[91] = t[219] ^ t[129];
  assign t[92] = t[130] ^ t[131];
  assign t[93] = t[132] & t[133];
  assign t[94] = t[39] ^ t[36];
  assign t[95] = t[134] ^ t[90];
  assign t[96] = t[80] ^ t[106];
  assign t[97] = t[118] ^ t[135];
  assign t[98] = t[136] ^ t[137];
  assign t[99] = t[138] ^ t[131];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind72(x, y);
 input [116:0] x;
 output y;

 wire [273:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[141] ^ t[142];
  assign t[101] = t[143] ^ t[144];
  assign t[102] = t[129] ^ t[59];
  assign t[103] = t[41] ^ t[85];
  assign t[104] = t[145] ^ t[146];
  assign t[105] = t[7] ? t[147] : t[232];
  assign t[106] = ~(t[69] ^ t[97]);
  assign t[107] = t[64] ^ t[148];
  assign t[108] = t[7] ? t[149] : t[233];
  assign t[109] = t[150] ^ t[63];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[151] & t[152];
  assign t[111] = ~(t[153] & t[154]);
  assign t[112] = t[155] ^ t[234];
  assign t[113] = ~(t[228]);
  assign t[114] = t[156] & t[155];
  assign t[115] = t[7] ? t[157] : t[235];
  assign t[116] = ~(t[82]);
  assign t[117] = t[229] ^ t[158];
  assign t[118] = ~t[159];
  assign t[119] = t[160] & t[161];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[7] ? t[162] : t[236];
  assign t[121] = ~(t[87] ^ t[163]);
  assign t[122] = t[78] ^ t[164];
  assign t[123] = t[21] ^ t[165];
  assign t[124] = ~(t[99] ^ t[102]);
  assign t[125] = t[92] ^ t[118];
  assign t[126] = t[27] ? x[56] : x[55];
  assign t[127] = ~(t[164]);
  assign t[128] = ~(t[115]);
  assign t[129] = t[115] ^ t[82];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[166] ^ t[145];
  assign t[131] = t[167] ^ t[168];
  assign t[132] = t[7] ? t[169] : t[237];
  assign t[133] = t[7] ? t[170] : t[238];
  assign t[134] = t[230] ^ t[171];
  assign t[135] = t[231] ^ t[172];
  assign t[136] = t[173] & t[174];
  assign t[137] = t[175] & t[148];
  assign t[138] = ~(t[136] ^ t[176]);
  assign t[139] = t[177] ^ t[178];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[96] ^ t[179];
  assign t[141] = t[180] ^ t[166];
  assign t[142] = t[181] & t[182];
  assign t[143] = t[180] ^ t[145];
  assign t[144] = t[183] & t[184];
  assign t[145] = t[185] ? t[186] : t[239];
  assign t[146] = t[167] ^ t[142];
  assign t[147] = t[232] ^ t[187];
  assign t[148] = t[7] ? t[188] : t[240];
  assign t[149] = t[233] ^ t[189];
  assign t[14] = ~(t[26]);
  assign t[150] = t[190] & t[191];
  assign t[151] = ~(t[125] ^ t[109]);
  assign t[152] = t[80] ^ t[94];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[192] | t[113]);
  assign t[155] = ~(t[241]);
  assign t[156] = ~(t[234]);
  assign t[157] = t[235] ^ t[193];
  assign t[158] = t[7] ? t[194] : t[242];
  assign t[159] = t[7] ? t[195] : t[243];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = ~(t[150] ^ t[196]);
  assign t[161] = t[62] ^ t[197];
  assign t[162] = t[236] ^ t[198];
  assign t[163] = t[53] ^ t[115];
  assign t[164] = t[117] ^ t[82];
  assign t[165] = t[177] ^ t[137];
  assign t[166] = t[185] ? t[199] : t[244];
  assign t[167] = t[200] ^ t[144];
  assign t[168] = t[201] & t[202];
  assign t[169] = t[237] ^ t[203];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[238] ^ t[204];
  assign t[171] = t[205] ? x[82] : x[81];
  assign t[172] = t[76] ? x[84] : x[83];
  assign t[173] = ~(t[178]);
  assign t[174] = ~(t[105]);
  assign t[175] = ~(t[95]);
  assign t[176] = t[64] ^ t[105];
  assign t[177] = t[105] ^ t[96];
  assign t[178] = t[148] ^ t[95];
  assign t[179] = t[97] ^ t[70];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[185] ? t[206] : t[245];
  assign t[181] = ~(t[141] ^ t[167]);
  assign t[182] = t[130] ^ t[184];
  assign t[183] = ~(t[166]);
  assign t[184] = t[185] ? t[207] : t[246];
  assign t[185] = ~(t[14]);
  assign t[186] = t[239] ^ t[208];
  assign t[187] = t[205] ? x[92] : x[91];
  assign t[188] = t[240] ^ t[209];
  assign t[189] = t[76] ? x[94] : x[93];
  assign t[18] = ~(t[32] ^ t[33]);
  assign t[190] = ~(t[197]);
  assign t[191] = ~(t[92]);
  assign t[192] = ~(t[225]);
  assign t[193] = t[27] ? x[96] : x[95];
  assign t[194] = t[242] ^ t[210];
  assign t[195] = t[243] ^ t[211];
  assign t[196] = t[80] ^ t[92];
  assign t[197] = t[94] ^ t[118];
  assign t[198] = t[27] ? x[98] : x[97];
  assign t[199] = t[244] ^ t[212];
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[213] & t[214];
  assign t[201] = ~(t[200] ^ t[215]);
  assign t[202] = t[143] ^ t[216];
  assign t[203] = t[76] ? x[100] : x[99];
  assign t[204] = t[76] ? x[102] : x[101];
  assign t[205] = ~(t[48]);
  assign t[206] = t[245] ^ t[217];
  assign t[207] = t[246] ^ t[218];
  assign t[208] = t[219] ? x[104] : x[103];
  assign t[209] = t[205] ? x[106] : x[105];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[27] ? x[108] : x[107];
  assign t[211] = t[27] ? x[110] : x[109];
  assign t[212] = t[219] ? x[112] : x[111];
  assign t[213] = ~(t[216]);
  assign t[214] = ~(t[180]);
  assign t[215] = t[130] ^ t[180];
  assign t[216] = t[184] ^ t[166];
  assign t[217] = t[219] ? x[114] : x[113];
  assign t[218] = t[219] ? x[116] : x[115];
  assign t[219] = ~(t[48]);
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[4];
  assign t[221] = t[248] ^ x[9];
  assign t[222] = t[249] ^ x[12];
  assign t[223] = t[250] ^ x[15];
  assign t[224] = t[251] ^ x[18];
  assign t[225] = t[252] ^ x[21];
  assign t[226] = t[253] ^ x[24];
  assign t[227] = t[254] ^ x[27];
  assign t[228] = t[255] ^ x[30];
  assign t[229] = t[256] ^ x[33];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[36];
  assign t[231] = t[258] ^ x[39];
  assign t[232] = t[259] ^ x[42];
  assign t[233] = t[260] ^ x[45];
  assign t[234] = t[261] ^ x[48];
  assign t[235] = t[262] ^ x[51];
  assign t[236] = t[263] ^ x[54];
  assign t[237] = t[264] ^ x[59];
  assign t[238] = t[265] ^ x[62];
  assign t[239] = t[266] ^ x[65];
  assign t[23] = ~(t[42] ^ t[20]);
  assign t[240] = t[267] ^ x[68];
  assign t[241] = t[268] ^ x[71];
  assign t[242] = t[269] ^ x[74];
  assign t[243] = t[270] ^ x[77];
  assign t[244] = t[271] ^ x[80];
  assign t[245] = t[272] ^ x[87];
  assign t[246] = t[273] ^ x[90];
  assign t[247] = (x[2] & x[3]);
  assign t[248] = (x[7] & x[8]);
  assign t[249] = (x[10] & x[11]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (x[13] & x[14]);
  assign t[251] = (x[16] & x[17]);
  assign t[252] = (x[19] & x[20]);
  assign t[253] = (x[22] & x[23]);
  assign t[254] = (x[25] & x[26]);
  assign t[255] = (x[28] & x[29]);
  assign t[256] = (x[31] & x[32]);
  assign t[257] = (x[34] & x[35]);
  assign t[258] = (x[37] & x[38]);
  assign t[259] = (x[40] & x[41]);
  assign t[25] = ~(t[34] ^ t[45]);
  assign t[260] = (x[43] & x[44]);
  assign t[261] = (x[46] & x[47]);
  assign t[262] = (x[49] & x[50]);
  assign t[263] = (x[52] & x[53]);
  assign t[264] = (x[57] & x[58]);
  assign t[265] = (x[60] & x[61]);
  assign t[266] = (x[63] & x[64]);
  assign t[267] = (x[66] & x[67]);
  assign t[268] = (x[69] & x[70]);
  assign t[269] = (x[72] & x[73]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[270] = (x[75] & x[76]);
  assign t[271] = (x[78] & x[79]);
  assign t[272] = (x[85] & x[86]);
  assign t[273] = (x[88] & x[89]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[221]);
  assign t[29] = ~(t[222]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[223]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[51] ^ t[13];
  assign t[33] = ~(t[52] ^ t[42]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] ^ t[56]);
  assign t[36] = t[224] ^ t[57];
  assign t[37] = t[58] ^ t[59];
  assign t[38] = t[60] ^ t[61];
  assign t[39] = ~(t[40] ^ t[45]);
  assign t[3] = t[7] ? t[8] : t[220];
  assign t[40] = t[62] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = ~(t[66] ^ t[34]);
  assign t[43] = ~(t[67] ^ t[68]);
  assign t[44] = t[69] ^ t[70];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = ~(t[73] & t[74]);
  assign t[47] = t[225] | t[75];
  assign t[48] = ~(t[76]);
  assign t[49] = ~(t[224]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[77] & t[226]);
  assign t[51] = t[78] ^ t[79];
  assign t[52] = t[80] ^ t[81];
  assign t[53] = t[82] ^ t[36];
  assign t[54] = t[58] ^ t[83];
  assign t[55] = t[84] ^ t[43];
  assign t[56] = ~(t[20] ^ t[85]);
  assign t[57] = t[7] ? t[86] : t[227];
  assign t[58] = t[87] ^ t[79];
  assign t[59] = t[88] & t[89];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[20] ^ t[51];
  assign t[61] = ~(t[90] ^ t[91]);
  assign t[62] = t[92] ^ t[71];
  assign t[63] = t[93] & t[94];
  assign t[64] = t[95] ^ t[96];
  assign t[65] = t[97] ^ t[98];
  assign t[66] = ~(t[99] ^ t[100]);
  assign t[67] = t[101] ^ t[102];
  assign t[68] = ~(t[103] ^ t[104]);
  assign t[69] = t[105] ^ t[95];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[106] & t[107];
  assign t[71] = t[108];
  assign t[72] = t[109] ^ t[110];
  assign t[73] = ~(t[75] & t[111]);
  assign t[74] = ~(t[228] ^ t[112]);
  assign t[75] = ~(t[113] & t[114]);
  assign t[76] = ~(t[47]);
  assign t[77] = ~(t[229]);
  assign t[78] = t[115] ^ t[36];
  assign t[79] = t[116] & t[117];
  assign t[7] = ~(t[14]);
  assign t[80] = t[118] ^ t[71];
  assign t[81] = t[109] ^ t[119];
  assign t[82] = t[223] ^ t[120];
  assign t[83] = t[121] & t[122];
  assign t[84] = ~(t[123] ^ t[124]);
  assign t[85] = t[125] ^ t[110];
  assign t[86] = t[227] ^ t[126];
  assign t[87] = t[127] & t[128];
  assign t[88] = ~(t[129] ^ t[58]);
  assign t[89] = t[53] ^ t[117];
  assign t[8] = t[220] ^ t[15];
  assign t[90] = ~(t[44] ^ t[104]);
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[132];
  assign t[93] = ~(t[118]);
  assign t[94] = t[133];
  assign t[95] = t[7] ? t[134] : t[230];
  assign t[96] = t[7] ? t[135] : t[231];
  assign t[97] = t[136] ^ t[137];
  assign t[98] = t[138] & t[139];
  assign t[99] = t[52] ^ t[140];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind73(x, y);
 input [116:0] x;
 output y;

 wire [264:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[220] ^ t[142];
  assign t[101] = t[221] ^ t[143];
  assign t[102] = t[222] ^ t[144];
  assign t[103] = t[223] ^ t[145];
  assign t[104] = ~(t[116] ^ t[56]);
  assign t[105] = t[34] ^ t[126];
  assign t[106] = t[224] ^ t[146];
  assign t[107] = t[147] & t[148];
  assign t[108] = t[149] & t[150];
  assign t[109] = ~(t[92] ^ t[71]);
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = t[151] ^ t[150];
  assign t[111] = ~(t[152] & t[153]);
  assign t[112] = t[154] ^ t[229];
  assign t[113] = ~(t[225]);
  assign t[114] = t[155] & t[154];
  assign t[115] = t[156] ^ t[61];
  assign t[116] = t[157] ^ t[55];
  assign t[117] = t[121] ^ t[158];
  assign t[118] = t[62] ^ t[159];
  assign t[119] = t[227] ^ t[160];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[161] ^ t[41];
  assign t[121] = t[82] ^ t[65];
  assign t[122] = t[228] ^ t[162];
  assign t[123] = ~(t[129]);
  assign t[124] = ~(t[157]);
  assign t[125] = ~(t[55]);
  assign t[126] = t[226] ^ t[163];
  assign t[127] = t[34] ^ t[157];
  assign t[128] = t[157] ^ t[42];
  assign t[129] = t[126] ^ t[55];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = ~(t[164] ^ t[165]);
  assign t[131] = t[166] ^ t[167];
  assign t[132] = t[168];
  assign t[133] = ~t[169];
  assign t[134] = t[170] ? x[62] : x[61];
  assign t[135] = t[170] ? x[64] : x[63];
  assign t[136] = ~(t[141]);
  assign t[137] = ~(t[156]);
  assign t[138] = ~(t[60]);
  assign t[139] = t[93] ? t[171] : t[230];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[38] ^ t[156];
  assign t[141] = t[139] ^ t[60];
  assign t[142] = t[172] ? x[69] : x[68];
  assign t[143] = t[76] ? x[71] : x[70];
  assign t[144] = t[172] ? x[73] : x[72];
  assign t[145] = t[27] ? x[75] : x[74];
  assign t[146] = t[76] ? x[77] : x[76];
  assign t[147] = ~(t[173]);
  assign t[148] = ~(t[132]);
  assign t[149] = ~(t[133]);
  assign t[14] = ~(t[26]);
  assign t[150] = t[174];
  assign t[151] = t[133] ^ t[44];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[175] | t[113]);
  assign t[154] = ~(t[231]);
  assign t[155] = ~(t[229]);
  assign t[156] = t[93] ? t[176] : t[232];
  assign t[157] = t[7] ? t[177] : t[233];
  assign t[158] = t[120] ^ t[178];
  assign t[159] = t[179] & t[180];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[172] ? x[88] : x[87];
  assign t[161] = t[181] & t[182];
  assign t[162] = t[27] ? x[90] : x[89];
  assign t[163] = t[7] ? t[183] : t[234];
  assign t[164] = t[184] ^ t[185];
  assign t[165] = ~(t[186] ^ t[25]);
  assign t[166] = t[151] ^ t[187];
  assign t[167] = t[65] ^ t[188];
  assign t[168] = t[7] ? t[189] : t[235];
  assign t[169] = t[7] ? t[190] : t[236];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = ~(t[48]);
  assign t[171] = t[230] ^ t[191];
  assign t[172] = ~(t[48]);
  assign t[173] = t[150] ^ t[133];
  assign t[174] = t[7] ? t[192] : t[237];
  assign t[175] = ~(t[216]);
  assign t[176] = t[232] ^ t[193];
  assign t[177] = t[233] ^ t[194];
  assign t[178] = t[195] & t[196];
  assign t[179] = ~(t[197] ^ t[62]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[38] ^ t[139];
  assign t[181] = ~(t[198]);
  assign t[182] = ~(t[64]);
  assign t[183] = t[234] ^ t[199];
  assign t[184] = t[24] ^ t[200];
  assign t[185] = ~(t[201] ^ t[22]);
  assign t[186] = t[202] ^ t[108];
  assign t[187] = t[71] ^ t[203];
  assign t[188] = t[120] ^ t[54];
  assign t[189] = t[235] ^ t[204];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[236] ^ t[205];
  assign t[191] = t[170] ? x[104] : x[103];
  assign t[192] = t[237] ^ t[206];
  assign t[193] = t[170] ? x[106] : x[105];
  assign t[194] = t[27] ? x[108] : x[107];
  assign t[195] = ~(t[161] ^ t[207]);
  assign t[196] = t[40] ^ t[198];
  assign t[197] = t[156] ^ t[60];
  assign t[198] = t[67] ^ t[82];
  assign t[199] = t[27] ? x[110] : x[109];
  assign t[19] = ~(t[20] ^ t[25]);
  assign t[1] = ~(t[4]);
  assign t[200] = t[128] ^ t[87];
  assign t[201] = ~(t[33] ^ t[81]);
  assign t[202] = t[132] ^ t[44];
  assign t[203] = t[208] & t[209];
  assign t[204] = t[76] ? x[112] : x[111];
  assign t[205] = t[27] ? x[114] : x[113];
  assign t[206] = t[76] ? x[116] : x[115];
  assign t[207] = t[121] ^ t[64];
  assign t[208] = ~(t[107] ^ t[210]);
  assign t[209] = t[202] ^ t[173];
  assign t[20] = t[34] ^ t[35];
  assign t[210] = t[151] ^ t[132];
  assign t[211] = t[238] ^ x[4];
  assign t[212] = t[239] ^ x[9];
  assign t[213] = t[240] ^ x[12];
  assign t[214] = t[241] ^ x[15];
  assign t[215] = t[242] ^ x[18];
  assign t[216] = t[243] ^ x[21];
  assign t[217] = t[244] ^ x[24];
  assign t[218] = t[245] ^ x[27];
  assign t[219] = t[246] ^ x[30];
  assign t[21] = ~(t[36] ^ t[37]);
  assign t[220] = t[247] ^ x[33];
  assign t[221] = t[248] ^ x[36];
  assign t[222] = t[249] ^ x[39];
  assign t[223] = t[250] ^ x[42];
  assign t[224] = t[251] ^ x[45];
  assign t[225] = t[252] ^ x[48];
  assign t[226] = t[253] ^ x[51];
  assign t[227] = t[254] ^ x[54];
  assign t[228] = t[255] ^ x[57];
  assign t[229] = t[256] ^ x[60];
  assign t[22] = t[38] ^ t[39];
  assign t[230] = t[257] ^ x[67];
  assign t[231] = t[258] ^ x[80];
  assign t[232] = t[259] ^ x[83];
  assign t[233] = t[260] ^ x[86];
  assign t[234] = t[261] ^ x[93];
  assign t[235] = t[262] ^ x[96];
  assign t[236] = t[263] ^ x[99];
  assign t[237] = t[264] ^ x[102];
  assign t[238] = (x[2] & x[3]);
  assign t[239] = (x[7] & x[8]);
  assign t[23] = t[40] ^ t[41];
  assign t[240] = (x[10] & x[11]);
  assign t[241] = (x[13] & x[14]);
  assign t[242] = (x[16] & x[17]);
  assign t[243] = (x[19] & x[20]);
  assign t[244] = (x[22] & x[23]);
  assign t[245] = (x[25] & x[26]);
  assign t[246] = (x[28] & x[29]);
  assign t[247] = (x[31] & x[32]);
  assign t[248] = (x[34] & x[35]);
  assign t[249] = (x[37] & x[38]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (x[40] & x[41]);
  assign t[251] = (x[43] & x[44]);
  assign t[252] = (x[46] & x[47]);
  assign t[253] = (x[49] & x[50]);
  assign t[254] = (x[52] & x[53]);
  assign t[255] = (x[55] & x[56]);
  assign t[256] = (x[58] & x[59]);
  assign t[257] = (x[65] & x[66]);
  assign t[258] = (x[78] & x[79]);
  assign t[259] = (x[81] & x[82]);
  assign t[25] = t[44] ^ t[45];
  assign t[260] = (x[84] & x[85]);
  assign t[261] = (x[91] & x[92]);
  assign t[262] = (x[94] & x[95]);
  assign t[263] = (x[97] & x[98]);
  assign t[264] = (x[100] & x[101]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[212]);
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[214]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = ~(t[51] ^ t[52]);
  assign t[33] = t[53] ^ t[54];
  assign t[34] = t[55] ^ t[42];
  assign t[35] = t[56] ^ t[57];
  assign t[36] = t[58] ^ t[32];
  assign t[37] = ~(t[24] ^ t[59]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[62] ^ t[63];
  assign t[3] = t[7] ? t[8] : t[211];
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[66] & t[67];
  assign t[42] = t[215] ^ t[68];
  assign t[43] = t[56] ^ t[69];
  assign t[44] = t[70];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = ~(t[73] & t[74]);
  assign t[47] = t[216] | t[75];
  assign t[48] = ~(t[76]);
  assign t[49] = ~(t[215]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[77] & t[217]);
  assign t[51] = t[78] ^ t[79];
  assign t[52] = ~(t[80] ^ t[81]);
  assign t[53] = t[64] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[214] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] & t[89];
  assign t[58] = ~(t[90] ^ t[91]);
  assign t[59] = t[92] ^ t[72];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[93] ? t[94] : t[218];
  assign t[61] = t[93] ? t[95] : t[219];
  assign t[62] = t[96] ^ t[97];
  assign t[63] = t[98] & t[99];
  assign t[64] = t[7] ? t[100] : t[220];
  assign t[65] = t[7] ? t[101] : t[221];
  assign t[66] = ~(t[82]);
  assign t[67] = t[7] ? t[102] : t[222];
  assign t[68] = t[7] ? t[103] : t[223];
  assign t[69] = t[104] & t[105];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[7] ? t[106] : t[224];
  assign t[71] = t[107] ^ t[108];
  assign t[72] = t[109] & t[110];
  assign t[73] = ~(t[75] & t[111]);
  assign t[74] = ~(t[225] ^ t[112]);
  assign t[75] = ~(t[113] & t[114]);
  assign t[76] = ~(t[47]);
  assign t[77] = ~(t[226]);
  assign t[78] = t[115] ^ t[97];
  assign t[79] = t[116] ^ t[69];
  assign t[7] = ~(t[14]);
  assign t[80] = t[117] ^ t[59];
  assign t[81] = t[61] ^ t[118];
  assign t[82] = t[7] ? t[119] : t[227];
  assign t[83] = ~(t[53] ^ t[120]);
  assign t[84] = t[121] ^ t[67];
  assign t[85] = t[7] ? t[122] : t[228];
  assign t[86] = t[123] & t[124];
  assign t[87] = t[125] & t[126];
  assign t[88] = ~(t[86] ^ t[127]);
  assign t[89] = t[128] ^ t[129];
  assign t[8] = t[211] ^ t[15];
  assign t[90] = t[130] ^ t[23];
  assign t[91] = ~(t[131] ^ t[79]);
  assign t[92] = t[132] ^ t[133];
  assign t[93] = ~(t[14]);
  assign t[94] = t[218] ^ t[134];
  assign t[95] = t[219] ^ t[135];
  assign t[96] = t[136] & t[137];
  assign t[97] = t[138] & t[139];
  assign t[98] = ~(t[96] ^ t[140]);
  assign t[99] = t[115] ^ t[141];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind74(x, y);
 input [116:0] x;
 output y;

 wire [262:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[216] ^ t[142];
  assign t[101] = t[217] ^ t[143];
  assign t[102] = t[26] ? t[144] : t[225];
  assign t[103] = ~(t[145] & t[146]);
  assign t[104] = t[147] ^ t[226];
  assign t[105] = ~(t[218]);
  assign t[106] = t[148] & t[147];
  assign t[107] = t[86] ^ t[126];
  assign t[108] = t[149] & t[150];
  assign t[109] = t[215] ^ t[151];
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = t[111] ^ t[61];
  assign t[111] = t[152] ^ t[153];
  assign t[112] = t[154] & t[155];
  assign t[113] = t[220] ^ t[156];
  assign t[114] = t[157] ^ t[58];
  assign t[115] = t[126] ^ t[77];
  assign t[116] = t[114] ^ t[158];
  assign t[117] = t[159] ^ t[128];
  assign t[118] = t[160] & t[161];
  assign t[119] = t[62] ^ t[162];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[140] ^ t[97];
  assign t[121] = t[159] ^ t[123];
  assign t[122] = t[163] & t[164];
  assign t[123] = t[7] ? t[165] : t[227];
  assign t[124] = t[129] ^ t[118];
  assign t[125] = t[221] ^ t[166];
  assign t[126] = t[26] ? t[167] : t[228];
  assign t[127] = t[222] ^ t[168];
  assign t[128] = t[7] ? t[169] : t[229];
  assign t[129] = t[170] ^ t[122];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[171] & t[172];
  assign t[131] = ~(t[14]);
  assign t[132] = t[223] ^ t[173];
  assign t[133] = t[131] ? t[174] : t[230];
  assign t[134] = t[211] ^ t[175];
  assign t[135] = t[224] ^ t[176];
  assign t[136] = ~(t[141]);
  assign t[137] = ~(t[41]);
  assign t[138] = ~(t[42]);
  assign t[139] = t[39] ^ t[41];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[41] ^ t[62];
  assign t[141] = t[67] ^ t[42];
  assign t[142] = t[177] ? x[71] : x[70];
  assign t[143] = t[177] ? x[73] : x[72];
  assign t[144] = t[225] ^ t[178];
  assign t[145] = ~(t[148] | t[147]);
  assign t[146] = ~(t[179] | t[105]);
  assign t[147] = ~(t[231]);
  assign t[148] = ~(t[226]);
  assign t[149] = ~(t[107] ^ t[114]);
  assign t[14] = ~(t[26]);
  assign t[150] = t[115] ^ t[88];
  assign t[151] = t[131] ? t[180] : t[232];
  assign t[152] = t[181] & t[182];
  assign t[153] = t[183] & t[134];
  assign t[154] = ~(t[152] ^ t[184]);
  assign t[155] = t[185] ^ t[186];
  assign t[156] = t[71] ? x[81] : x[80];
  assign t[157] = t[187] & t[188];
  assign t[158] = t[189] & t[190];
  assign t[159] = t[7] ? t[191] : t[233];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = ~(t[117] ^ t[129]);
  assign t[161] = t[89] ^ t[164];
  assign t[162] = t[63] ^ t[25];
  assign t[163] = ~(t[128]);
  assign t[164] = t[7] ? t[192] : t[234];
  assign t[165] = t[227] ^ t[193];
  assign t[166] = t[27] ? x[89] : x[88];
  assign t[167] = t[228] ^ t[194];
  assign t[168] = t[71] ? x[91] : x[90];
  assign t[169] = t[229] ^ t[195];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[196] & t[197];
  assign t[171] = ~(t[170] ^ t[198]);
  assign t[172] = t[121] ^ t[199];
  assign t[173] = t[200] ? x[93] : x[92];
  assign t[174] = t[230] ^ t[201];
  assign t[175] = t[131] ? t[202] : t[235];
  assign t[176] = t[177] ? x[98] : x[97];
  assign t[177] = ~(t[47]);
  assign t[178] = t[177] ? x[100] : x[99];
  assign t[179] = ~(t[213]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[232] ^ t[203];
  assign t[181] = ~(t[186]);
  assign t[182] = ~(t[91]);
  assign t[183] = ~(t[92]);
  assign t[184] = t[75] ^ t[91];
  assign t[185] = t[91] ^ t[109];
  assign t[186] = t[134] ^ t[92];
  assign t[187] = ~(t[204]);
  assign t[188] = ~(t[86]);
  assign t[189] = ~(t[157] ^ t[205]);
  assign t[18] = ~(t[23] ^ t[32]);
  assign t[190] = t[57] ^ t[204];
  assign t[191] = t[233] ^ t[206];
  assign t[192] = t[234] ^ t[207];
  assign t[193] = t[177] ? x[102] : x[101];
  assign t[194] = t[27] ? x[104] : x[103];
  assign t[195] = t[177] ? x[106] : x[105];
  assign t[196] = ~(t[199]);
  assign t[197] = ~(t[159]);
  assign t[198] = t[89] ^ t[159];
  assign t[199] = t[164] ^ t[128];
  assign t[19] = ~(t[33] ^ t[34]);
  assign t[1] = ~(t[4]);
  assign t[200] = ~(t[47]);
  assign t[201] = t[200] ? x[108] : x[107];
  assign t[202] = t[235] ^ t[208];
  assign t[203] = t[200] ? x[110] : x[109];
  assign t[204] = t[88] ^ t[126];
  assign t[205] = t[115] ^ t[86];
  assign t[206] = t[177] ? x[112] : x[111];
  assign t[207] = t[177] ? x[114] : x[113];
  assign t[208] = t[200] ? x[116] : x[115];
  assign t[209] = t[236] ^ x[4];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[237] ^ x[9];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[37] ^ t[13]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[60];
  assign t[228] = t[255] ^ x[63];
  assign t[229] = t[256] ^ x[66];
  assign t[22] = ~(t[37] ^ t[38]);
  assign t[230] = t[257] ^ x[69];
  assign t[231] = t[258] ^ x[76];
  assign t[232] = t[259] ^ x[79];
  assign t[233] = t[260] ^ x[84];
  assign t[234] = t[261] ^ x[87];
  assign t[235] = t[262] ^ x[96];
  assign t[236] = (x[2] & x[3]);
  assign t[237] = (x[7] & x[8]);
  assign t[238] = (x[10] & x[11]);
  assign t[239] = (x[13] & x[14]);
  assign t[23] = t[39] ^ t[40];
  assign t[240] = (x[16] & x[17]);
  assign t[241] = (x[19] & x[20]);
  assign t[242] = (x[22] & x[23]);
  assign t[243] = (x[25] & x[26]);
  assign t[244] = (x[28] & x[29]);
  assign t[245] = (x[31] & x[32]);
  assign t[246] = (x[34] & x[35]);
  assign t[247] = (x[37] & x[38]);
  assign t[248] = (x[40] & x[41]);
  assign t[249] = (x[43] & x[44]);
  assign t[24] = t[41] ^ t[42];
  assign t[250] = (x[46] & x[47]);
  assign t[251] = (x[49] & x[50]);
  assign t[252] = (x[52] & x[53]);
  assign t[253] = (x[55] & x[56]);
  assign t[254] = (x[58] & x[59]);
  assign t[255] = (x[61] & x[62]);
  assign t[256] = (x[64] & x[65]);
  assign t[257] = (x[67] & x[68]);
  assign t[258] = (x[74] & x[75]);
  assign t[259] = (x[77] & x[78]);
  assign t[25] = t[43] & t[44];
  assign t[260] = (x[82] & x[83]);
  assign t[261] = (x[85] & x[86]);
  assign t[262] = (x[94] & x[95]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[210]);
  assign t[29] = ~(t[211]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[212]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = ~(t[50] ^ t[51]);
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[34] = t[12] ^ t[54];
  assign t[35] = ~(t[55] ^ t[56]);
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ t[52];
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[42] ^ t[62];
  assign t[3] = t[7] ? t[8] : t[209];
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65];
  assign t[42] = ~t[66];
  assign t[43] = ~(t[24] ^ t[63]);
  assign t[44] = t[39] ^ t[67];
  assign t[45] = ~(t[68] & t[69]);
  assign t[46] = t[213] | t[70];
  assign t[47] = ~(t[71]);
  assign t[48] = ~(t[214]);
  assign t[49] = ~(t[72] & t[215]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[73] ^ t[74]);
  assign t[51] = t[75] ^ t[76];
  assign t[52] = t[77] ^ t[78];
  assign t[53] = t[79] ^ t[80];
  assign t[54] = ~(t[81] ^ t[82]);
  assign t[55] = t[83] ^ t[32];
  assign t[56] = ~(t[84] ^ t[85]);
  assign t[57] = t[86] ^ t[77];
  assign t[58] = t[87] & t[88];
  assign t[59] = t[89] ^ t[90];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[91] ^ t[92];
  assign t[61] = t[93] & t[94];
  assign t[62] = ~t[95];
  assign t[63] = t[96] ^ t[97];
  assign t[64] = t[98] & t[99];
  assign t[65] = t[7] ? t[100] : t[216];
  assign t[66] = t[7] ? t[101] : t[217];
  assign t[67] = t[102];
  assign t[68] = ~(t[70] & t[103]);
  assign t[69] = ~(t[218] ^ t[104]);
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[105] & t[106]);
  assign t[71] = ~(t[46]);
  assign t[72] = ~(t[219]);
  assign t[73] = t[107] ^ t[108];
  assign t[74] = t[109] ^ t[110];
  assign t[75] = t[92] ^ t[109];
  assign t[76] = t[111] ^ t[112];
  assign t[77] = t[26] ? t[113] : t[220];
  assign t[78] = t[114] ^ t[108];
  assign t[79] = t[115] ^ t[116];
  assign t[7] = ~(t[14]);
  assign t[80] = t[117] ^ t[118];
  assign t[81] = t[51] ^ t[36];
  assign t[82] = ~(t[119] ^ t[85]);
  assign t[83] = t[119] ^ t[120];
  assign t[84] = t[121] ^ t[122];
  assign t[85] = t[123] ^ t[124];
  assign t[86] = t[26] ? t[125] : t[221];
  assign t[87] = ~(t[126]);
  assign t[88] = t[26] ? t[127] : t[222];
  assign t[89] = t[128] ^ t[123];
  assign t[8] = t[209] ^ t[15];
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[131] ? t[132] : t[223];
  assign t[92] = t[210] ^ t[133];
  assign t[93] = ~(t[60] ^ t[111]);
  assign t[94] = t[75] ^ t[134];
  assign t[95] = t[7] ? t[135] : t[224];
  assign t[96] = t[136] & t[137];
  assign t[97] = t[138] & t[67];
  assign t[98] = ~(t[96] ^ t[139]);
  assign t[99] = t[140] ^ t[141];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind75(x, y);
 input [116:0] x;
 output y;

 wire [264:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[140] ^ t[104];
  assign t[101] = t[141] & t[142];
  assign t[102] = t[219] ^ t[143];
  assign t[103] = t[122] ^ t[66];
  assign t[104] = t[144] & t[145];
  assign t[105] = ~t[146];
  assign t[106] = t[118] ^ t[53];
  assign t[107] = t[147] ^ t[120];
  assign t[108] = ~(t[148] & t[149]);
  assign t[109] = t[150] ^ t[225];
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = ~(t[220]);
  assign t[111] = t[151] & t[150];
  assign t[112] = ~(t[14]);
  assign t[113] = t[222] ^ t[152];
  assign t[114] = t[212] ^ t[153];
  assign t[115] = t[112] ? t[154] : t[226];
  assign t[116] = t[7] ? t[155] : t[227];
  assign t[117] = t[7] ? t[156] : t[228];
  assign t[118] = t[157] ^ t[158];
  assign t[119] = t[159];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[26] ? t[160] : t[229];
  assign t[121] = t[161] & t[162];
  assign t[122] = t[7] ? t[163] : t[230];
  assign t[123] = ~(t[85] ^ t[100]);
  assign t[124] = t[64] ^ t[145];
  assign t[125] = t[223] ^ t[164];
  assign t[126] = t[165] & t[166];
  assign t[127] = ~(t[134] ^ t[88]);
  assign t[128] = t[136] ^ t[78];
  assign t[129] = t[74] ? x[65] : x[64];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[167] & t[168];
  assign t[131] = t[169] & t[170];
  assign t[132] = ~(t[107] ^ t[91]);
  assign t[133] = t[83] ^ t[170];
  assign t[134] = t[76] ^ t[114];
  assign t[135] = t[171] & t[172];
  assign t[136] = t[114] ^ t[56];
  assign t[137] = t[88] ^ t[173];
  assign t[138] = t[147] ^ t[58];
  assign t[139] = t[224] ^ t[174];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[175] & t[176];
  assign t[141] = ~(t[140] ^ t[177]);
  assign t[142] = t[103] ^ t[178];
  assign t[143] = t[179] ? x[67] : x[66];
  assign t[144] = ~(t[99]);
  assign t[145] = t[7] ? t[180] : t[231];
  assign t[146] = t[7] ? t[181] : t[232];
  assign t[147] = t[26] ? t[182] : t[233];
  assign t[148] = ~(t[151] | t[150]);
  assign t[149] = ~(t[183] | t[110]);
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[234]);
  assign t[151] = ~(t[225]);
  assign t[152] = t[184] ? x[81] : x[80];
  assign t[153] = t[112] ? t[185] : t[235];
  assign t[154] = t[226] ^ t[186];
  assign t[155] = t[227] ^ t[187];
  assign t[156] = t[228] ^ t[188];
  assign t[157] = t[189] & t[190];
  assign t[158] = t[191] & t[119];
  assign t[159] = t[26] ? t[192] : t[236];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[229] ^ t[193];
  assign t[161] = ~(t[130] ^ t[194]);
  assign t[162] = t[138] ^ t[195];
  assign t[163] = t[230] ^ t[196];
  assign t[164] = t[184] ? x[89] : x[88];
  assign t[165] = ~(t[197]);
  assign t[166] = ~(t[76]);
  assign t[167] = ~(t[195]);
  assign t[168] = ~(t[147]);
  assign t[169] = ~(t[120]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[26] ? t[198] : t[237];
  assign t[171] = ~(t[157] ^ t[199]);
  assign t[172] = t[200] ^ t[201];
  assign t[173] = t[202] & t[203];
  assign t[174] = t[179] ? x[94] : x[93];
  assign t[175] = ~(t[178]);
  assign t[176] = ~(t[122]);
  assign t[177] = t[64] ^ t[122];
  assign t[178] = t[145] ^ t[99];
  assign t[179] = ~(t[47]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[231] ^ t[204];
  assign t[181] = t[232] ^ t[205];
  assign t[182] = t[233] ^ t[206];
  assign t[183] = ~(t[215]);
  assign t[184] = ~(t[47]);
  assign t[185] = t[235] ^ t[207];
  assign t[186] = t[184] ? x[96] : x[95];
  assign t[187] = t[179] ? x[98] : x[97];
  assign t[188] = t[179] ? x[100] : x[99];
  assign t[189] = ~(t[201]);
  assign t[18] = t[32] ^ t[33];
  assign t[190] = ~(t[79]);
  assign t[191] = ~(t[80]);
  assign t[192] = t[236] ^ t[208];
  assign t[193] = t[27] ? x[102] : x[101];
  assign t[194] = t[83] ^ t[147];
  assign t[195] = t[170] ^ t[120];
  assign t[196] = t[179] ? x[104] : x[103];
  assign t[197] = t[78] ^ t[114];
  assign t[198] = t[237] ^ t[209];
  assign t[199] = t[95] ^ t[79];
  assign t[19] = ~(t[34] ^ t[35]);
  assign t[1] = ~(t[4]);
  assign t[200] = t[79] ^ t[105];
  assign t[201] = t[119] ^ t[80];
  assign t[202] = ~(t[126] ^ t[210]);
  assign t[203] = t[50] ^ t[197];
  assign t[204] = t[179] ? x[106] : x[105];
  assign t[205] = t[179] ? x[108] : x[107];
  assign t[206] = t[27] ? x[110] : x[109];
  assign t[207] = t[184] ? x[112] : x[111];
  assign t[208] = t[179] ? x[114] : x[113];
  assign t[209] = t[74] ? x[116] : x[115];
  assign t[20] = ~(t[36] ^ t[34]);
  assign t[210] = t[136] ^ t[76];
  assign t[211] = t[238] ^ x[4];
  assign t[212] = t[239] ^ x[9];
  assign t[213] = t[240] ^ x[12];
  assign t[214] = t[241] ^ x[15];
  assign t[215] = t[242] ^ x[18];
  assign t[216] = t[243] ^ x[21];
  assign t[217] = t[244] ^ x[24];
  assign t[218] = t[245] ^ x[27];
  assign t[219] = t[246] ^ x[30];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[33];
  assign t[221] = t[248] ^ x[36];
  assign t[222] = t[249] ^ x[39];
  assign t[223] = t[250] ^ x[42];
  assign t[224] = t[251] ^ x[45];
  assign t[225] = t[252] ^ x[48];
  assign t[226] = t[253] ^ x[51];
  assign t[227] = t[254] ^ x[54];
  assign t[228] = t[255] ^ x[57];
  assign t[229] = t[256] ^ x[60];
  assign t[22] = t[21] ^ t[33];
  assign t[230] = t[257] ^ x[63];
  assign t[231] = t[258] ^ x[70];
  assign t[232] = t[259] ^ x[73];
  assign t[233] = t[260] ^ x[76];
  assign t[234] = t[261] ^ x[79];
  assign t[235] = t[262] ^ x[84];
  assign t[236] = t[263] ^ x[87];
  assign t[237] = t[264] ^ x[92];
  assign t[238] = (x[2] & x[3]);
  assign t[239] = (x[7] & x[8]);
  assign t[23] = ~(t[39] ^ t[40]);
  assign t[240] = (x[10] & x[11]);
  assign t[241] = (x[13] & x[14]);
  assign t[242] = (x[16] & x[17]);
  assign t[243] = (x[19] & x[20]);
  assign t[244] = (x[22] & x[23]);
  assign t[245] = (x[25] & x[26]);
  assign t[246] = (x[28] & x[29]);
  assign t[247] = (x[31] & x[32]);
  assign t[248] = (x[34] & x[35]);
  assign t[249] = (x[37] & x[38]);
  assign t[24] = ~(t[41] ^ t[42]);
  assign t[250] = (x[40] & x[41]);
  assign t[251] = (x[43] & x[44]);
  assign t[252] = (x[46] & x[47]);
  assign t[253] = (x[49] & x[50]);
  assign t[254] = (x[52] & x[53]);
  assign t[255] = (x[55] & x[56]);
  assign t[256] = (x[58] & x[59]);
  assign t[257] = (x[61] & x[62]);
  assign t[258] = (x[68] & x[69]);
  assign t[259] = (x[71] & x[72]);
  assign t[25] = ~(t[43] ^ t[44]);
  assign t[260] = (x[74] & x[75]);
  assign t[261] = (x[77] & x[78]);
  assign t[262] = (x[82] & x[83]);
  assign t[263] = (x[85] & x[86]);
  assign t[264] = (x[90] & x[91]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[212]);
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[214]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = t[50] ^ t[51];
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] ^ t[57];
  assign t[36] = t[58] ^ t[59];
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[38] = ~(t[62] ^ t[63]);
  assign t[39] = t[64] ^ t[65];
  assign t[3] = t[7] ? t[8] : t[211];
  assign t[40] = t[66] ^ t[67];
  assign t[41] = t[68] ^ t[54];
  assign t[42] = ~(t[37] ^ t[69]);
  assign t[43] = t[10] ^ t[70];
  assign t[44] = ~(t[61] ^ t[40]);
  assign t[45] = ~(t[71] & t[72]);
  assign t[46] = t[215] | t[73];
  assign t[47] = ~(t[74]);
  assign t[48] = ~(t[216]);
  assign t[49] = ~(t[75] & t[217]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[76] ^ t[56];
  assign t[51] = t[77] & t[78];
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] & t[82];
  assign t[54] = t[83] ^ t[84];
  assign t[55] = t[85] ^ t[86];
  assign t[56] = t[217] ^ t[87];
  assign t[57] = t[88] ^ t[89];
  assign t[58] = t[26] ? t[90] : t[218];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = ~(t[93] ^ t[94]);
  assign t[61] = t[95] ^ t[96];
  assign t[62] = t[97] ^ t[98];
  assign t[63] = ~(t[69] ^ t[40]);
  assign t[64] = t[99] ^ t[66];
  assign t[65] = t[100] ^ t[101];
  assign t[66] = t[7] ? t[102] : t[219];
  assign t[67] = t[100] ^ t[86];
  assign t[68] = t[103] ^ t[104];
  assign t[69] = t[105] ^ t[106];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[107] ^ t[92];
  assign t[71] = ~(t[73] & t[108]);
  assign t[72] = ~(t[220] ^ t[109]);
  assign t[73] = ~(t[110] & t[111]);
  assign t[74] = ~(t[46]);
  assign t[75] = ~(t[221]);
  assign t[76] = t[112] ? t[113] : t[222];
  assign t[77] = ~(t[114]);
  assign t[78] = t[213] ^ t[115];
  assign t[79] = t[116];
  assign t[7] = ~(t[14]);
  assign t[80] = ~t[117];
  assign t[81] = ~(t[52] ^ t[118]);
  assign t[82] = t[95] ^ t[119];
  assign t[83] = t[120] ^ t[58];
  assign t[84] = t[91] ^ t[121];
  assign t[85] = t[122] ^ t[99];
  assign t[86] = t[123] & t[124];
  assign t[87] = t[112] ? t[125] : t[223];
  assign t[88] = t[126] ^ t[51];
  assign t[89] = t[127] & t[128];
  assign t[8] = t[211] ^ t[15];
  assign t[90] = t[218] ^ t[129];
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[132] & t[133];
  assign t[93] = t[39] ^ t[36];
  assign t[94] = t[134] ^ t[89];
  assign t[95] = t[80] ^ t[105];
  assign t[96] = t[118] ^ t[135];
  assign t[97] = t[136] ^ t[137];
  assign t[98] = t[138] ^ t[131];
  assign t[99] = t[7] ? t[139] : t[224];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind76(x, y);
 input [116:0] x;
 output y;

 wire [271:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[127] ^ t[58];
  assign t[101] = t[42] ^ t[83];
  assign t[102] = t[143] ^ t[144];
  assign t[103] = t[30] ? t[145] : t[233];
  assign t[104] = ~(t[68] ^ t[95]);
  assign t[105] = t[63] ^ t[146];
  assign t[106] = t[227] ^ t[147];
  assign t[107] = t[148] ^ t[62];
  assign t[108] = t[149] & t[150];
  assign t[109] = ~(t[151] & t[152]);
  assign t[10] = ~(t[219]);
  assign t[110] = t[153] ^ t[234];
  assign t[111] = ~(t[228]);
  assign t[112] = t[154] & t[153];
  assign t[113] = t[155];
  assign t[114] = ~(t[80]);
  assign t[115] = t[156];
  assign t[116] = t[8] ? t[157] : t[235];
  assign t[117] = t[158] & t[159];
  assign t[118] = t[8] ? t[160] : t[236];
  assign t[119] = ~(t[85] ^ t[161]);
  assign t[11] = ~(t[220]);
  assign t[120] = t[76] ^ t[162];
  assign t[121] = t[25] ^ t[163];
  assign t[122] = ~(t[97] ^ t[100]);
  assign t[123] = t[90] ^ t[116];
  assign t[124] = t[164] ? x[62] : x[61];
  assign t[125] = ~(t[162]);
  assign t[126] = ~(t[113]);
  assign t[127] = t[113] ^ t[80];
  assign t[128] = t[165] ^ t[143];
  assign t[129] = t[166] ^ t[167];
  assign t[12] = ~(t[221]);
  assign t[130] = t[229] ^ t[168];
  assign t[131] = t[230] ^ t[169];
  assign t[132] = t[231] ^ t[170];
  assign t[133] = t[232] ^ t[171];
  assign t[134] = t[172] & t[173];
  assign t[135] = t[174] & t[146];
  assign t[136] = ~(t[134] ^ t[175]);
  assign t[137] = t[176] ^ t[177];
  assign t[138] = t[94] ^ t[178];
  assign t[139] = t[179] ^ t[165];
  assign t[13] = ~(t[20] | t[21]);
  assign t[140] = t[180] & t[181];
  assign t[141] = t[179] ^ t[143];
  assign t[142] = t[182] & t[183];
  assign t[143] = t[223] ^ t[184];
  assign t[144] = t[166] ^ t[140];
  assign t[145] = t[233] ^ t[185];
  assign t[146] = t[30] ? t[186] : t[237];
  assign t[147] = t[164] ? x[67] : x[66];
  assign t[148] = t[187] & t[188];
  assign t[149] = ~(t[123] ^ t[107]);
  assign t[14] = t[22] ^ t[23];
  assign t[150] = t[78] ^ t[92];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[189] | t[111]);
  assign t[153] = ~(t[238]);
  assign t[154] = ~(t[234]);
  assign t[155] = t[8] ? t[190] : t[239];
  assign t[156] = t[30] ? t[191] : t[240];
  assign t[157] = t[235] ^ t[192];
  assign t[158] = ~(t[148] ^ t[193]);
  assign t[159] = t[61] ^ t[194];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = t[236] ^ t[195];
  assign t[161] = t[52] ^ t[113];
  assign t[162] = t[115] ^ t[80];
  assign t[163] = t[176] ^ t[135];
  assign t[164] = ~(t[49]);
  assign t[165] = t[219] ^ t[196];
  assign t[166] = t[197] ^ t[142];
  assign t[167] = t[198] & t[199];
  assign t[168] = t[164] ? x[78] : x[77];
  assign t[169] = t[164] ? x[80] : x[79];
  assign t[16] = ~(t[26] ^ t[27]);
  assign t[170] = t[31] ? x[82] : x[81];
  assign t[171] = t[75] ? x[84] : x[83];
  assign t[172] = ~(t[177]);
  assign t[173] = ~(t[103]);
  assign t[174] = ~(t[93]);
  assign t[175] = t[63] ^ t[103];
  assign t[176] = t[103] ^ t[94];
  assign t[177] = t[146] ^ t[93];
  assign t[178] = t[95] ^ t[69];
  assign t[179] = t[200] ? t[201] : t[241];
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[180] = ~(t[139] ^ t[166]);
  assign t[181] = t[128] ^ t[183];
  assign t[182] = ~(t[165]);
  assign t[183] = t[220] ^ t[202];
  assign t[184] = t[200] ? t[203] : t[242];
  assign t[185] = t[31] ? x[92] : x[91];
  assign t[186] = t[237] ^ t[204];
  assign t[187] = ~(t[194]);
  assign t[188] = ~(t[90]);
  assign t[189] = ~(t[225]);
  assign t[18] = ~(t[30]);
  assign t[190] = t[239] ^ t[205];
  assign t[191] = t[240] ^ t[206];
  assign t[192] = t[164] ? x[94] : x[93];
  assign t[193] = t[78] ^ t[90];
  assign t[194] = t[92] ^ t[116];
  assign t[195] = t[164] ? x[96] : x[95];
  assign t[196] = t[200] ? t[207] : t[243];
  assign t[197] = t[208] & t[209];
  assign t[198] = ~(t[197] ^ t[210]);
  assign t[199] = t[141] ^ t[211];
  assign t[19] = t[31] ? x[15] : x[14];
  assign t[1] = ~(t[4] | t[5]);
  assign t[200] = ~(t[18]);
  assign t[201] = t[241] ^ t[212];
  assign t[202] = t[200] ? t[213] : t[244];
  assign t[203] = t[242] ^ t[214];
  assign t[204] = t[75] ? x[104] : x[103];
  assign t[205] = t[164] ? x[106] : x[105];
  assign t[206] = t[164] ? x[108] : x[107];
  assign t[207] = t[243] ^ t[215];
  assign t[208] = ~(t[211]);
  assign t[209] = ~(t[179]);
  assign t[20] = ~(t[222]);
  assign t[210] = t[128] ^ t[179];
  assign t[211] = t[183] ^ t[165];
  assign t[212] = t[216] ? x[110] : x[109];
  assign t[213] = t[244] ^ t[217];
  assign t[214] = t[216] ? x[112] : x[111];
  assign t[215] = t[216] ? x[114] : x[113];
  assign t[216] = ~(t[49]);
  assign t[217] = t[216] ? x[116] : x[115];
  assign t[218] = t[245] ^ x[4];
  assign t[219] = t[246] ^ x[7];
  assign t[21] = ~(t[32] & t[223]);
  assign t[220] = t[247] ^ x[10];
  assign t[221] = t[248] ^ x[13];
  assign t[222] = t[249] ^ x[18];
  assign t[223] = t[250] ^ x[21];
  assign t[224] = t[251] ^ x[24];
  assign t[225] = t[252] ^ x[27];
  assign t[226] = t[253] ^ x[30];
  assign t[227] = t[254] ^ x[33];
  assign t[228] = t[255] ^ x[36];
  assign t[229] = t[256] ^ x[39];
  assign t[22] = ~(t[33] ^ t[34]);
  assign t[230] = t[257] ^ x[42];
  assign t[231] = t[258] ^ x[45];
  assign t[232] = t[259] ^ x[48];
  assign t[233] = t[260] ^ x[51];
  assign t[234] = t[261] ^ x[54];
  assign t[235] = t[262] ^ x[57];
  assign t[236] = t[263] ^ x[60];
  assign t[237] = t[264] ^ x[65];
  assign t[238] = t[265] ^ x[70];
  assign t[239] = t[266] ^ x[73];
  assign t[23] = t[35] ^ t[36];
  assign t[240] = t[267] ^ x[76];
  assign t[241] = t[268] ^ x[87];
  assign t[242] = t[269] ^ x[90];
  assign t[243] = t[270] ^ x[99];
  assign t[244] = t[271] ^ x[102];
  assign t[245] = (x[2] & x[3]);
  assign t[246] = (x[5] & x[6]);
  assign t[247] = (x[8] & x[9]);
  assign t[248] = (x[11] & x[12]);
  assign t[249] = (x[16] & x[17]);
  assign t[24] = t[37] ^ t[38];
  assign t[250] = (x[19] & x[20]);
  assign t[251] = (x[22] & x[23]);
  assign t[252] = (x[25] & x[26]);
  assign t[253] = (x[28] & x[29]);
  assign t[254] = (x[31] & x[32]);
  assign t[255] = (x[34] & x[35]);
  assign t[256] = (x[37] & x[38]);
  assign t[257] = (x[40] & x[41]);
  assign t[258] = (x[43] & x[44]);
  assign t[259] = (x[46] & x[47]);
  assign t[25] = ~(t[39] ^ t[40]);
  assign t[260] = (x[49] & x[50]);
  assign t[261] = (x[52] & x[53]);
  assign t[262] = (x[55] & x[56]);
  assign t[263] = (x[58] & x[59]);
  assign t[264] = (x[63] & x[64]);
  assign t[265] = (x[68] & x[69]);
  assign t[266] = (x[71] & x[72]);
  assign t[267] = (x[74] & x[75]);
  assign t[268] = (x[85] & x[86]);
  assign t[269] = (x[88] & x[89]);
  assign t[26] = t[41] ^ t[42];
  assign t[270] = (x[97] & x[98]);
  assign t[271] = (x[100] & x[101]);
  assign t[27] = ~(t[43] ^ t[24]);
  assign t[28] = t[44] ^ t[45];
  assign t[29] = ~(t[35] ^ t[46]);
  assign t[2] = ~(t[6] ^ t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = ~(t[49]);
  assign t[32] = ~(t[224]);
  assign t[33] = t[50] ^ t[17];
  assign t[34] = ~(t[51] ^ t[43]);
  assign t[35] = t[52] ^ t[53];
  assign t[36] = ~(t[54] ^ t[55]);
  assign t[37] = ~t[56];
  assign t[38] = t[57] ^ t[58];
  assign t[39] = t[59] ^ t[60];
  assign t[3] = t[8] ? t[9] : t[218];
  assign t[40] = ~(t[41] ^ t[46]);
  assign t[41] = t[61] ^ t[62];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] ^ t[35]);
  assign t[44] = ~(t[66] ^ t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = t[70] ^ t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[225] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = ~(t[10] & t[11]);
  assign t[50] = t[76] ^ t[77];
  assign t[51] = t[78] ^ t[79];
  assign t[52] = t[80] ^ t[37];
  assign t[53] = t[57] ^ t[81];
  assign t[54] = t[82] ^ t[44];
  assign t[55] = ~(t[24] ^ t[83]);
  assign t[56] = t[8] ? t[84] : t[226];
  assign t[57] = t[85] ^ t[77];
  assign t[58] = t[86] & t[87];
  assign t[59] = t[24] ^ t[50];
  assign t[5] = ~(t[12] & t[13]);
  assign t[60] = ~(t[88] ^ t[89]);
  assign t[61] = t[90] ^ t[70];
  assign t[62] = t[91] & t[92];
  assign t[63] = t[93] ^ t[94];
  assign t[64] = t[95] ^ t[96];
  assign t[65] = ~(t[97] ^ t[98]);
  assign t[66] = t[99] ^ t[100];
  assign t[67] = ~(t[101] ^ t[102]);
  assign t[68] = t[103] ^ t[93];
  assign t[69] = t[104] & t[105];
  assign t[6] = ~(t[14] ^ t[15]);
  assign t[70] = t[8] ? t[106] : t[227];
  assign t[71] = t[107] ^ t[108];
  assign t[72] = ~(t[74] & t[109]);
  assign t[73] = ~(t[228] ^ t[110]);
  assign t[74] = ~(t[111] & t[112]);
  assign t[75] = ~(t[48]);
  assign t[76] = t[113] ^ t[37];
  assign t[77] = t[114] & t[115];
  assign t[78] = t[116] ^ t[70];
  assign t[79] = t[107] ^ t[117];
  assign t[7] = ~(t[16] ^ t[17]);
  assign t[80] = ~t[118];
  assign t[81] = t[119] & t[120];
  assign t[82] = ~(t[121] ^ t[122]);
  assign t[83] = t[123] ^ t[108];
  assign t[84] = t[226] ^ t[124];
  assign t[85] = t[125] & t[126];
  assign t[86] = ~(t[127] ^ t[57]);
  assign t[87] = t[52] ^ t[115];
  assign t[88] = ~(t[45] ^ t[102]);
  assign t[89] = t[128] ^ t[129];
  assign t[8] = ~(t[18]);
  assign t[90] = t[8] ? t[130] : t[229];
  assign t[91] = ~(t[116]);
  assign t[92] = t[8] ? t[131] : t[230];
  assign t[93] = t[30] ? t[132] : t[231];
  assign t[94] = t[30] ? t[133] : t[232];
  assign t[95] = t[134] ^ t[135];
  assign t[96] = t[136] & t[137];
  assign t[97] = t[51] ^ t[138];
  assign t[98] = t[139] ^ t[140];
  assign t[99] = t[141] ^ t[142];
  assign t[9] = t[218] ^ t[19];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind77(x, y);
 input [116:0] x;
 output y;

 wire [262:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[221] ^ t[143];
  assign t[101] = ~(t[113] ^ t[55]);
  assign t[102] = t[35] ^ t[123];
  assign t[103] = t[144] ? x[59] : x[58];
  assign t[104] = t[145] & t[146];
  assign t[105] = t[147] & t[148];
  assign t[106] = ~(t[90] ^ t[70]);
  assign t[107] = t[149] ^ t[148];
  assign t[108] = ~(t[150] & t[151]);
  assign t[109] = t[152] ^ t[227];
  assign t[10] = ~(t[210]);
  assign t[110] = ~(t[222]);
  assign t[111] = t[153] & t[152];
  assign t[112] = t[154] ^ t[60];
  assign t[113] = t[155] ^ t[54];
  assign t[114] = t[118] ^ t[156];
  assign t[115] = t[61] ^ t[157];
  assign t[116] = t[223] ^ t[158];
  assign t[117] = t[159] ^ t[42];
  assign t[118] = t[80] ^ t[64];
  assign t[119] = t[224] ^ t[160];
  assign t[11] = ~(t[211]);
  assign t[120] = ~(t[126]);
  assign t[121] = ~(t[155]);
  assign t[122] = ~(t[54]);
  assign t[123] = t[161];
  assign t[124] = t[35] ^ t[155];
  assign t[125] = t[155] ^ t[43];
  assign t[126] = t[123] ^ t[54];
  assign t[127] = ~(t[162] ^ t[163]);
  assign t[128] = t[164] ^ t[165];
  assign t[129] = t[8] ? t[166] : t[228];
  assign t[12] = ~(t[212]);
  assign t[130] = t[8] ? t[167] : t[229];
  assign t[131] = ~(t[18]);
  assign t[132] = t[225] ^ t[168];
  assign t[133] = t[226] ^ t[169];
  assign t[134] = ~(t[139]);
  assign t[135] = ~(t[154]);
  assign t[136] = ~(t[59]);
  assign t[137] = t[211] ^ t[170];
  assign t[138] = t[39] ^ t[154];
  assign t[139] = t[137] ^ t[59];
  assign t[13] = ~(t[20] | t[21]);
  assign t[140] = t[31] ? x[70] : x[69];
  assign t[141] = t[75] ? x[72] : x[71];
  assign t[142] = t[75] ? x[74] : x[73];
  assign t[143] = t[144] ? x[76] : x[75];
  assign t[144] = ~(t[49]);
  assign t[145] = ~(t[171]);
  assign t[146] = ~(t[129]);
  assign t[147] = ~(t[130]);
  assign t[148] = t[8] ? t[172] : t[230];
  assign t[149] = t[130] ^ t[45];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = ~(t[153] | t[152]);
  assign t[151] = ~(t[173] | t[110]);
  assign t[152] = ~(t[231]);
  assign t[153] = ~(t[227]);
  assign t[154] = t[131] ? t[174] : t[232];
  assign t[155] = t[175];
  assign t[156] = t[117] ^ t[176];
  assign t[157] = t[177] & t[178];
  assign t[158] = t[31] ? x[87] : x[86];
  assign t[159] = t[179] & t[180];
  assign t[15] = t[24] ^ t[25];
  assign t[160] = t[144] ? x[89] : x[88];
  assign t[161] = t[30] ? t[181] : t[233];
  assign t[162] = t[182] ^ t[183];
  assign t[163] = ~(t[184] ^ t[29]);
  assign t[164] = t[149] ^ t[185];
  assign t[165] = t[64] ^ t[186];
  assign t[166] = t[228] ^ t[187];
  assign t[167] = t[229] ^ t[188];
  assign t[168] = t[189] ? x[94] : x[93];
  assign t[169] = t[189] ? x[96] : x[95];
  assign t[16] = t[26] ^ t[27];
  assign t[170] = t[131] ? t[190] : t[234];
  assign t[171] = t[148] ^ t[130];
  assign t[172] = t[230] ^ t[191];
  assign t[173] = ~(t[217]);
  assign t[174] = t[232] ^ t[192];
  assign t[175] = t[8] ? t[193] : t[235];
  assign t[176] = t[194] & t[195];
  assign t[177] = ~(t[196] ^ t[61]);
  assign t[178] = t[39] ^ t[137];
  assign t[179] = ~(t[197]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[180] = ~(t[63]);
  assign t[181] = t[233] ^ t[198];
  assign t[182] = t[28] ^ t[199];
  assign t[183] = ~(t[200] ^ t[26]);
  assign t[184] = t[201] ^ t[105];
  assign t[185] = t[70] ^ t[202];
  assign t[186] = t[117] ^ t[53];
  assign t[187] = t[144] ? x[104] : x[103];
  assign t[188] = t[144] ? x[106] : x[105];
  assign t[189] = ~(t[49]);
  assign t[18] = ~(t[30]);
  assign t[190] = t[234] ^ t[203];
  assign t[191] = t[144] ? x[108] : x[107];
  assign t[192] = t[189] ? x[110] : x[109];
  assign t[193] = t[235] ^ t[204];
  assign t[194] = ~(t[159] ^ t[205]);
  assign t[195] = t[41] ^ t[197];
  assign t[196] = t[154] ^ t[59];
  assign t[197] = t[66] ^ t[80];
  assign t[198] = t[144] ? x[112] : x[111];
  assign t[199] = t[125] ^ t[85];
  assign t[19] = t[31] ? x[15] : x[14];
  assign t[1] = ~(t[4] | t[5]);
  assign t[200] = ~(t[34] ^ t[79]);
  assign t[201] = t[129] ^ t[45];
  assign t[202] = t[206] & t[207];
  assign t[203] = t[189] ? x[114] : x[113];
  assign t[204] = t[144] ? x[116] : x[115];
  assign t[205] = t[118] ^ t[63];
  assign t[206] = ~(t[104] ^ t[208]);
  assign t[207] = t[201] ^ t[171];
  assign t[208] = t[149] ^ t[129];
  assign t[209] = t[236] ^ x[4];
  assign t[20] = ~(t[213]);
  assign t[210] = t[237] ^ x[7];
  assign t[211] = t[238] ^ x[10];
  assign t[212] = t[239] ^ x[13];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[32] & t[214]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[62];
  assign t[228] = t[255] ^ x[65];
  assign t[229] = t[256] ^ x[68];
  assign t[22] = t[33] ^ t[34];
  assign t[230] = t[257] ^ x[79];
  assign t[231] = t[258] ^ x[82];
  assign t[232] = t[259] ^ x[85];
  assign t[233] = t[260] ^ x[92];
  assign t[234] = t[261] ^ x[99];
  assign t[235] = t[262] ^ x[102];
  assign t[236] = (x[2] & x[3]);
  assign t[237] = (x[5] & x[6]);
  assign t[238] = (x[8] & x[9]);
  assign t[239] = (x[11] & x[12]);
  assign t[23] = ~(t[24] ^ t[29]);
  assign t[240] = (x[16] & x[17]);
  assign t[241] = (x[19] & x[20]);
  assign t[242] = (x[22] & x[23]);
  assign t[243] = (x[25] & x[26]);
  assign t[244] = (x[28] & x[29]);
  assign t[245] = (x[31] & x[32]);
  assign t[246] = (x[34] & x[35]);
  assign t[247] = (x[37] & x[38]);
  assign t[248] = (x[40] & x[41]);
  assign t[249] = (x[43] & x[44]);
  assign t[24] = t[35] ^ t[36];
  assign t[250] = (x[46] & x[47]);
  assign t[251] = (x[49] & x[50]);
  assign t[252] = (x[52] & x[53]);
  assign t[253] = (x[55] & x[56]);
  assign t[254] = (x[60] & x[61]);
  assign t[255] = (x[63] & x[64]);
  assign t[256] = (x[66] & x[67]);
  assign t[257] = (x[77] & x[78]);
  assign t[258] = (x[80] & x[81]);
  assign t[259] = (x[83] & x[84]);
  assign t[25] = ~(t[37] ^ t[38]);
  assign t[260] = (x[90] & x[91]);
  assign t[261] = (x[97] & x[98]);
  assign t[262] = (x[100] & x[101]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = t[41] ^ t[42];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[6] ^ t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = ~(t[49]);
  assign t[32] = ~(t[215]);
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[34] = t[52] ^ t[53];
  assign t[35] = t[54] ^ t[43];
  assign t[36] = t[55] ^ t[56];
  assign t[37] = t[57] ^ t[33];
  assign t[38] = ~(t[28] ^ t[58]);
  assign t[39] = t[59] ^ t[60];
  assign t[3] = t[8] ? t[9] : t[209];
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = ~t[67];
  assign t[44] = t[55] ^ t[68];
  assign t[45] = t[8] ? t[69] : t[216];
  assign t[46] = t[70] ^ t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[217] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = ~(t[10] & t[11]);
  assign t[50] = t[76] ^ t[77];
  assign t[51] = ~(t[78] ^ t[79]);
  assign t[52] = t[63] ^ t[80];
  assign t[53] = t[81] & t[82];
  assign t[54] = ~t[83];
  assign t[55] = t[84] ^ t[85];
  assign t[56] = t[86] & t[87];
  assign t[57] = ~(t[88] ^ t[89]);
  assign t[58] = t[90] ^ t[71];
  assign t[59] = t[210] ^ t[91];
  assign t[5] = ~(t[12] & t[13]);
  assign t[60] = t[214] ^ t[92];
  assign t[61] = t[93] ^ t[94];
  assign t[62] = t[95] & t[96];
  assign t[63] = t[30] ? t[97] : t[218];
  assign t[64] = t[30] ? t[98] : t[219];
  assign t[65] = ~(t[80]);
  assign t[66] = t[30] ? t[99] : t[220];
  assign t[67] = t[8] ? t[100] : t[221];
  assign t[68] = t[101] & t[102];
  assign t[69] = t[216] ^ t[103];
  assign t[6] = ~(t[14] ^ t[15]);
  assign t[70] = t[104] ^ t[105];
  assign t[71] = t[106] & t[107];
  assign t[72] = ~(t[74] & t[108]);
  assign t[73] = ~(t[222] ^ t[109]);
  assign t[74] = ~(t[110] & t[111]);
  assign t[75] = ~(t[48]);
  assign t[76] = t[112] ^ t[94];
  assign t[77] = t[113] ^ t[68];
  assign t[78] = t[114] ^ t[58];
  assign t[79] = t[60] ^ t[115];
  assign t[7] = ~(t[16] ^ t[17]);
  assign t[80] = t[30] ? t[116] : t[223];
  assign t[81] = ~(t[52] ^ t[117]);
  assign t[82] = t[118] ^ t[66];
  assign t[83] = t[8] ? t[119] : t[224];
  assign t[84] = t[120] & t[121];
  assign t[85] = t[122] & t[123];
  assign t[86] = ~(t[84] ^ t[124]);
  assign t[87] = t[125] ^ t[126];
  assign t[88] = t[127] ^ t[27];
  assign t[89] = ~(t[128] ^ t[77]);
  assign t[8] = ~(t[18]);
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[131] ? t[132] : t[225];
  assign t[92] = t[131] ? t[133] : t[226];
  assign t[93] = t[134] & t[135];
  assign t[94] = t[136] & t[137];
  assign t[95] = ~(t[93] ^ t[138]);
  assign t[96] = t[112] ^ t[139];
  assign t[97] = t[218] ^ t[140];
  assign t[98] = t[219] ^ t[141];
  assign t[99] = t[220] ^ t[142];
  assign t[9] = t[209] ^ t[19];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind78(x, y);
 input [116:0] x;
 output y;

 wire [260:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[218] ^ t[140];
  assign t[101] = ~(t[141] & t[142]);
  assign t[102] = t[143] ^ t[221];
  assign t[103] = ~(t[219]);
  assign t[104] = t[144] & t[143];
  assign t[105] = t[84] ^ t[124];
  assign t[106] = t[145] & t[146];
  assign t[107] = t[147];
  assign t[108] = t[109] ^ t[60];
  assign t[109] = t[148] ^ t[149];
  assign t[10] = ~(t[208]);
  assign t[110] = t[150] & t[151];
  assign t[111] = t[152] ? t[153] : t[222];
  assign t[112] = t[154] ^ t[57];
  assign t[113] = t[124] ^ t[75];
  assign t[114] = t[112] ^ t[155];
  assign t[115] = t[156] ^ t[126];
  assign t[116] = t[157] & t[158];
  assign t[117] = t[61] ^ t[159];
  assign t[118] = t[137] ^ t[95];
  assign t[119] = t[156] ^ t[121];
  assign t[11] = ~(t[209]);
  assign t[120] = t[160] & t[161];
  assign t[121] = t[8] ? t[162] : t[223];
  assign t[122] = t[127] ^ t[116];
  assign t[123] = t[220] ^ t[163];
  assign t[124] = t[210] ^ t[164];
  assign t[125] = t[30] ? t[165] : t[224];
  assign t[126] = t[8] ? t[166] : t[225];
  assign t[127] = t[167] ^ t[120];
  assign t[128] = t[168] & t[169];
  assign t[129] = t[30] ? t[170] : t[226];
  assign t[12] = ~(t[210]);
  assign t[130] = t[30] ? t[171] : t[227];
  assign t[131] = t[172];
  assign t[132] = t[139] ? x[72] : x[71];
  assign t[133] = ~(t[138]);
  assign t[134] = ~(t[42]);
  assign t[135] = ~(t[43]);
  assign t[136] = t[40] ^ t[42];
  assign t[137] = t[42] ^ t[61];
  assign t[138] = t[66] ^ t[43];
  assign t[139] = ~(t[48]);
  assign t[13] = ~(t[20] | t[21]);
  assign t[140] = t[139] ? x[74] : x[73];
  assign t[141] = ~(t[144] | t[143]);
  assign t[142] = ~(t[173] | t[103]);
  assign t[143] = ~(t[228]);
  assign t[144] = ~(t[221]);
  assign t[145] = ~(t[105] ^ t[112]);
  assign t[146] = t[113] ^ t[86];
  assign t[147] = t[30] ? t[174] : t[229];
  assign t[148] = t[175] & t[176];
  assign t[149] = t[177] & t[131];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = ~(t[148] ^ t[178]);
  assign t[151] = t[179] ^ t[180];
  assign t[152] = ~(t[18]);
  assign t[153] = t[222] ^ t[181];
  assign t[154] = t[182] & t[183];
  assign t[155] = t[184] & t[185];
  assign t[156] = t[8] ? t[186] : t[230];
  assign t[157] = ~(t[115] ^ t[127]);
  assign t[158] = t[87] ^ t[161];
  assign t[159] = t[62] ^ t[29];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[126]);
  assign t[161] = t[8] ? t[187] : t[231];
  assign t[162] = t[223] ^ t[188];
  assign t[163] = t[139] ? x[88] : x[87];
  assign t[164] = t[30] ? t[189] : t[232];
  assign t[165] = t[224] ^ t[190];
  assign t[166] = t[225] ^ t[191];
  assign t[167] = t[192] & t[193];
  assign t[168] = ~(t[167] ^ t[194]);
  assign t[169] = t[119] ^ t[195];
  assign t[16] = ~(t[26] ^ t[27]);
  assign t[170] = t[226] ^ t[196];
  assign t[171] = t[227] ^ t[197];
  assign t[172] = t[30] ? t[198] : t[233];
  assign t[173] = ~(t[216]);
  assign t[174] = t[229] ^ t[199];
  assign t[175] = ~(t[180]);
  assign t[176] = ~(t[89]);
  assign t[177] = ~(t[90]);
  assign t[178] = t[73] ^ t[89];
  assign t[179] = t[89] ^ t[107];
  assign t[17] = t[28] ^ t[29];
  assign t[180] = t[131] ^ t[90];
  assign t[181] = t[200] ? x[96] : x[95];
  assign t[182] = ~(t[201]);
  assign t[183] = ~(t[84]);
  assign t[184] = ~(t[154] ^ t[202]);
  assign t[185] = t[56] ^ t[201];
  assign t[186] = t[230] ^ t[203];
  assign t[187] = t[231] ^ t[204];
  assign t[188] = t[31] ? x[98] : x[97];
  assign t[189] = t[232] ^ t[205];
  assign t[18] = ~(t[30]);
  assign t[190] = t[70] ? x[100] : x[99];
  assign t[191] = t[31] ? x[102] : x[101];
  assign t[192] = ~(t[195]);
  assign t[193] = ~(t[156]);
  assign t[194] = t[87] ^ t[156];
  assign t[195] = t[161] ^ t[126];
  assign t[196] = t[70] ? x[104] : x[103];
  assign t[197] = t[200] ? x[106] : x[105];
  assign t[198] = t[233] ^ t[206];
  assign t[199] = t[70] ? x[108] : x[107];
  assign t[19] = t[31] ? x[15] : x[14];
  assign t[1] = ~(t[4] | t[5]);
  assign t[200] = ~(t[48]);
  assign t[201] = t[86] ^ t[124];
  assign t[202] = t[113] ^ t[84];
  assign t[203] = t[31] ? x[110] : x[109];
  assign t[204] = t[31] ? x[112] : x[111];
  assign t[205] = t[139] ? x[114] : x[113];
  assign t[206] = t[200] ? x[116] : x[115];
  assign t[207] = t[234] ^ x[4];
  assign t[208] = t[235] ^ x[7];
  assign t[209] = t[236] ^ x[10];
  assign t[20] = ~(t[211]);
  assign t[210] = t[237] ^ x[13];
  assign t[211] = t[238] ^ x[18];
  assign t[212] = t[239] ^ x[21];
  assign t[213] = t[240] ^ x[24];
  assign t[214] = t[241] ^ x[27];
  assign t[215] = t[242] ^ x[30];
  assign t[216] = t[243] ^ x[33];
  assign t[217] = t[244] ^ x[36];
  assign t[218] = t[245] ^ x[39];
  assign t[219] = t[246] ^ x[42];
  assign t[21] = ~(t[32] & t[212]);
  assign t[220] = t[247] ^ x[45];
  assign t[221] = t[248] ^ x[52];
  assign t[222] = t[249] ^ x[55];
  assign t[223] = t[250] ^ x[58];
  assign t[224] = t[251] ^ x[61];
  assign t[225] = t[252] ^ x[64];
  assign t[226] = t[253] ^ x[67];
  assign t[227] = t[254] ^ x[70];
  assign t[228] = t[255] ^ x[77];
  assign t[229] = t[256] ^ x[80];
  assign t[22] = ~(t[27] ^ t[33]);
  assign t[230] = t[257] ^ x[83];
  assign t[231] = t[258] ^ x[86];
  assign t[232] = t[259] ^ x[91];
  assign t[233] = t[260] ^ x[94];
  assign t[234] = (x[2] & x[3]);
  assign t[235] = (x[5] & x[6]);
  assign t[236] = (x[8] & x[9]);
  assign t[237] = (x[11] & x[12]);
  assign t[238] = (x[16] & x[17]);
  assign t[239] = (x[19] & x[20]);
  assign t[23] = ~(t[34] ^ t[35]);
  assign t[240] = (x[22] & x[23]);
  assign t[241] = (x[25] & x[26]);
  assign t[242] = (x[28] & x[29]);
  assign t[243] = (x[31] & x[32]);
  assign t[244] = (x[34] & x[35]);
  assign t[245] = (x[37] & x[38]);
  assign t[246] = (x[40] & x[41]);
  assign t[247] = (x[43] & x[44]);
  assign t[248] = (x[50] & x[51]);
  assign t[249] = (x[53] & x[54]);
  assign t[24] = t[36] ^ t[37];
  assign t[250] = (x[56] & x[57]);
  assign t[251] = (x[59] & x[60]);
  assign t[252] = (x[62] & x[63]);
  assign t[253] = (x[65] & x[66]);
  assign t[254] = (x[68] & x[69]);
  assign t[255] = (x[75] & x[76]);
  assign t[256] = (x[78] & x[79]);
  assign t[257] = (x[81] & x[82]);
  assign t[258] = (x[84] & x[85]);
  assign t[259] = (x[89] & x[90]);
  assign t[25] = ~(t[38] ^ t[17]);
  assign t[260] = (x[92] & x[93]);
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[27] = t[40] ^ t[41];
  assign t[28] = t[42] ^ t[43];
  assign t[29] = t[44] & t[45];
  assign t[2] = ~(t[6] ^ t[7]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[31] = ~(t[48]);
  assign t[32] = ~(t[213]);
  assign t[33] = ~(t[49] ^ t[50]);
  assign t[34] = ~(t[51] ^ t[52]);
  assign t[35] = t[16] ^ t[53];
  assign t[36] = ~(t[54] ^ t[55]);
  assign t[37] = t[56] ^ t[57];
  assign t[38] = t[58] ^ t[51];
  assign t[39] = t[59] ^ t[60];
  assign t[3] = t[8] ? t[9] : t[207];
  assign t[40] = t[43] ^ t[61];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[8] ? t[64] : t[214];
  assign t[43] = t[8] ? t[65] : t[215];
  assign t[44] = ~(t[28] ^ t[62]);
  assign t[45] = t[40] ^ t[66];
  assign t[46] = ~(t[67] & t[68]);
  assign t[47] = t[216] | t[69];
  assign t[48] = ~(t[70]);
  assign t[49] = ~(t[71] ^ t[72]);
  assign t[4] = ~(t[10] & t[11]);
  assign t[50] = t[73] ^ t[74];
  assign t[51] = t[75] ^ t[76];
  assign t[52] = t[77] ^ t[78];
  assign t[53] = ~(t[79] ^ t[80]);
  assign t[54] = t[81] ^ t[33];
  assign t[55] = ~(t[82] ^ t[83]);
  assign t[56] = t[84] ^ t[75];
  assign t[57] = t[85] & t[86];
  assign t[58] = t[87] ^ t[88];
  assign t[59] = t[89] ^ t[90];
  assign t[5] = ~(t[12] & t[13]);
  assign t[60] = t[91] & t[92];
  assign t[61] = t[8] ? t[93] : t[217];
  assign t[62] = t[94] ^ t[95];
  assign t[63] = t[96] & t[97];
  assign t[64] = t[214] ^ t[98];
  assign t[65] = t[215] ^ t[99];
  assign t[66] = t[8] ? t[100] : t[218];
  assign t[67] = ~(t[69] & t[101]);
  assign t[68] = ~(t[219] ^ t[102]);
  assign t[69] = ~(t[103] & t[104]);
  assign t[6] = t[14] ^ t[15];
  assign t[70] = ~(t[47]);
  assign t[71] = t[105] ^ t[106];
  assign t[72] = t[107] ^ t[108];
  assign t[73] = t[90] ^ t[107];
  assign t[74] = t[109] ^ t[110];
  assign t[75] = t[211] ^ t[111];
  assign t[76] = t[112] ^ t[106];
  assign t[77] = t[113] ^ t[114];
  assign t[78] = t[115] ^ t[116];
  assign t[79] = t[50] ^ t[37];
  assign t[7] = ~(t[16] ^ t[17]);
  assign t[80] = ~(t[117] ^ t[83]);
  assign t[81] = t[117] ^ t[118];
  assign t[82] = t[119] ^ t[120];
  assign t[83] = t[121] ^ t[122];
  assign t[84] = t[30] ? t[123] : t[220];
  assign t[85] = ~(t[124]);
  assign t[86] = t[213] ^ t[125];
  assign t[87] = t[126] ^ t[121];
  assign t[88] = t[127] ^ t[128];
  assign t[89] = ~t[129];
  assign t[8] = ~(t[18]);
  assign t[90] = t[130];
  assign t[91] = ~(t[59] ^ t[109]);
  assign t[92] = t[73] ^ t[131];
  assign t[93] = t[217] ^ t[132];
  assign t[94] = t[133] & t[134];
  assign t[95] = t[135] & t[66];
  assign t[96] = ~(t[94] ^ t[136]);
  assign t[97] = t[137] ^ t[138];
  assign t[98] = t[139] ? x[47] : x[46];
  assign t[99] = t[139] ? x[49] : x[48];
  assign t[9] = t[207] ^ t[19];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind79(x, y);
 input [116:0] x;
 output y;

 wire [262:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[119] ^ t[137];
  assign t[101] = t[138] ^ t[139];
  assign t[102] = t[140] ^ t[133];
  assign t[103] = t[106] ? t[141] : t[225];
  assign t[104] = t[142] ^ t[109];
  assign t[105] = t[143] & t[144];
  assign t[106] = ~(t[145]);
  assign t[107] = t[219] ^ t[146];
  assign t[108] = t[123] ^ t[70];
  assign t[109] = t[147] & t[148];
  assign t[10] = ~(t[210]);
  assign t[110] = t[106] ? t[149] : t[226];
  assign t[111] = t[119] ^ t[57];
  assign t[112] = t[150] ^ t[121];
  assign t[113] = ~(t[213]);
  assign t[114] = t[8] ? t[151] : t[227];
  assign t[115] = t[152];
  assign t[116] = t[8] ? t[153] : t[228];
  assign t[117] = t[221] ^ t[154];
  assign t[118] = t[222] ^ t[155];
  assign t[119] = t[156] ^ t[157];
  assign t[11] = ~(t[211]);
  assign t[120] = t[106] ? t[158] : t[229];
  assign t[121] = t[212] ^ t[159];
  assign t[122] = t[160] & t[161];
  assign t[123] = t[106] ? t[162] : t[230];
  assign t[124] = ~(t[89] ^ t[104]);
  assign t[125] = t[68] ^ t[148];
  assign t[126] = t[223] ^ t[163];
  assign t[127] = t[164] & t[165];
  assign t[128] = ~(t[136] ^ t[92]);
  assign t[129] = t[138] ^ t[82];
  assign t[12] = ~(t[212]);
  assign t[130] = ~(t[145]);
  assign t[131] = t[224] ^ t[166];
  assign t[132] = t[167] & t[168];
  assign t[133] = t[169] & t[170];
  assign t[134] = ~(t[112] ^ t[95]);
  assign t[135] = t[87] ^ t[170];
  assign t[136] = t[80] ^ t[115];
  assign t[137] = t[171] & t[172];
  assign t[138] = t[115] ^ t[60];
  assign t[139] = t[92] ^ t[173];
  assign t[13] = ~(t[21] | t[22]);
  assign t[140] = t[150] ^ t[62];
  assign t[141] = t[225] ^ t[174];
  assign t[142] = t[175] & t[176];
  assign t[143] = ~(t[142] ^ t[177]);
  assign t[144] = t[108] ^ t[178];
  assign t[145] = ~(t[8]);
  assign t[146] = t[34] ? x[71] : x[70];
  assign t[147] = ~(t[103]);
  assign t[148] = t[106] ? t[179] : t[231];
  assign t[149] = t[226] ^ t[180];
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = t[8] ? t[181] : t[232];
  assign t[151] = t[227] ^ t[182];
  assign t[152] = t[8] ? t[183] : t[233];
  assign t[153] = t[228] ^ t[184];
  assign t[154] = t[185] ? x[82] : x[81];
  assign t[155] = t[185] ? x[84] : x[83];
  assign t[156] = t[186] & t[187];
  assign t[157] = t[188] & t[120];
  assign t[158] = t[229] ^ t[189];
  assign t[159] = t[8] ? t[190] : t[234];
  assign t[15] = ~(t[25] ^ t[26]);
  assign t[160] = ~(t[132] ^ t[191]);
  assign t[161] = t[140] ^ t[192];
  assign t[162] = t[230] ^ t[193];
  assign t[163] = t[79] ? x[89] : x[88];
  assign t[164] = ~(t[194]);
  assign t[165] = ~(t[80]);
  assign t[166] = t[195] ? x[91] : x[90];
  assign t[167] = ~(t[192]);
  assign t[168] = ~(t[150]);
  assign t[169] = ~(t[121]);
  assign t[16] = ~(t[27] ^ t[28]);
  assign t[170] = t[217] ^ t[196];
  assign t[171] = ~(t[156] ^ t[197]);
  assign t[172] = t[198] ^ t[199];
  assign t[173] = t[200] & t[201];
  assign t[174] = t[34] ? x[93] : x[92];
  assign t[175] = ~(t[178]);
  assign t[176] = ~(t[123]);
  assign t[177] = t[68] ^ t[123];
  assign t[178] = t[148] ^ t[103];
  assign t[179] = t[231] ^ t[202];
  assign t[17] = ~(t[29] ^ t[30]);
  assign t[180] = t[185] ? x[95] : x[94];
  assign t[181] = t[232] ^ t[203];
  assign t[182] = t[79] ? x[97] : x[96];
  assign t[183] = t[233] ^ t[204];
  assign t[184] = t[195] ? x[99] : x[98];
  assign t[185] = ~(t[53]);
  assign t[186] = ~(t[199]);
  assign t[187] = ~(t[83]);
  assign t[188] = ~(t[84]);
  assign t[189] = t[185] ? x[101] : x[100];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[234] ^ t[205];
  assign t[191] = t[87] ^ t[150];
  assign t[192] = t[170] ^ t[121];
  assign t[193] = t[34] ? x[103] : x[102];
  assign t[194] = t[82] ^ t[115];
  assign t[195] = ~(t[53]);
  assign t[196] = t[8] ? t[206] : t[235];
  assign t[197] = t[99] ^ t[83];
  assign t[198] = t[83] ^ t[110];
  assign t[199] = t[120] ^ t[84];
  assign t[19] = t[213] | t[33];
  assign t[1] = ~(t[4] | t[5]);
  assign t[200] = ~(t[127] ^ t[207]);
  assign t[201] = t[54] ^ t[194];
  assign t[202] = t[34] ? x[108] : x[107];
  assign t[203] = t[185] ? x[110] : x[109];
  assign t[204] = t[195] ? x[112] : x[111];
  assign t[205] = t[185] ? x[114] : x[113];
  assign t[206] = t[235] ^ t[208];
  assign t[207] = t[138] ^ t[80];
  assign t[208] = t[79] ? x[116] : x[115];
  assign t[209] = t[236] ^ x[4];
  assign t[20] = t[34] ? x[18] : x[17];
  assign t[210] = t[237] ^ x[7];
  assign t[211] = t[238] ^ x[10];
  assign t[212] = t[239] ^ x[13];
  assign t[213] = t[240] ^ x[16];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[214]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[60];
  assign t[228] = t[255] ^ x[63];
  assign t[229] = t[256] ^ x[66];
  assign t[22] = ~(t[35] & t[215]);
  assign t[230] = t[257] ^ x[69];
  assign t[231] = t[258] ^ x[74];
  assign t[232] = t[259] ^ x[77];
  assign t[233] = t[260] ^ x[80];
  assign t[234] = t[261] ^ x[87];
  assign t[235] = t[262] ^ x[106];
  assign t[236] = (x[2] & x[3]);
  assign t[237] = (x[5] & x[6]);
  assign t[238] = (x[8] & x[9]);
  assign t[239] = (x[11] & x[12]);
  assign t[23] = t[36] ^ t[37];
  assign t[240] = (x[14] & x[15]);
  assign t[241] = (x[19] & x[20]);
  assign t[242] = (x[22] & x[23]);
  assign t[243] = (x[25] & x[26]);
  assign t[244] = (x[28] & x[29]);
  assign t[245] = (x[31] & x[32]);
  assign t[246] = (x[34] & x[35]);
  assign t[247] = (x[37] & x[38]);
  assign t[248] = (x[40] & x[41]);
  assign t[249] = (x[43] & x[44]);
  assign t[24] = ~(t[38] ^ t[39]);
  assign t[250] = (x[46] & x[47]);
  assign t[251] = (x[49] & x[50]);
  assign t[252] = (x[52] & x[53]);
  assign t[253] = (x[55] & x[56]);
  assign t[254] = (x[58] & x[59]);
  assign t[255] = (x[61] & x[62]);
  assign t[256] = (x[64] & x[65]);
  assign t[257] = (x[67] & x[68]);
  assign t[258] = (x[72] & x[73]);
  assign t[259] = (x[75] & x[76]);
  assign t[25] = ~(t[40] ^ t[38]);
  assign t[260] = (x[78] & x[79]);
  assign t[261] = (x[85] & x[86]);
  assign t[262] = (x[104] & x[105]);
  assign t[26] = t[41] ^ t[42];
  assign t[27] = t[26] ^ t[37];
  assign t[28] = ~(t[43] ^ t[44]);
  assign t[29] = ~(t[45] ^ t[46]);
  assign t[2] = ~(t[6] ^ t[7]);
  assign t[30] = ~(t[47] ^ t[48]);
  assign t[31] = ~(t[33] & t[49]);
  assign t[32] = ~(t[216] ^ t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = ~(t[53]);
  assign t[35] = ~(t[217]);
  assign t[36] = t[54] ^ t[55];
  assign t[37] = t[56] ^ t[57];
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[60] ^ t[61];
  assign t[3] = t[8] ? t[9] : t[209];
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[64] ^ t[65]);
  assign t[42] = ~(t[66] ^ t[67]);
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = t[72] ^ t[58];
  assign t[46] = ~(t[41] ^ t[73]);
  assign t[47] = t[14] ^ t[74];
  assign t[48] = ~(t[65] ^ t[44]);
  assign t[49] = ~(t[75] & t[76]);
  assign t[4] = ~(t[10] & t[11]);
  assign t[50] = t[77] ^ t[218];
  assign t[51] = ~(t[216]);
  assign t[52] = t[78] & t[77];
  assign t[53] = ~(t[79]);
  assign t[54] = t[80] ^ t[60];
  assign t[55] = t[81] & t[82];
  assign t[56] = t[83] ^ t[84];
  assign t[57] = t[85] & t[86];
  assign t[58] = t[87] ^ t[88];
  assign t[59] = t[89] ^ t[90];
  assign t[5] = ~(t[12] & t[13]);
  assign t[60] = t[91];
  assign t[61] = t[92] ^ t[93];
  assign t[62] = t[214] ^ t[94];
  assign t[63] = t[95] ^ t[96];
  assign t[64] = ~(t[97] ^ t[98]);
  assign t[65] = t[99] ^ t[100];
  assign t[66] = t[101] ^ t[102];
  assign t[67] = ~(t[73] ^ t[44]);
  assign t[68] = t[103] ^ t[70];
  assign t[69] = t[104] ^ t[105];
  assign t[6] = ~(t[14] ^ t[15]);
  assign t[70] = t[106] ? t[107] : t[219];
  assign t[71] = t[104] ^ t[90];
  assign t[72] = t[108] ^ t[109];
  assign t[73] = t[110] ^ t[111];
  assign t[74] = t[112] ^ t[96];
  assign t[75] = ~(t[78] | t[77]);
  assign t[76] = ~(t[113] | t[51]);
  assign t[77] = ~(t[220]);
  assign t[78] = ~(t[218]);
  assign t[79] = ~(t[19]);
  assign t[7] = ~(t[16] ^ t[17]);
  assign t[80] = ~t[114];
  assign t[81] = ~(t[115]);
  assign t[82] = t[116];
  assign t[83] = t[106] ? t[117] : t[221];
  assign t[84] = t[106] ? t[118] : t[222];
  assign t[85] = ~(t[56] ^ t[119]);
  assign t[86] = t[99] ^ t[120];
  assign t[87] = t[121] ^ t[62];
  assign t[88] = t[95] ^ t[122];
  assign t[89] = t[123] ^ t[103];
  assign t[8] = ~(t[18] & t[19]);
  assign t[90] = t[124] & t[125];
  assign t[91] = t[8] ? t[126] : t[223];
  assign t[92] = t[127] ^ t[55];
  assign t[93] = t[128] & t[129];
  assign t[94] = t[130] ? t[131] : t[224];
  assign t[95] = t[132] ^ t[133];
  assign t[96] = t[134] & t[135];
  assign t[97] = t[43] ^ t[40];
  assign t[98] = t[136] ^ t[93];
  assign t[99] = t[84] ^ t[110];
  assign t[9] = t[209] ^ t[20];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind80(x, y);
 input [116:0] x;
 output y;

 wire [271:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[127] ^ t[58];
  assign t[101] = t[42] ^ t[83];
  assign t[102] = t[143] ^ t[144];
  assign t[103] = t[30] ? t[145] : t[232];
  assign t[104] = ~(t[68] ^ t[95]);
  assign t[105] = t[63] ^ t[146];
  assign t[106] = t[227] ^ t[147];
  assign t[107] = t[148] ^ t[62];
  assign t[108] = t[149] & t[150];
  assign t[109] = ~(t[151] & t[152]);
  assign t[10] = ~(t[219]);
  assign t[110] = t[153] ^ t[233];
  assign t[111] = ~(t[228]);
  assign t[112] = t[154] & t[153];
  assign t[113] = t[8] ? t[155] : t[234];
  assign t[114] = ~(t[80]);
  assign t[115] = t[8] ? t[156] : t[235];
  assign t[116] = t[8] ? t[157] : t[236];
  assign t[117] = t[158] & t[159];
  assign t[118] = t[229] ^ t[160];
  assign t[119] = ~(t[85] ^ t[161]);
  assign t[11] = ~(t[220]);
  assign t[120] = t[76] ^ t[162];
  assign t[121] = t[25] ^ t[163];
  assign t[122] = ~(t[97] ^ t[100]);
  assign t[123] = t[90] ^ t[116];
  assign t[124] = ~(t[49]);
  assign t[125] = ~(t[162]);
  assign t[126] = ~(t[113]);
  assign t[127] = t[113] ^ t[80];
  assign t[128] = t[164] ^ t[143];
  assign t[129] = t[165] ^ t[166];
  assign t[12] = ~(t[221]);
  assign t[130] = t[230] ^ t[167];
  assign t[131] = t[231] ^ t[168];
  assign t[132] = t[30] ? t[169] : t[237];
  assign t[133] = t[170] ? t[171] : t[238];
  assign t[134] = t[172] & t[173];
  assign t[135] = t[174] & t[146];
  assign t[136] = ~(t[134] ^ t[175]);
  assign t[137] = t[176] ^ t[177];
  assign t[138] = t[94] ^ t[178];
  assign t[139] = t[179] ^ t[164];
  assign t[13] = ~(t[20] | t[21]);
  assign t[140] = t[180] & t[181];
  assign t[141] = t[179] ^ t[143];
  assign t[142] = t[182] & t[183];
  assign t[143] = t[184];
  assign t[144] = t[165] ^ t[140];
  assign t[145] = t[232] ^ t[185];
  assign t[146] = t[224] ^ t[186];
  assign t[147] = t[31] ? x[70] : x[69];
  assign t[148] = t[187] & t[188];
  assign t[149] = ~(t[123] ^ t[107]);
  assign t[14] = t[22] ^ t[23];
  assign t[150] = t[78] ^ t[92];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[189] | t[111]);
  assign t[153] = ~(t[239]);
  assign t[154] = ~(t[233]);
  assign t[155] = t[234] ^ t[190];
  assign t[156] = t[235] ^ t[191];
  assign t[157] = t[236] ^ t[192];
  assign t[158] = ~(t[148] ^ t[193]);
  assign t[159] = t[61] ^ t[194];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = t[124] ? x[75] : x[74];
  assign t[161] = t[52] ^ t[113];
  assign t[162] = t[115] ^ t[80];
  assign t[163] = t[176] ^ t[135];
  assign t[164] = t[195];
  assign t[165] = t[196] ^ t[142];
  assign t[166] = t[197] & t[198];
  assign t[167] = t[31] ? x[77] : x[76];
  assign t[168] = t[31] ? x[79] : x[78];
  assign t[169] = t[237] ^ t[199];
  assign t[16] = ~(t[26] ^ t[27]);
  assign t[170] = ~(t[18]);
  assign t[171] = t[238] ^ t[200];
  assign t[172] = ~(t[177]);
  assign t[173] = ~(t[103]);
  assign t[174] = ~(t[93]);
  assign t[175] = t[63] ^ t[103];
  assign t[176] = t[103] ^ t[94];
  assign t[177] = t[146] ^ t[93];
  assign t[178] = t[95] ^ t[69];
  assign t[179] = ~t[201];
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[180] = ~(t[139] ^ t[165]);
  assign t[181] = t[128] ^ t[183];
  assign t[182] = ~(t[164]);
  assign t[183] = t[202];
  assign t[184] = t[30] ? t[203] : t[240];
  assign t[185] = t[124] ? x[84] : x[83];
  assign t[186] = t[30] ? t[204] : t[241];
  assign t[187] = ~(t[194]);
  assign t[188] = ~(t[90]);
  assign t[189] = ~(t[226]);
  assign t[18] = ~(t[30]);
  assign t[190] = t[124] ? x[89] : x[88];
  assign t[191] = t[124] ? x[91] : x[90];
  assign t[192] = t[31] ? x[93] : x[92];
  assign t[193] = t[78] ^ t[90];
  assign t[194] = t[92] ^ t[116];
  assign t[195] = t[30] ? t[205] : t[242];
  assign t[196] = t[206] & t[207];
  assign t[197] = ~(t[196] ^ t[208]);
  assign t[198] = t[141] ^ t[209];
  assign t[199] = t[124] ? x[98] : x[97];
  assign t[19] = t[31] ? x[15] : x[14];
  assign t[1] = ~(t[4] | t[5]);
  assign t[200] = t[210] ? x[100] : x[99];
  assign t[201] = t[30] ? t[211] : t[243];
  assign t[202] = t[30] ? t[212] : t[244];
  assign t[203] = t[240] ^ t[213];
  assign t[204] = t[241] ^ t[214];
  assign t[205] = t[242] ^ t[215];
  assign t[206] = ~(t[209]);
  assign t[207] = ~(t[179]);
  assign t[208] = t[128] ^ t[179];
  assign t[209] = t[183] ^ t[164];
  assign t[20] = ~(t[222]);
  assign t[210] = ~(t[49]);
  assign t[211] = t[243] ^ t[216];
  assign t[212] = t[244] ^ t[217];
  assign t[213] = t[75] ? x[108] : x[107];
  assign t[214] = t[75] ? x[110] : x[109];
  assign t[215] = t[210] ? x[112] : x[111];
  assign t[216] = t[75] ? x[114] : x[113];
  assign t[217] = t[210] ? x[116] : x[115];
  assign t[218] = t[245] ^ x[4];
  assign t[219] = t[246] ^ x[7];
  assign t[21] = ~(t[32] & t[223]);
  assign t[220] = t[247] ^ x[10];
  assign t[221] = t[248] ^ x[13];
  assign t[222] = t[249] ^ x[18];
  assign t[223] = t[250] ^ x[21];
  assign t[224] = t[251] ^ x[24];
  assign t[225] = t[252] ^ x[27];
  assign t[226] = t[253] ^ x[30];
  assign t[227] = t[254] ^ x[33];
  assign t[228] = t[255] ^ x[36];
  assign t[229] = t[256] ^ x[39];
  assign t[22] = ~(t[33] ^ t[34]);
  assign t[230] = t[257] ^ x[44];
  assign t[231] = t[258] ^ x[47];
  assign t[232] = t[259] ^ x[50];
  assign t[233] = t[260] ^ x[53];
  assign t[234] = t[261] ^ x[56];
  assign t[235] = t[262] ^ x[59];
  assign t[236] = t[263] ^ x[62];
  assign t[237] = t[264] ^ x[65];
  assign t[238] = t[265] ^ x[68];
  assign t[239] = t[266] ^ x[73];
  assign t[23] = t[35] ^ t[36];
  assign t[240] = t[267] ^ x[82];
  assign t[241] = t[268] ^ x[87];
  assign t[242] = t[269] ^ x[96];
  assign t[243] = t[270] ^ x[103];
  assign t[244] = t[271] ^ x[106];
  assign t[245] = (x[2] & x[3]);
  assign t[246] = (x[5] & x[6]);
  assign t[247] = (x[8] & x[9]);
  assign t[248] = (x[11] & x[12]);
  assign t[249] = (x[16] & x[17]);
  assign t[24] = t[37] ^ t[38];
  assign t[250] = (x[19] & x[20]);
  assign t[251] = (x[22] & x[23]);
  assign t[252] = (x[25] & x[26]);
  assign t[253] = (x[28] & x[29]);
  assign t[254] = (x[31] & x[32]);
  assign t[255] = (x[34] & x[35]);
  assign t[256] = (x[37] & x[38]);
  assign t[257] = (x[42] & x[43]);
  assign t[258] = (x[45] & x[46]);
  assign t[259] = (x[48] & x[49]);
  assign t[25] = ~(t[39] ^ t[40]);
  assign t[260] = (x[51] & x[52]);
  assign t[261] = (x[54] & x[55]);
  assign t[262] = (x[57] & x[58]);
  assign t[263] = (x[60] & x[61]);
  assign t[264] = (x[63] & x[64]);
  assign t[265] = (x[66] & x[67]);
  assign t[266] = (x[71] & x[72]);
  assign t[267] = (x[80] & x[81]);
  assign t[268] = (x[85] & x[86]);
  assign t[269] = (x[94] & x[95]);
  assign t[26] = t[41] ^ t[42];
  assign t[270] = (x[101] & x[102]);
  assign t[271] = (x[104] & x[105]);
  assign t[27] = ~(t[43] ^ t[24]);
  assign t[28] = t[44] ^ t[45];
  assign t[29] = ~(t[35] ^ t[46]);
  assign t[2] = ~(t[6] ^ t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = ~(t[49]);
  assign t[32] = ~(t[224]);
  assign t[33] = t[50] ^ t[17];
  assign t[34] = ~(t[51] ^ t[43]);
  assign t[35] = t[52] ^ t[53];
  assign t[36] = ~(t[54] ^ t[55]);
  assign t[37] = t[8] ? t[56] : t[225];
  assign t[38] = t[57] ^ t[58];
  assign t[39] = t[59] ^ t[60];
  assign t[3] = t[8] ? t[9] : t[218];
  assign t[40] = ~(t[41] ^ t[46]);
  assign t[41] = t[61] ^ t[62];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] ^ t[35]);
  assign t[44] = ~(t[66] ^ t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = t[70] ^ t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[226] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = ~(t[10] & t[11]);
  assign t[50] = t[76] ^ t[77];
  assign t[51] = t[78] ^ t[79];
  assign t[52] = t[80] ^ t[37];
  assign t[53] = t[57] ^ t[81];
  assign t[54] = t[82] ^ t[44];
  assign t[55] = ~(t[24] ^ t[83]);
  assign t[56] = t[225] ^ t[84];
  assign t[57] = t[85] ^ t[77];
  assign t[58] = t[86] & t[87];
  assign t[59] = t[24] ^ t[50];
  assign t[5] = ~(t[12] & t[13]);
  assign t[60] = ~(t[88] ^ t[89]);
  assign t[61] = t[90] ^ t[70];
  assign t[62] = t[91] & t[92];
  assign t[63] = t[93] ^ t[94];
  assign t[64] = t[95] ^ t[96];
  assign t[65] = ~(t[97] ^ t[98]);
  assign t[66] = t[99] ^ t[100];
  assign t[67] = ~(t[101] ^ t[102]);
  assign t[68] = t[103] ^ t[93];
  assign t[69] = t[104] & t[105];
  assign t[6] = ~(t[14] ^ t[15]);
  assign t[70] = t[8] ? t[106] : t[227];
  assign t[71] = t[107] ^ t[108];
  assign t[72] = ~(t[74] & t[109]);
  assign t[73] = ~(t[228] ^ t[110]);
  assign t[74] = ~(t[111] & t[112]);
  assign t[75] = ~(t[48]);
  assign t[76] = t[113] ^ t[37];
  assign t[77] = t[114] & t[115];
  assign t[78] = t[116] ^ t[70];
  assign t[79] = t[107] ^ t[117];
  assign t[7] = ~(t[16] ^ t[17]);
  assign t[80] = t[8] ? t[118] : t[229];
  assign t[81] = t[119] & t[120];
  assign t[82] = ~(t[121] ^ t[122]);
  assign t[83] = t[123] ^ t[108];
  assign t[84] = t[124] ? x[41] : x[40];
  assign t[85] = t[125] & t[126];
  assign t[86] = ~(t[127] ^ t[57]);
  assign t[87] = t[52] ^ t[115];
  assign t[88] = ~(t[45] ^ t[102]);
  assign t[89] = t[128] ^ t[129];
  assign t[8] = ~(t[18]);
  assign t[90] = t[8] ? t[130] : t[230];
  assign t[91] = ~(t[116]);
  assign t[92] = t[8] ? t[131] : t[231];
  assign t[93] = t[221] ^ t[132];
  assign t[94] = t[222] ^ t[133];
  assign t[95] = t[134] ^ t[135];
  assign t[96] = t[136] & t[137];
  assign t[97] = t[51] ^ t[138];
  assign t[98] = t[139] ^ t[140];
  assign t[99] = t[141] ^ t[142];
  assign t[9] = t[218] ^ t[19];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind81(x, y);
 input [116:0] x;
 output y;

 wire [262:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[143] ? x[56] : x[55];
  assign t[101] = ~(t[113] ^ t[55]);
  assign t[102] = t[35] ^ t[123];
  assign t[103] = t[31] ? x[58] : x[57];
  assign t[104] = t[144] & t[145];
  assign t[105] = t[146] & t[147];
  assign t[106] = ~(t[90] ^ t[70]);
  assign t[107] = t[148] ^ t[147];
  assign t[108] = ~(t[149] & t[150]);
  assign t[109] = t[151] ^ t[226];
  assign t[10] = ~(t[210]);
  assign t[110] = ~(t[221]);
  assign t[111] = t[152] & t[151];
  assign t[112] = t[153] ^ t[60];
  assign t[113] = t[154] ^ t[54];
  assign t[114] = t[118] ^ t[155];
  assign t[115] = t[61] ^ t[156];
  assign t[116] = t[30] ? t[157] : t[227];
  assign t[117] = t[158] ^ t[42];
  assign t[118] = t[80] ^ t[64];
  assign t[119] = t[143] ? x[66] : x[65];
  assign t[11] = ~(t[211]);
  assign t[120] = ~(t[126]);
  assign t[121] = ~(t[154]);
  assign t[122] = ~(t[54]);
  assign t[123] = t[8] ? t[159] : t[228];
  assign t[124] = t[35] ^ t[154];
  assign t[125] = t[154] ^ t[43];
  assign t[126] = t[123] ^ t[54];
  assign t[127] = ~(t[160] ^ t[161]);
  assign t[128] = t[162] ^ t[163];
  assign t[129] = t[8] ? t[164] : t[229];
  assign t[12] = ~(t[212]);
  assign t[130] = t[8] ? t[165] : t[230];
  assign t[131] = t[222] ^ t[166];
  assign t[132] = t[223] ^ t[167];
  assign t[133] = ~(t[138]);
  assign t[134] = ~(t[153]);
  assign t[135] = ~(t[59]);
  assign t[136] = t[168];
  assign t[137] = t[39] ^ t[153];
  assign t[138] = t[136] ^ t[59];
  assign t[139] = t[143] ? x[77] : x[76];
  assign t[13] = ~(t[20] | t[21]);
  assign t[140] = ~(t[18]);
  assign t[141] = t[224] ^ t[169];
  assign t[142] = t[225] ^ t[170];
  assign t[143] = ~(t[49]);
  assign t[144] = ~(t[171]);
  assign t[145] = ~(t[129]);
  assign t[146] = ~(t[130]);
  assign t[147] = t[8] ? t[172] : t[231];
  assign t[148] = t[130] ^ t[45];
  assign t[149] = ~(t[152] | t[151]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = ~(t[173] | t[110]);
  assign t[151] = ~(t[232]);
  assign t[152] = ~(t[226]);
  assign t[153] = ~t[174];
  assign t[154] = t[8] ? t[175] : t[233];
  assign t[155] = t[117] ^ t[176];
  assign t[156] = t[177] & t[178];
  assign t[157] = t[227] ^ t[179];
  assign t[158] = t[180] & t[181];
  assign t[159] = t[228] ^ t[182];
  assign t[15] = t[24] ^ t[25];
  assign t[160] = t[183] ^ t[184];
  assign t[161] = ~(t[185] ^ t[29]);
  assign t[162] = t[148] ^ t[186];
  assign t[163] = t[64] ^ t[187];
  assign t[164] = t[229] ^ t[188];
  assign t[165] = t[230] ^ t[189];
  assign t[166] = t[190] ? x[88] : x[87];
  assign t[167] = t[75] ? x[90] : x[89];
  assign t[168] = t[30] ? t[191] : t[234];
  assign t[169] = t[190] ? x[95] : x[94];
  assign t[16] = t[26] ^ t[27];
  assign t[170] = t[75] ? x[97] : x[96];
  assign t[171] = t[147] ^ t[130];
  assign t[172] = t[231] ^ t[192];
  assign t[173] = ~(t[218]);
  assign t[174] = t[30] ? t[193] : t[235];
  assign t[175] = t[233] ^ t[194];
  assign t[176] = t[195] & t[196];
  assign t[177] = ~(t[197] ^ t[61]);
  assign t[178] = t[39] ^ t[136];
  assign t[179] = t[143] ? x[102] : x[101];
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[180] = ~(t[198]);
  assign t[181] = ~(t[63]);
  assign t[182] = t[143] ? x[104] : x[103];
  assign t[183] = t[28] ^ t[199];
  assign t[184] = ~(t[200] ^ t[26]);
  assign t[185] = t[201] ^ t[105];
  assign t[186] = t[70] ^ t[202];
  assign t[187] = t[117] ^ t[53];
  assign t[188] = t[31] ? x[106] : x[105];
  assign t[189] = t[31] ? x[108] : x[107];
  assign t[18] = ~(t[30]);
  assign t[190] = ~(t[49]);
  assign t[191] = t[234] ^ t[203];
  assign t[192] = t[31] ? x[110] : x[109];
  assign t[193] = t[235] ^ t[204];
  assign t[194] = t[143] ? x[112] : x[111];
  assign t[195] = ~(t[158] ^ t[205]);
  assign t[196] = t[41] ^ t[198];
  assign t[197] = t[153] ^ t[59];
  assign t[198] = t[66] ^ t[80];
  assign t[199] = t[125] ^ t[85];
  assign t[19] = t[31] ? x[15] : x[14];
  assign t[1] = ~(t[4] | t[5]);
  assign t[200] = ~(t[34] ^ t[79]);
  assign t[201] = t[129] ^ t[45];
  assign t[202] = t[206] & t[207];
  assign t[203] = t[190] ? x[114] : x[113];
  assign t[204] = t[75] ? x[116] : x[115];
  assign t[205] = t[118] ^ t[63];
  assign t[206] = ~(t[104] ^ t[208]);
  assign t[207] = t[201] ^ t[171];
  assign t[208] = t[148] ^ t[129];
  assign t[209] = t[236] ^ x[4];
  assign t[20] = ~(t[213]);
  assign t[210] = t[237] ^ x[7];
  assign t[211] = t[238] ^ x[10];
  assign t[212] = t[239] ^ x[13];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[32] & t[214]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[61];
  assign t[227] = t[254] ^ x[64];
  assign t[228] = t[255] ^ x[69];
  assign t[229] = t[256] ^ x[72];
  assign t[22] = t[33] ^ t[34];
  assign t[230] = t[257] ^ x[75];
  assign t[231] = t[258] ^ x[80];
  assign t[232] = t[259] ^ x[83];
  assign t[233] = t[260] ^ x[86];
  assign t[234] = t[261] ^ x[93];
  assign t[235] = t[262] ^ x[100];
  assign t[236] = (x[2] & x[3]);
  assign t[237] = (x[5] & x[6]);
  assign t[238] = (x[8] & x[9]);
  assign t[239] = (x[11] & x[12]);
  assign t[23] = ~(t[24] ^ t[29]);
  assign t[240] = (x[16] & x[17]);
  assign t[241] = (x[19] & x[20]);
  assign t[242] = (x[22] & x[23]);
  assign t[243] = (x[25] & x[26]);
  assign t[244] = (x[28] & x[29]);
  assign t[245] = (x[31] & x[32]);
  assign t[246] = (x[34] & x[35]);
  assign t[247] = (x[37] & x[38]);
  assign t[248] = (x[40] & x[41]);
  assign t[249] = (x[43] & x[44]);
  assign t[24] = t[35] ^ t[36];
  assign t[250] = (x[46] & x[47]);
  assign t[251] = (x[49] & x[50]);
  assign t[252] = (x[52] & x[53]);
  assign t[253] = (x[59] & x[60]);
  assign t[254] = (x[62] & x[63]);
  assign t[255] = (x[67] & x[68]);
  assign t[256] = (x[70] & x[71]);
  assign t[257] = (x[73] & x[74]);
  assign t[258] = (x[78] & x[79]);
  assign t[259] = (x[81] & x[82]);
  assign t[25] = ~(t[37] ^ t[38]);
  assign t[260] = (x[84] & x[85]);
  assign t[261] = (x[91] & x[92]);
  assign t[262] = (x[98] & x[99]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = t[41] ^ t[42];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[6] ^ t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = ~(t[49]);
  assign t[32] = ~(t[215]);
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[34] = t[52] ^ t[53];
  assign t[35] = t[54] ^ t[43];
  assign t[36] = t[55] ^ t[56];
  assign t[37] = t[57] ^ t[33];
  assign t[38] = ~(t[28] ^ t[58]);
  assign t[39] = t[59] ^ t[60];
  assign t[3] = t[8] ? t[9] : t[209];
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[8] ? t[67] : t[216];
  assign t[44] = t[55] ^ t[68];
  assign t[45] = t[8] ? t[69] : t[217];
  assign t[46] = t[70] ^ t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[218] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = ~(t[10] & t[11]);
  assign t[50] = t[76] ^ t[77];
  assign t[51] = ~(t[78] ^ t[79]);
  assign t[52] = t[63] ^ t[80];
  assign t[53] = t[81] & t[82];
  assign t[54] = t[8] ? t[83] : t[219];
  assign t[55] = t[84] ^ t[85];
  assign t[56] = t[86] & t[87];
  assign t[57] = ~(t[88] ^ t[89]);
  assign t[58] = t[90] ^ t[71];
  assign t[59] = t[91];
  assign t[5] = ~(t[12] & t[13]);
  assign t[60] = t[92];
  assign t[61] = t[93] ^ t[94];
  assign t[62] = t[95] & t[96];
  assign t[63] = t[30] ? t[97] : t[220];
  assign t[64] = t[213] ^ t[98];
  assign t[65] = ~(t[80]);
  assign t[66] = t[215] ^ t[99];
  assign t[67] = t[216] ^ t[100];
  assign t[68] = t[101] & t[102];
  assign t[69] = t[217] ^ t[103];
  assign t[6] = ~(t[14] ^ t[15]);
  assign t[70] = t[104] ^ t[105];
  assign t[71] = t[106] & t[107];
  assign t[72] = ~(t[74] & t[108]);
  assign t[73] = ~(t[221] ^ t[109]);
  assign t[74] = ~(t[110] & t[111]);
  assign t[75] = ~(t[48]);
  assign t[76] = t[112] ^ t[94];
  assign t[77] = t[113] ^ t[68];
  assign t[78] = t[114] ^ t[58];
  assign t[79] = t[60] ^ t[115];
  assign t[7] = ~(t[16] ^ t[17]);
  assign t[80] = t[212] ^ t[116];
  assign t[81] = ~(t[52] ^ t[117]);
  assign t[82] = t[118] ^ t[66];
  assign t[83] = t[219] ^ t[119];
  assign t[84] = t[120] & t[121];
  assign t[85] = t[122] & t[123];
  assign t[86] = ~(t[84] ^ t[124]);
  assign t[87] = t[125] ^ t[126];
  assign t[88] = t[127] ^ t[27];
  assign t[89] = ~(t[128] ^ t[77]);
  assign t[8] = ~(t[18]);
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[30] ? t[131] : t[222];
  assign t[92] = t[30] ? t[132] : t[223];
  assign t[93] = t[133] & t[134];
  assign t[94] = t[135] & t[136];
  assign t[95] = ~(t[93] ^ t[137]);
  assign t[96] = t[112] ^ t[138];
  assign t[97] = t[220] ^ t[139];
  assign t[98] = t[140] ? t[141] : t[224];
  assign t[99] = t[30] ? t[142] : t[225];
  assign t[9] = t[209] ^ t[19];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind82(x, y);
 input [116:0] x;
 output y;

 wire [247:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[87]);
  assign t[101] = t[8] ? t[136] : t[211];
  assign t[102] = t[87] ^ t[26];
  assign t[103] = t[75] ? x[61] : x[60];
  assign t[104] = t[205] ^ t[137];
  assign t[105] = t[138] & t[139];
  assign t[106] = t[140] & t[71];
  assign t[107] = t[199] ^ t[141];
  assign t[108] = t[8] ? t[142] : t[212];
  assign t[109] = ~(t[143] & t[144]);
  assign t[10] = ~(t[195]);
  assign t[110] = t[145] ^ t[213];
  assign t[111] = ~(t[206]);
  assign t[112] = t[146] & t[145];
  assign t[113] = t[147] ^ t[64];
  assign t[114] = ~(t[148] ^ t[39]);
  assign t[115] = t[149] ^ t[150];
  assign t[116] = t[43] ^ t[107];
  assign t[117] = t[69] ^ t[29];
  assign t[118] = t[30] ? t[151] : t[214];
  assign t[119] = t[30] ? t[152] : t[215];
  assign t[11] = ~(t[196]);
  assign t[120] = t[153];
  assign t[121] = t[30] ? t[154] : t[216];
  assign t[122] = t[155] & t[156];
  assign t[123] = t[157] ^ t[53];
  assign t[124] = t[158] & t[159];
  assign t[125] = t[207] ^ t[160];
  assign t[126] = t[208] ^ t[161];
  assign t[127] = t[209] ^ t[162];
  assign t[128] = t[93] ? t[163] : t[217];
  assign t[129] = t[210] ^ t[164];
  assign t[12] = ~(t[197]);
  assign t[130] = t[165] & t[166];
  assign t[131] = t[167] ? x[81] : x[80];
  assign t[132] = t[168] & t[169];
  assign t[133] = ~(t[170] ^ t[95]);
  assign t[134] = t[149] ^ t[90];
  assign t[135] = t[101] ^ t[87];
  assign t[136] = t[211] ^ t[171];
  assign t[137] = t[31] ? x[83] : x[82];
  assign t[138] = ~(t[172]);
  assign t[139] = ~(t[43]);
  assign t[13] = ~(t[20] | t[21]);
  assign t[140] = ~(t[44]);
  assign t[141] = t[8] ? t[173] : t[218];
  assign t[142] = t[212] ^ t[174];
  assign t[143] = ~(t[146] | t[145]);
  assign t[144] = ~(t[175] | t[111]);
  assign t[145] = ~(t[219]);
  assign t[146] = ~(t[213]);
  assign t[147] = t[86] ^ t[26];
  assign t[148] = t[176] ^ t[124];
  assign t[149] = t[128] ^ t[60];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[95] ^ t[177];
  assign t[151] = t[214] ^ t[178];
  assign t[152] = t[215] ^ t[179];
  assign t[153] = t[30] ? t[180] : t[220];
  assign t[154] = t[216] ^ t[181];
  assign t[155] = ~(t[105] ^ t[182]);
  assign t[156] = t[116] ^ t[172];
  assign t[157] = t[183] & t[184];
  assign t[158] = ~(t[176] ^ t[123]);
  assign t[159] = t[91] ^ t[83];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = t[97] ? x[94] : x[93];
  assign t[161] = t[97] ? x[96] : x[95];
  assign t[162] = t[167] ? x[98] : x[97];
  assign t[163] = t[217] ^ t[185];
  assign t[164] = t[167] ? x[100] : x[99];
  assign t[165] = ~(t[157] ^ t[186]);
  assign t[166] = t[52] ^ t[187];
  assign t[167] = ~(t[49]);
  assign t[168] = ~(t[188]);
  assign t[169] = ~(t[88]);
  assign t[16] = t[26] ^ t[27];
  assign t[170] = t[88] ^ t[128];
  assign t[171] = t[97] ? x[102] : x[101];
  assign t[172] = t[71] ^ t[44];
  assign t[173] = t[218] ^ t[189];
  assign t[174] = t[31] ? x[104] : x[103];
  assign t[175] = ~(t[203]);
  assign t[176] = t[80] ^ t[120];
  assign t[177] = t[190] & t[191];
  assign t[178] = t[75] ? x[106] : x[105];
  assign t[179] = t[75] ? x[108] : x[107];
  assign t[17] = t[28] ^ t[29];
  assign t[180] = t[220] ^ t[192];
  assign t[181] = t[97] ? x[110] : x[109];
  assign t[182] = t[70] ^ t[43];
  assign t[183] = ~(t[187]);
  assign t[184] = ~(t[80]);
  assign t[185] = t[167] ? x[112] : x[111];
  assign t[186] = t[91] ^ t[80];
  assign t[187] = t[83] ^ t[120];
  assign t[188] = t[90] ^ t[128];
  assign t[189] = t[75] ? x[114] : x[113];
  assign t[18] = ~(t[30]);
  assign t[190] = ~(t[132] ^ t[193]);
  assign t[191] = t[57] ^ t[188];
  assign t[192] = t[31] ? x[116] : x[115];
  assign t[193] = t[149] ^ t[88];
  assign t[194] = t[221] ^ x[4];
  assign t[195] = t[222] ^ x[7];
  assign t[196] = t[223] ^ x[10];
  assign t[197] = t[224] ^ x[13];
  assign t[198] = t[225] ^ x[18];
  assign t[199] = t[226] ^ x[21];
  assign t[19] = t[31] ? x[15] : x[14];
  assign t[1] = ~(t[4] | t[5]);
  assign t[200] = t[227] ^ x[24];
  assign t[201] = t[228] ^ x[27];
  assign t[202] = t[229] ^ x[30];
  assign t[203] = t[230] ^ x[33];
  assign t[204] = t[231] ^ x[36];
  assign t[205] = t[232] ^ x[41];
  assign t[206] = t[233] ^ x[44];
  assign t[207] = t[234] ^ x[47];
  assign t[208] = t[235] ^ x[50];
  assign t[209] = t[236] ^ x[53];
  assign t[20] = ~(t[198]);
  assign t[210] = t[237] ^ x[56];
  assign t[211] = t[238] ^ x[59];
  assign t[212] = t[239] ^ x[64];
  assign t[213] = t[240] ^ x[67];
  assign t[214] = t[241] ^ x[70];
  assign t[215] = t[242] ^ x[73];
  assign t[216] = t[243] ^ x[76];
  assign t[217] = t[244] ^ x[79];
  assign t[218] = t[245] ^ x[86];
  assign t[219] = t[246] ^ x[89];
  assign t[21] = ~(t[32] & t[199]);
  assign t[220] = t[247] ^ x[92];
  assign t[221] = (x[2] & x[3]);
  assign t[222] = (x[5] & x[6]);
  assign t[223] = (x[8] & x[9]);
  assign t[224] = (x[11] & x[12]);
  assign t[225] = (x[16] & x[17]);
  assign t[226] = (x[19] & x[20]);
  assign t[227] = (x[22] & x[23]);
  assign t[228] = (x[25] & x[26]);
  assign t[229] = (x[28] & x[29]);
  assign t[22] = t[33] ^ t[34];
  assign t[230] = (x[31] & x[32]);
  assign t[231] = (x[34] & x[35]);
  assign t[232] = (x[39] & x[40]);
  assign t[233] = (x[42] & x[43]);
  assign t[234] = (x[45] & x[46]);
  assign t[235] = (x[48] & x[49]);
  assign t[236] = (x[51] & x[52]);
  assign t[237] = (x[54] & x[55]);
  assign t[238] = (x[57] & x[58]);
  assign t[239] = (x[62] & x[63]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (x[65] & x[66]);
  assign t[241] = (x[68] & x[69]);
  assign t[242] = (x[71] & x[72]);
  assign t[243] = (x[74] & x[75]);
  assign t[244] = (x[77] & x[78]);
  assign t[245] = (x[84] & x[85]);
  assign t[246] = (x[87] & x[88]);
  assign t[247] = (x[90] & x[91]);
  assign t[24] = t[37] ^ t[36];
  assign t[25] = ~(t[38] ^ t[39]);
  assign t[26] = t[8] ? t[40] : t[200];
  assign t[27] = t[41] ^ t[42];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[45] & t[46];
  assign t[2] = ~(t[6] ^ t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = ~(t[49]);
  assign t[32] = ~(t[201]);
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[34] = t[52] ^ t[53];
  assign t[35] = t[54] ^ t[55];
  assign t[36] = t[56] ^ t[42];
  assign t[37] = t[57] ^ t[58];
  assign t[38] = t[59] ^ t[17];
  assign t[39] = t[60] ^ t[61];
  assign t[3] = t[8] ? t[9] : t[194];
  assign t[40] = t[200] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[8] ? t[67] : t[202];
  assign t[44] = t[195] ^ t[68];
  assign t[45] = ~(t[28] ^ t[69]);
  assign t[46] = t[70] ^ t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[203] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = ~(t[10] & t[11]);
  assign t[50] = t[76] ^ t[77];
  assign t[51] = ~(t[78] ^ t[79]);
  assign t[52] = t[80] ^ t[81];
  assign t[53] = t[82] & t[83];
  assign t[54] = t[70] ^ t[84];
  assign t[55] = t[81] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ^ t[60];
  assign t[58] = t[89] & t[90];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = ~(t[12] & t[13]);
  assign t[60] = t[93] ? t[94] : t[204];
  assign t[61] = t[95] ^ t[96];
  assign t[62] = t[97] ? x[38] : x[37];
  assign t[63] = t[98] & t[99];
  assign t[64] = t[100] & t[101];
  assign t[65] = ~(t[56] ^ t[41]);
  assign t[66] = t[102] ^ t[101];
  assign t[67] = t[202] ^ t[103];
  assign t[68] = t[30] ? t[104] : t[205];
  assign t[69] = t[105] ^ t[106];
  assign t[6] = t[14] ^ t[15];
  assign t[70] = t[44] ^ t[107];
  assign t[71] = t[196] ^ t[108];
  assign t[72] = ~(t[74] & t[109]);
  assign t[73] = ~(t[206] ^ t[110]);
  assign t[74] = ~(t[111] & t[112]);
  assign t[75] = ~(t[48]);
  assign t[76] = t[16] ^ t[113];
  assign t[77] = ~(t[114] ^ t[115]);
  assign t[78] = t[116] ^ t[106];
  assign t[79] = t[107] ^ t[117];
  assign t[7] = ~(t[16] ^ t[17]);
  assign t[80] = ~t[118];
  assign t[81] = ~t[119];
  assign t[82] = ~(t[120]);
  assign t[83] = t[121];
  assign t[84] = t[69] ^ t[122];
  assign t[85] = t[123] ^ t[124];
  assign t[86] = t[8] ? t[125] : t[207];
  assign t[87] = t[8] ? t[126] : t[208];
  assign t[88] = t[93] ? t[127] : t[209];
  assign t[89] = ~(t[128]);
  assign t[8] = ~(t[18]);
  assign t[90] = t[93] ? t[129] : t[210];
  assign t[91] = t[120] ^ t[81];
  assign t[92] = t[123] ^ t[130];
  assign t[93] = ~(t[18]);
  assign t[94] = t[204] ^ t[131];
  assign t[95] = t[132] ^ t[58];
  assign t[96] = t[133] & t[134];
  assign t[97] = ~(t[49]);
  assign t[98] = ~(t[135]);
  assign t[99] = ~(t[86]);
  assign t[9] = t[194] ^ t[19];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind83(x, y);
 input [116:0] x;
 output y;

 wire [249:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[98] ^ t[134]);
  assign t[101] = t[135] ^ t[136];
  assign t[102] = t[207] ^ t[137];
  assign t[103] = t[138] & t[139];
  assign t[104] = t[140] & t[125];
  assign t[105] = t[141] & t[142];
  assign t[106] = t[7] ? t[143] : t[211];
  assign t[107] = t[197] ^ t[144];
  assign t[108] = ~(t[69] ^ t[145]);
  assign t[109] = t[146] ^ t[147];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[146] ^ t[148];
  assign t[111] = t[149] ^ t[62];
  assign t[112] = t[90] ^ t[40];
  assign t[113] = t[34] ^ t[150];
  assign t[114] = t[204] ^ t[151];
  assign t[115] = t[145] ^ t[70];
  assign t[116] = ~(t[152] & t[153]);
  assign t[117] = t[154] ^ t[212];
  assign t[118] = ~(t[208]);
  assign t[119] = t[155] & t[154];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = ~(t[49]);
  assign t[121] = t[7] ? t[156] : t[213];
  assign t[122] = t[210] ^ t[157];
  assign t[123] = t[26] ? t[158] : t[214];
  assign t[124] = t[26] ? t[159] : t[215];
  assign t[125] = t[160];
  assign t[126] = t[161] ? x[69] : x[68];
  assign t[127] = ~(t[111] ^ t[63]);
  assign t[128] = t[38] ^ t[133];
  assign t[129] = t[161] ? x[71] : x[70];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = ~(t[136]);
  assign t[131] = ~(t[149]);
  assign t[132] = ~(t[62]);
  assign t[133] = t[94] ? t[162] : t[216];
  assign t[134] = t[38] ^ t[149];
  assign t[135] = t[149] ^ t[60];
  assign t[136] = t[133] ^ t[62];
  assign t[137] = t[79] ? x[76] : x[75];
  assign t[138] = ~(t[163]);
  assign t[139] = ~(t[90]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[91]);
  assign t[141] = ~(t[103] ^ t[164]);
  assign t[142] = t[112] ^ t[163];
  assign t[143] = t[211] ^ t[165];
  assign t[144] = t[26] ? t[166] : t[217];
  assign t[145] = t[167] ^ t[168];
  assign t[146] = t[107] ^ t[114];
  assign t[147] = t[198] ^ t[169];
  assign t[148] = t[145] ^ t[170];
  assign t[149] = t[94] ? t[171] : t[218];
  assign t[14] = ~(t[26]);
  assign t[150] = t[172] & t[173];
  assign t[151] = t[7] ? t[174] : t[219];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[175] | t[118]);
  assign t[154] = ~(t[220]);
  assign t[155] = ~(t[212]);
  assign t[156] = t[213] ^ t[176];
  assign t[157] = t[120] ? x[90] : x[89];
  assign t[158] = t[214] ^ t[177];
  assign t[159] = t[215] ^ t[178];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[26] ? t[179] : t[221];
  assign t[161] = ~(t[49]);
  assign t[162] = t[216] ^ t[180];
  assign t[163] = t[125] ^ t[91];
  assign t[164] = t[67] ^ t[90];
  assign t[165] = t[79] ? x[95] : x[94];
  assign t[166] = t[217] ^ t[181];
  assign t[167] = t[182] & t[183];
  assign t[168] = t[184] & t[147];
  assign t[169] = t[7] ? t[185] : t[222];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[186] & t[187];
  assign t[171] = t[218] ^ t[188];
  assign t[172] = ~(t[189] ^ t[34]);
  assign t[173] = t[18] ^ t[86];
  assign t[174] = t[219] ^ t[190];
  assign t[175] = ~(t[202]);
  assign t[176] = t[120] ? x[100] : x[99];
  assign t[177] = t[79] ? x[102] : x[101];
  assign t[178] = t[27] ? x[104] : x[103];
  assign t[179] = t[221] ^ t[191];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[161] ? x[106] : x[105];
  assign t[181] = t[27] ? x[108] : x[107];
  assign t[182] = ~(t[192]);
  assign t[183] = ~(t[106]);
  assign t[184] = ~(t[107]);
  assign t[185] = t[222] ^ t[193];
  assign t[186] = ~(t[167] ^ t[194]);
  assign t[187] = t[195] ^ t[192];
  assign t[188] = t[161] ? x[110] : x[109];
  assign t[189] = t[121] ^ t[32];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[79] ? x[112] : x[111];
  assign t[191] = t[120] ? x[114] : x[113];
  assign t[192] = t[147] ^ t[107];
  assign t[193] = t[27] ? x[116] : x[115];
  assign t[194] = t[146] ^ t[106];
  assign t[195] = t[106] ^ t[114];
  assign t[196] = t[223] ^ x[4];
  assign t[197] = t[224] ^ x[9];
  assign t[198] = t[225] ^ x[12];
  assign t[199] = t[226] ^ x[15];
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[18];
  assign t[201] = t[228] ^ x[21];
  assign t[202] = t[229] ^ x[24];
  assign t[203] = t[230] ^ x[27];
  assign t[204] = t[231] ^ x[30];
  assign t[205] = t[232] ^ x[33];
  assign t[206] = t[233] ^ x[36];
  assign t[207] = t[234] ^ x[39];
  assign t[208] = t[235] ^ x[42];
  assign t[209] = t[236] ^ x[45];
  assign t[20] = ~(t[36] ^ t[37]);
  assign t[210] = t[237] ^ x[52];
  assign t[211] = t[238] ^ x[55];
  assign t[212] = t[239] ^ x[58];
  assign t[213] = t[240] ^ x[61];
  assign t[214] = t[241] ^ x[64];
  assign t[215] = t[242] ^ x[67];
  assign t[216] = t[243] ^ x[74];
  assign t[217] = t[244] ^ x[79];
  assign t[218] = t[245] ^ x[82];
  assign t[219] = t[246] ^ x[85];
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[247] ^ x[88];
  assign t[221] = t[248] ^ x[93];
  assign t[222] = t[249] ^ x[98];
  assign t[223] = (x[2] & x[3]);
  assign t[224] = (x[7] & x[8]);
  assign t[225] = (x[10] & x[11]);
  assign t[226] = (x[13] & x[14]);
  assign t[227] = (x[16] & x[17]);
  assign t[228] = (x[19] & x[20]);
  assign t[229] = (x[22] & x[23]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (x[25] & x[26]);
  assign t[231] = (x[28] & x[29]);
  assign t[232] = (x[31] & x[32]);
  assign t[233] = (x[34] & x[35]);
  assign t[234] = (x[37] & x[38]);
  assign t[235] = (x[40] & x[41]);
  assign t[236] = (x[43] & x[44]);
  assign t[237] = (x[50] & x[51]);
  assign t[238] = (x[53] & x[54]);
  assign t[239] = (x[56] & x[57]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (x[59] & x[60]);
  assign t[241] = (x[62] & x[63]);
  assign t[242] = (x[65] & x[66]);
  assign t[243] = (x[72] & x[73]);
  assign t[244] = (x[77] & x[78]);
  assign t[245] = (x[80] & x[81]);
  assign t[246] = (x[83] & x[84]);
  assign t[247] = (x[86] & x[87]);
  assign t[248] = (x[91] & x[92]);
  assign t[249] = (x[96] & x[97]);
  assign t[24] = ~(t[44] ^ t[10]);
  assign t[25] = ~(t[45] ^ t[46]);
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49]);
  assign t[28] = ~(t[197]);
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[199]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = t[7] ? t[52] : t[200];
  assign t[33] = t[7] ? t[53] : t[201];
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] & t[57];
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[62] ^ t[60];
  assign t[39] = t[63] ^ t[64];
  assign t[3] = t[7] ? t[8] : t[196];
  assign t[40] = ~t[65];
  assign t[41] = t[66] ^ t[59];
  assign t[42] = t[67] ^ t[68];
  assign t[43] = t[69] ^ t[70];
  assign t[44] = ~(t[71] ^ t[72]);
  assign t[45] = t[21] ^ t[73];
  assign t[46] = ~(t[74] ^ t[75]);
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = t[202] | t[78];
  assign t[49] = ~(t[79]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[203]);
  assign t[51] = ~(t[80] & t[204]);
  assign t[52] = t[200] ^ t[81];
  assign t[53] = t[201] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[85] & t[86];
  assign t[56] = ~(t[54] ^ t[87]);
  assign t[57] = t[88] ^ t[89];
  assign t[58] = t[90] ^ t[91];
  assign t[59] = t[92] & t[93];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[94] ? t[95] : t[205];
  assign t[61] = t[63] ^ t[96];
  assign t[62] = t[94] ? t[97] : t[206];
  assign t[63] = t[98] ^ t[99];
  assign t[64] = t[100] & t[101];
  assign t[65] = t[26] ? t[102] : t[207];
  assign t[66] = t[103] ^ t[104];
  assign t[67] = t[91] ^ t[40];
  assign t[68] = t[66] ^ t[105];
  assign t[69] = t[106] ^ t[107];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[108] & t[109];
  assign t[71] = t[110] ^ t[22];
  assign t[72] = t[111] ^ t[96];
  assign t[73] = t[112] ^ t[104];
  assign t[74] = t[33] ^ t[113];
  assign t[75] = t[114] ^ t[115];
  assign t[76] = ~(t[78] & t[116]);
  assign t[77] = ~(t[208] ^ t[117]);
  assign t[78] = ~(t[118] & t[119]);
  assign t[79] = ~(t[48]);
  assign t[7] = ~(t[14]);
  assign t[80] = ~(t[209]);
  assign t[81] = t[120] ? x[47] : x[46];
  assign t[82] = t[120] ? x[49] : x[48];
  assign t[83] = ~(t[89]);
  assign t[84] = ~(t[121]);
  assign t[85] = ~(t[32]);
  assign t[86] = t[7] ? t[122] : t[210];
  assign t[87] = t[18] ^ t[121];
  assign t[88] = t[121] ^ t[33];
  assign t[89] = t[86] ^ t[32];
  assign t[8] = t[196] ^ t[15];
  assign t[90] = ~t[123];
  assign t[91] = t[124];
  assign t[92] = ~(t[58] ^ t[66]);
  assign t[93] = t[67] ^ t[125];
  assign t[94] = ~(t[14]);
  assign t[95] = t[205] ^ t[126];
  assign t[96] = t[127] & t[128];
  assign t[97] = t[206] ^ t[129];
  assign t[98] = t[130] & t[131];
  assign t[99] = t[132] & t[133];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind84(x, y);
 input [116:0] x;
 output y;

 wire [260:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[137] ^ t[120];
  assign t[101] = t[138] & t[139];
  assign t[102] = t[217] ^ t[140];
  assign t[103] = t[141] ^ t[142];
  assign t[104] = t[41] ^ t[143];
  assign t[105] = t[144] ^ t[145];
  assign t[106] = ~t[146];
  assign t[107] = ~(t[71] ^ t[100]);
  assign t[108] = t[65] ^ t[147];
  assign t[109] = t[148] & t[149];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = ~(t[150] & t[151]);
  assign t[111] = t[152] ^ t[223];
  assign t[112] = ~(t[218]);
  assign t[113] = t[153] & t[152];
  assign t[114] = t[99] ^ t[154];
  assign t[115] = t[155] ^ t[156];
  assign t[116] = t[157] & t[158];
  assign t[117] = t[156] ^ t[144];
  assign t[118] = t[159] ^ t[160];
  assign t[119] = t[106] ^ t[99];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[161] & t[147];
  assign t[121] = t[162] ? x[56] : x[55];
  assign t[122] = t[162] ? x[58] : x[57];
  assign t[123] = t[163] & t[164];
  assign t[124] = t[165] & t[87];
  assign t[125] = t[220] ^ t[166];
  assign t[126] = t[221] ^ t[167];
  assign t[127] = ~(t[130]);
  assign t[128] = ~(t[95]);
  assign t[129] = t[36] ^ t[95];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[97] ^ t[58];
  assign t[131] = t[78] ? x[60] : x[59];
  assign t[132] = t[95] ^ t[58];
  assign t[133] = t[222] ^ t[168];
  assign t[134] = t[7] ? t[169] : t[224];
  assign t[135] = t[26] ? t[170] : t[225];
  assign t[136] = t[26] ? t[171] : t[226];
  assign t[137] = t[172] & t[173];
  assign t[138] = ~(t[137] ^ t[174]);
  assign t[139] = t[119] ^ t[175];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[162] ? x[71] : x[70];
  assign t[141] = t[155] ^ t[144];
  assign t[142] = t[176] & t[177];
  assign t[143] = t[132] ^ t[62];
  assign t[144] = t[178] ? t[179] : t[227];
  assign t[145] = t[159] ^ t[116];
  assign t[146] = t[26] ? t[180] : t[228];
  assign t[147] = t[181];
  assign t[148] = ~(t[123] ^ t[182]);
  assign t[149] = t[183] ^ t[184];
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[153] | t[152]);
  assign t[151] = ~(t[185] | t[112]);
  assign t[152] = ~(t[229]);
  assign t[153] = ~(t[223]);
  assign t[154] = t[100] ^ t[72];
  assign t[155] = t[178] ? t[186] : t[230];
  assign t[156] = t[178] ? t[187] : t[231];
  assign t[157] = ~(t[115] ^ t[159]);
  assign t[158] = t[117] ^ t[177];
  assign t[159] = t[188] ^ t[142];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[189] & t[190];
  assign t[161] = ~(t[98]);
  assign t[162] = ~(t[48]);
  assign t[163] = ~(t[184]);
  assign t[164] = ~(t[54]);
  assign t[165] = ~(t[55]);
  assign t[166] = t[162] ? x[88] : x[87];
  assign t[167] = t[27] ? x[90] : x[89];
  assign t[168] = t[78] ? x[92] : x[91];
  assign t[169] = t[224] ^ t[191];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[225] ^ t[192];
  assign t[171] = t[226] ^ t[193];
  assign t[172] = ~(t[175]);
  assign t[173] = ~(t[106]);
  assign t[174] = t[65] ^ t[106];
  assign t[175] = t[147] ^ t[98];
  assign t[176] = ~(t[156]);
  assign t[177] = t[178] ? t[194] : t[232];
  assign t[178] = ~(t[14]);
  assign t[179] = t[227] ^ t[195];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[228] ^ t[196];
  assign t[181] = t[26] ? t[197] : t[233];
  assign t[182] = t[73] ^ t[54];
  assign t[183] = t[54] ^ t[67];
  assign t[184] = t[87] ^ t[55];
  assign t[185] = ~(t[212]);
  assign t[186] = t[230] ^ t[198];
  assign t[187] = t[231] ^ t[199];
  assign t[188] = t[200] & t[201];
  assign t[189] = ~(t[188] ^ t[202]);
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[141] ^ t[203];
  assign t[191] = t[27] ? x[100] : x[99];
  assign t[192] = t[27] ? x[102] : x[101];
  assign t[193] = t[78] ? x[104] : x[103];
  assign t[194] = t[232] ^ t[204];
  assign t[195] = t[205] ? x[106] : x[105];
  assign t[196] = t[78] ? x[108] : x[107];
  assign t[197] = t[233] ^ t[206];
  assign t[198] = t[205] ? x[110] : x[109];
  assign t[199] = t[205] ? x[112] : x[111];
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = ~(t[203]);
  assign t[201] = ~(t[155]);
  assign t[202] = t[117] ^ t[155];
  assign t[203] = t[177] ^ t[156];
  assign t[204] = t[205] ? x[114] : x[113];
  assign t[205] = ~(t[48]);
  assign t[206] = t[162] ? x[116] : x[115];
  assign t[207] = t[234] ^ x[4];
  assign t[208] = t[235] ^ x[9];
  assign t[209] = t[236] ^ x[12];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[15];
  assign t[211] = t[238] ^ x[18];
  assign t[212] = t[239] ^ x[21];
  assign t[213] = t[240] ^ x[24];
  assign t[214] = t[241] ^ x[27];
  assign t[215] = t[242] ^ x[30];
  assign t[216] = t[243] ^ x[33];
  assign t[217] = t[244] ^ x[36];
  assign t[218] = t[245] ^ x[39];
  assign t[219] = t[246] ^ x[42];
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[247] ^ x[45];
  assign t[221] = t[248] ^ x[48];
  assign t[222] = t[249] ^ x[51];
  assign t[223] = t[250] ^ x[54];
  assign t[224] = t[251] ^ x[63];
  assign t[225] = t[252] ^ x[66];
  assign t[226] = t[253] ^ x[69];
  assign t[227] = t[254] ^ x[74];
  assign t[228] = t[255] ^ x[77];
  assign t[229] = t[256] ^ x[80];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[83];
  assign t[231] = t[258] ^ x[86];
  assign t[232] = t[259] ^ x[95];
  assign t[233] = t[260] ^ x[98];
  assign t[234] = (x[2] & x[3]);
  assign t[235] = (x[7] & x[8]);
  assign t[236] = (x[10] & x[11]);
  assign t[237] = (x[13] & x[14]);
  assign t[238] = (x[16] & x[17]);
  assign t[239] = (x[19] & x[20]);
  assign t[23] = ~(t[32] ^ t[42]);
  assign t[240] = (x[22] & x[23]);
  assign t[241] = (x[25] & x[26]);
  assign t[242] = (x[28] & x[29]);
  assign t[243] = (x[31] & x[32]);
  assign t[244] = (x[34] & x[35]);
  assign t[245] = (x[37] & x[38]);
  assign t[246] = (x[40] & x[41]);
  assign t[247] = (x[43] & x[44]);
  assign t[248] = (x[46] & x[47]);
  assign t[249] = (x[49] & x[50]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (x[52] & x[53]);
  assign t[251] = (x[61] & x[62]);
  assign t[252] = (x[64] & x[65]);
  assign t[253] = (x[67] & x[68]);
  assign t[254] = (x[72] & x[73]);
  assign t[255] = (x[75] & x[76]);
  assign t[256] = (x[78] & x[79]);
  assign t[257] = (x[81] & x[82]);
  assign t[258] = (x[84] & x[85]);
  assign t[259] = (x[93] & x[94]);
  assign t[25] = ~(t[45] ^ t[21]);
  assign t[260] = (x[96] & x[97]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[208]);
  assign t[29] = ~(t[209]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[210]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = ~(t[51] ^ t[45]);
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] & t[57];
  assign t[36] = t[58] ^ t[38];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[211] ^ t[61];
  assign t[39] = t[59] ^ t[62];
  assign t[3] = t[7] ? t[8] : t[207];
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] ^ t[68];
  assign t[43] = ~(t[69] ^ t[70]);
  assign t[44] = t[71] ^ t[72];
  assign t[45] = t[73] ^ t[74];
  assign t[46] = ~(t[75] & t[76]);
  assign t[47] = t[212] | t[77];
  assign t[48] = ~(t[78]);
  assign t[49] = ~(t[213]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[79] & t[211]);
  assign t[51] = ~(t[80] ^ t[81]);
  assign t[52] = t[82] ^ t[83];
  assign t[53] = ~(t[42] ^ t[21]);
  assign t[54] = t[7] ? t[84] : t[214];
  assign t[55] = t[7] ? t[85] : t[215];
  assign t[56] = ~(t[34] ^ t[86]);
  assign t[57] = t[73] ^ t[87];
  assign t[58] = t[208] ^ t[88];
  assign t[59] = t[89] ^ t[64];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[90] & t[91];
  assign t[61] = t[7] ? t[92] : t[216];
  assign t[62] = t[93] & t[94];
  assign t[63] = t[95] ^ t[38];
  assign t[64] = t[96] & t[97];
  assign t[65] = t[98] ^ t[99];
  assign t[66] = t[100] ^ t[101];
  assign t[67] = t[7] ? t[102] : t[217];
  assign t[68] = t[86] ^ t[35];
  assign t[69] = t[103] ^ t[19];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[104] ^ t[105]);
  assign t[71] = t[106] ^ t[98];
  assign t[72] = t[107] & t[108];
  assign t[73] = t[55] ^ t[67];
  assign t[74] = t[86] ^ t[109];
  assign t[75] = ~(t[77] & t[110]);
  assign t[76] = ~(t[218] ^ t[111]);
  assign t[77] = ~(t[112] & t[113]);
  assign t[78] = ~(t[47]);
  assign t[79] = ~(t[219]);
  assign t[7] = ~(t[14]);
  assign t[80] = t[20] ^ t[114];
  assign t[81] = t[115] ^ t[116];
  assign t[82] = t[117] ^ t[118];
  assign t[83] = t[119] ^ t[120];
  assign t[84] = t[214] ^ t[121];
  assign t[85] = t[215] ^ t[122];
  assign t[86] = t[123] ^ t[124];
  assign t[87] = t[7] ? t[125] : t[220];
  assign t[88] = t[26] ? t[126] : t[221];
  assign t[89] = t[127] & t[128];
  assign t[8] = t[207] ^ t[15];
  assign t[90] = ~(t[89] ^ t[129]);
  assign t[91] = t[63] ^ t[130];
  assign t[92] = t[216] ^ t[131];
  assign t[93] = ~(t[132] ^ t[59]);
  assign t[94] = t[36] ^ t[97];
  assign t[95] = t[7] ? t[133] : t[222];
  assign t[96] = ~(t[58]);
  assign t[97] = t[209] ^ t[134];
  assign t[98] = t[135];
  assign t[99] = ~t[136];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind85(x, y);
 input [116:0] x;
 output y;

 wire [242:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[124] ^ t[59];
  assign t[101] = t[134] ? t[135] : t[204];
  assign t[102] = t[134] ? t[136] : t[205];
  assign t[103] = ~(t[68] ^ t[137]);
  assign t[104] = t[138] ^ t[139];
  assign t[105] = t[140] & t[141];
  assign t[106] = ~(t[105] ^ t[142]);
  assign t[107] = t[18] ^ t[143];
  assign t[108] = ~(t[144] & t[145]);
  assign t[109] = t[146] ^ t[206];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = ~(t[202]);
  assign t[111] = t[147] & t[146];
  assign t[112] = ~(t[49]);
  assign t[113] = t[112] ? x[65] : x[64];
  assign t[114] = t[101] ^ t[120];
  assign t[115] = t[148] & t[139];
  assign t[116] = t[32] ^ t[54];
  assign t[117] = t[149] & t[150];
  assign t[118] = t[125] ^ t[151];
  assign t[119] = t[152] ^ t[89];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[134] ? t[153] : t[207];
  assign t[121] = t[137] ^ t[69];
  assign t[122] = t[26] ? t[154] : t[208];
  assign t[123] = t[26] ? t[155] : t[209];
  assign t[124] = t[156] ^ t[157];
  assign t[125] = t[86] ^ t[99];
  assign t[126] = t[158];
  assign t[127] = ~(t[152] ^ t[41]);
  assign t[128] = t[22] ^ t[95];
  assign t[129] = t[27] ? x[76] : x[75];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[75] ? x[78] : x[77];
  assign t[131] = t[7] ? t[159] : t[210];
  assign t[132] = t[7] ? t[160] : t[211];
  assign t[133] = t[26] ? t[161] : t[212];
  assign t[134] = ~(t[14]);
  assign t[135] = t[204] ^ t[162];
  assign t[136] = t[205] ^ t[163];
  assign t[137] = t[164] ^ t[115];
  assign t[138] = t[102] ^ t[120];
  assign t[139] = t[134] ? t[165] : t[213];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = ~(t[143]);
  assign t[141] = ~(t[32]);
  assign t[142] = t[45] ^ t[32];
  assign t[143] = t[35] ^ t[54];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[166] | t[110]);
  assign t[146] = ~(t[214]);
  assign t[147] = ~(t[206]);
  assign t[148] = ~(t[102]);
  assign t[149] = ~(t[116] ^ t[70]);
  assign t[14] = ~(t[26]);
  assign t[150] = t[45] ^ t[35];
  assign t[151] = t[124] ^ t[167];
  assign t[152] = t[131] ^ t[39];
  assign t[153] = t[207] ^ t[168];
  assign t[154] = t[208] ^ t[169];
  assign t[155] = t[209] ^ t[170];
  assign t[156] = t[171] & t[172];
  assign t[157] = t[173] & t[126];
  assign t[158] = t[26] ? t[174] : t[215];
  assign t[159] = t[210] ^ t[175];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[211] ^ t[176];
  assign t[161] = t[212] ^ t[177];
  assign t[162] = t[178] ? x[98] : x[97];
  assign t[163] = t[178] ? x[100] : x[99];
  assign t[164] = t[179] & t[180];
  assign t[165] = t[213] ^ t[181];
  assign t[166] = ~(t[197]);
  assign t[167] = t[182] & t[183];
  assign t[168] = t[178] ? x[102] : x[101];
  assign t[169] = t[75] ? x[104] : x[103];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[27] ? x[106] : x[105];
  assign t[171] = ~(t[184]);
  assign t[172] = ~(t[85]);
  assign t[173] = ~(t[86]);
  assign t[174] = t[215] ^ t[185];
  assign t[175] = t[75] ? x[108] : x[107];
  assign t[176] = t[27] ? x[110] : x[109];
  assign t[177] = t[75] ? x[112] : x[111];
  assign t[178] = ~(t[49]);
  assign t[179] = ~(t[186]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = ~(t[101]);
  assign t[181] = t[178] ? x[114] : x[113];
  assign t[182] = ~(t[156] ^ t[187]);
  assign t[183] = t[188] ^ t[184];
  assign t[184] = t[126] ^ t[86];
  assign t[185] = t[112] ? x[116] : x[115];
  assign t[186] = t[139] ^ t[102];
  assign t[187] = t[125] ^ t[85];
  assign t[188] = t[85] ^ t[99];
  assign t[189] = t[216] ^ x[4];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[217] ^ x[9];
  assign t[191] = t[218] ^ x[12];
  assign t[192] = t[219] ^ x[15];
  assign t[193] = t[220] ^ x[18];
  assign t[194] = t[221] ^ x[21];
  assign t[195] = t[222] ^ x[24];
  assign t[196] = t[223] ^ x[27];
  assign t[197] = t[224] ^ x[30];
  assign t[198] = t[225] ^ x[33];
  assign t[199] = t[226] ^ x[36];
  assign t[19] = t[34] & t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[39];
  assign t[201] = t[228] ^ x[42];
  assign t[202] = t[229] ^ x[45];
  assign t[203] = t[230] ^ x[48];
  assign t[204] = t[231] ^ x[57];
  assign t[205] = t[232] ^ x[60];
  assign t[206] = t[233] ^ x[63];
  assign t[207] = t[234] ^ x[68];
  assign t[208] = t[235] ^ x[71];
  assign t[209] = t[236] ^ x[74];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[81];
  assign t[211] = t[238] ^ x[84];
  assign t[212] = t[239] ^ x[87];
  assign t[213] = t[240] ^ x[90];
  assign t[214] = t[241] ^ x[93];
  assign t[215] = t[242] ^ x[96];
  assign t[216] = (x[2] & x[3]);
  assign t[217] = (x[7] & x[8]);
  assign t[218] = (x[10] & x[11]);
  assign t[219] = (x[13] & x[14]);
  assign t[21] = ~(t[25] ^ t[38]);
  assign t[220] = (x[16] & x[17]);
  assign t[221] = (x[19] & x[20]);
  assign t[222] = (x[22] & x[23]);
  assign t[223] = (x[25] & x[26]);
  assign t[224] = (x[28] & x[29]);
  assign t[225] = (x[31] & x[32]);
  assign t[226] = (x[34] & x[35]);
  assign t[227] = (x[37] & x[38]);
  assign t[228] = (x[40] & x[41]);
  assign t[229] = (x[43] & x[44]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (x[46] & x[47]);
  assign t[231] = (x[55] & x[56]);
  assign t[232] = (x[58] & x[59]);
  assign t[233] = (x[61] & x[62]);
  assign t[234] = (x[66] & x[67]);
  assign t[235] = (x[69] & x[70]);
  assign t[236] = (x[72] & x[73]);
  assign t[237] = (x[79] & x[80]);
  assign t[238] = (x[82] & x[83]);
  assign t[239] = (x[85] & x[86]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (x[88] & x[89]);
  assign t[241] = (x[91] & x[92]);
  assign t[242] = (x[94] & x[95]);
  assign t[24] = ~(t[43] ^ t[44]);
  assign t[25] = t[45] ^ t[46];
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49]);
  assign t[28] = ~(t[190]);
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[192]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = t[7] ? t[52] : t[193];
  assign t[33] = t[7] ? t[53] : t[194];
  assign t[34] = ~(t[54]);
  assign t[35] = t[7] ? t[55] : t[195];
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[37] = t[58] ^ t[59];
  assign t[38] = t[40] ^ t[60];
  assign t[39] = t[190] ^ t[61];
  assign t[3] = t[7] ? t[8] : t[189];
  assign t[40] = t[196] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[12] ^ t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[54] ^ t[33];
  assign t[46] = t[70] ^ t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[197] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[198]);
  assign t[51] = ~(t[76] & t[196]);
  assign t[52] = t[193] ^ t[77];
  assign t[53] = t[194] ^ t[78];
  assign t[54] = t[7] ? t[79] : t[199];
  assign t[55] = t[195] ^ t[80];
  assign t[56] = t[81] ^ t[82];
  assign t[57] = ~(t[83] ^ t[84]);
  assign t[58] = t[85] ^ t[86];
  assign t[59] = t[87] & t[88];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[41] ^ t[89];
  assign t[61] = t[26] ? t[90] : t[200];
  assign t[62] = t[7] ? t[91] : t[201];
  assign t[63] = t[92] & t[93];
  assign t[64] = t[94] & t[95];
  assign t[65] = ~(t[63] ^ t[96]);
  assign t[66] = t[97] ^ t[98];
  assign t[67] = t[99] ^ t[100];
  assign t[68] = t[101] ^ t[102];
  assign t[69] = t[103] & t[104];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[105] ^ t[19];
  assign t[71] = t[106] & t[107];
  assign t[72] = ~(t[74] & t[108]);
  assign t[73] = ~(t[202] ^ t[109]);
  assign t[74] = ~(t[110] & t[111]);
  assign t[75] = ~(t[48]);
  assign t[76] = ~(t[203]);
  assign t[77] = t[112] ? x[50] : x[49];
  assign t[78] = t[112] ? x[52] : x[51];
  assign t[79] = t[199] ^ t[113];
  assign t[7] = ~(t[14]);
  assign t[80] = t[112] ? x[54] : x[53];
  assign t[81] = t[114] ^ t[115];
  assign t[82] = t[116] ^ t[117];
  assign t[83] = t[118] ^ t[119];
  assign t[84] = t[120] ^ t[121];
  assign t[85] = ~t[122];
  assign t[86] = t[123];
  assign t[87] = ~(t[58] ^ t[124]);
  assign t[88] = t[125] ^ t[126];
  assign t[89] = t[127] & t[128];
  assign t[8] = t[189] ^ t[15];
  assign t[90] = t[200] ^ t[129];
  assign t[91] = t[201] ^ t[130];
  assign t[92] = ~(t[98]);
  assign t[93] = ~(t[131]);
  assign t[94] = ~(t[39]);
  assign t[95] = t[191] ^ t[132];
  assign t[96] = t[22] ^ t[131];
  assign t[97] = t[131] ^ t[40];
  assign t[98] = t[95] ^ t[39];
  assign t[99] = ~t[133];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind86(x, y);
 input [116:0] x;
 output y;

 wire [247:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[87]);
  assign t[101] = t[200] ^ t[137];
  assign t[102] = t[87] ^ t[26];
  assign t[103] = t[204] ^ t[138];
  assign t[104] = t[205] ^ t[139];
  assign t[105] = t[140] & t[141];
  assign t[106] = t[142] & t[71];
  assign t[107] = t[143];
  assign t[108] = t[8] ? t[144] : t[213];
  assign t[109] = ~(t[145] & t[146]);
  assign t[10] = ~(t[195]);
  assign t[110] = t[147] ^ t[214];
  assign t[111] = ~(t[206]);
  assign t[112] = t[148] & t[147];
  assign t[113] = t[149] ^ t[64];
  assign t[114] = ~(t[150] ^ t[39]);
  assign t[115] = t[151] ^ t[152];
  assign t[116] = t[43] ^ t[107];
  assign t[117] = t[69] ^ t[29];
  assign t[118] = t[207] ^ t[153];
  assign t[119] = t[208] ^ t[154];
  assign t[11] = ~(t[196]);
  assign t[120] = t[8] ? t[155] : t[215];
  assign t[121] = t[209] ^ t[156];
  assign t[122] = t[157] & t[158];
  assign t[123] = t[159] ^ t[53];
  assign t[124] = t[160] & t[161];
  assign t[125] = t[210] ^ t[162];
  assign t[126] = t[8] ? t[163] : t[216];
  assign t[127] = t[211] ^ t[164];
  assign t[128] = t[93] ? t[165] : t[217];
  assign t[129] = t[212] ^ t[166];
  assign t[12] = ~(t[197]);
  assign t[130] = t[167] & t[168];
  assign t[131] = t[169] ? x[79] : x[78];
  assign t[132] = t[170] & t[171];
  assign t[133] = ~(t[172] ^ t[95]);
  assign t[134] = t[151] ^ t[90];
  assign t[135] = ~(t[49]);
  assign t[136] = t[101] ^ t[87];
  assign t[137] = t[8] ? t[173] : t[218];
  assign t[138] = t[75] ? x[84] : x[83];
  assign t[139] = t[135] ? x[86] : x[85];
  assign t[13] = ~(t[20] | t[21]);
  assign t[140] = ~(t[174]);
  assign t[141] = ~(t[43]);
  assign t[142] = ~(t[44]);
  assign t[143] = t[8] ? t[175] : t[219];
  assign t[144] = t[213] ^ t[176];
  assign t[145] = ~(t[148] | t[147]);
  assign t[146] = ~(t[177] | t[111]);
  assign t[147] = ~(t[220]);
  assign t[148] = ~(t[214]);
  assign t[149] = t[86] ^ t[26];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[178] ^ t[124];
  assign t[151] = t[128] ^ t[60];
  assign t[152] = t[95] ^ t[179];
  assign t[153] = t[31] ? x[94] : x[93];
  assign t[154] = t[75] ? x[96] : x[95];
  assign t[155] = t[215] ^ t[180];
  assign t[156] = t[31] ? x[98] : x[97];
  assign t[157] = ~(t[105] ^ t[181]);
  assign t[158] = t[116] ^ t[174];
  assign t[159] = t[182] & t[183];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[178] ^ t[123]);
  assign t[161] = t[91] ^ t[83];
  assign t[162] = t[135] ? x[100] : x[99];
  assign t[163] = t[216] ^ t[184];
  assign t[164] = t[169] ? x[102] : x[101];
  assign t[165] = t[217] ^ t[185];
  assign t[166] = t[169] ? x[104] : x[103];
  assign t[167] = ~(t[159] ^ t[186]);
  assign t[168] = t[52] ^ t[187];
  assign t[169] = ~(t[49]);
  assign t[16] = t[26] ^ t[27];
  assign t[170] = ~(t[188]);
  assign t[171] = ~(t[88]);
  assign t[172] = t[88] ^ t[128];
  assign t[173] = t[218] ^ t[189];
  assign t[174] = t[71] ^ t[44];
  assign t[175] = t[219] ^ t[190];
  assign t[176] = t[75] ? x[106] : x[105];
  assign t[177] = ~(t[202]);
  assign t[178] = t[80] ^ t[120];
  assign t[179] = t[191] & t[192];
  assign t[17] = t[28] ^ t[29];
  assign t[180] = t[31] ? x[108] : x[107];
  assign t[181] = t[70] ^ t[43];
  assign t[182] = ~(t[187]);
  assign t[183] = ~(t[80]);
  assign t[184] = t[135] ? x[110] : x[109];
  assign t[185] = t[169] ? x[112] : x[111];
  assign t[186] = t[91] ^ t[80];
  assign t[187] = t[83] ^ t[120];
  assign t[188] = t[90] ^ t[128];
  assign t[189] = t[135] ? x[114] : x[113];
  assign t[18] = ~(t[30]);
  assign t[190] = t[75] ? x[116] : x[115];
  assign t[191] = ~(t[132] ^ t[193]);
  assign t[192] = t[57] ^ t[188];
  assign t[193] = t[151] ^ t[88];
  assign t[194] = t[221] ^ x[4];
  assign t[195] = t[222] ^ x[7];
  assign t[196] = t[223] ^ x[10];
  assign t[197] = t[224] ^ x[13];
  assign t[198] = t[225] ^ x[18];
  assign t[199] = t[226] ^ x[21];
  assign t[19] = t[31] ? x[15] : x[14];
  assign t[1] = ~(t[4] | t[5]);
  assign t[200] = t[227] ^ x[24];
  assign t[201] = t[228] ^ x[27];
  assign t[202] = t[229] ^ x[30];
  assign t[203] = t[230] ^ x[33];
  assign t[204] = t[231] ^ x[36];
  assign t[205] = t[232] ^ x[39];
  assign t[206] = t[233] ^ x[42];
  assign t[207] = t[234] ^ x[45];
  assign t[208] = t[235] ^ x[48];
  assign t[209] = t[236] ^ x[51];
  assign t[20] = ~(t[198]);
  assign t[210] = t[237] ^ x[54];
  assign t[211] = t[238] ^ x[57];
  assign t[212] = t[239] ^ x[60];
  assign t[213] = t[240] ^ x[65];
  assign t[214] = t[241] ^ x[68];
  assign t[215] = t[242] ^ x[71];
  assign t[216] = t[243] ^ x[74];
  assign t[217] = t[244] ^ x[77];
  assign t[218] = t[245] ^ x[82];
  assign t[219] = t[246] ^ x[89];
  assign t[21] = ~(t[32] & t[199]);
  assign t[220] = t[247] ^ x[92];
  assign t[221] = (x[2] & x[3]);
  assign t[222] = (x[5] & x[6]);
  assign t[223] = (x[8] & x[9]);
  assign t[224] = (x[11] & x[12]);
  assign t[225] = (x[16] & x[17]);
  assign t[226] = (x[19] & x[20]);
  assign t[227] = (x[22] & x[23]);
  assign t[228] = (x[25] & x[26]);
  assign t[229] = (x[28] & x[29]);
  assign t[22] = t[33] ^ t[34];
  assign t[230] = (x[31] & x[32]);
  assign t[231] = (x[34] & x[35]);
  assign t[232] = (x[37] & x[38]);
  assign t[233] = (x[40] & x[41]);
  assign t[234] = (x[43] & x[44]);
  assign t[235] = (x[46] & x[47]);
  assign t[236] = (x[49] & x[50]);
  assign t[237] = (x[52] & x[53]);
  assign t[238] = (x[55] & x[56]);
  assign t[239] = (x[58] & x[59]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (x[63] & x[64]);
  assign t[241] = (x[66] & x[67]);
  assign t[242] = (x[69] & x[70]);
  assign t[243] = (x[72] & x[73]);
  assign t[244] = (x[75] & x[76]);
  assign t[245] = (x[80] & x[81]);
  assign t[246] = (x[87] & x[88]);
  assign t[247] = (x[90] & x[91]);
  assign t[24] = t[37] ^ t[36];
  assign t[25] = ~(t[38] ^ t[39]);
  assign t[26] = t[198] ^ t[40];
  assign t[27] = t[41] ^ t[42];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[45] & t[46];
  assign t[2] = ~(t[6] ^ t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = ~(t[49]);
  assign t[32] = ~(t[200]);
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[34] = t[52] ^ t[53];
  assign t[35] = t[54] ^ t[55];
  assign t[36] = t[56] ^ t[42];
  assign t[37] = t[57] ^ t[58];
  assign t[38] = t[59] ^ t[17];
  assign t[39] = t[60] ^ t[61];
  assign t[3] = t[8] ? t[9] : t[194];
  assign t[40] = t[8] ? t[62] : t[201];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[67];
  assign t[44] = ~t[68];
  assign t[45] = ~(t[28] ^ t[69]);
  assign t[46] = t[70] ^ t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[202] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = ~(t[10] & t[11]);
  assign t[50] = t[76] ^ t[77];
  assign t[51] = ~(t[78] ^ t[79]);
  assign t[52] = t[80] ^ t[81];
  assign t[53] = t[82] & t[83];
  assign t[54] = t[70] ^ t[84];
  assign t[55] = t[81] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ^ t[60];
  assign t[58] = t[89] & t[90];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = ~(t[12] & t[13]);
  assign t[60] = t[93] ? t[94] : t[203];
  assign t[61] = t[95] ^ t[96];
  assign t[62] = t[201] ^ t[97];
  assign t[63] = t[98] & t[99];
  assign t[64] = t[100] & t[101];
  assign t[65] = ~(t[56] ^ t[41]);
  assign t[66] = t[102] ^ t[101];
  assign t[67] = t[8] ? t[103] : t[204];
  assign t[68] = t[8] ? t[104] : t[205];
  assign t[69] = t[105] ^ t[106];
  assign t[6] = t[14] ^ t[15];
  assign t[70] = t[44] ^ t[107];
  assign t[71] = t[108];
  assign t[72] = ~(t[74] & t[109]);
  assign t[73] = ~(t[206] ^ t[110]);
  assign t[74] = ~(t[111] & t[112]);
  assign t[75] = ~(t[48]);
  assign t[76] = t[16] ^ t[113];
  assign t[77] = ~(t[114] ^ t[115]);
  assign t[78] = t[116] ^ t[106];
  assign t[79] = t[107] ^ t[117];
  assign t[7] = ~(t[16] ^ t[17]);
  assign t[80] = t[8] ? t[118] : t[207];
  assign t[81] = t[8] ? t[119] : t[208];
  assign t[82] = ~(t[120]);
  assign t[83] = t[8] ? t[121] : t[209];
  assign t[84] = t[69] ^ t[122];
  assign t[85] = t[123] ^ t[124];
  assign t[86] = t[8] ? t[125] : t[210];
  assign t[87] = t[197] ^ t[126];
  assign t[88] = t[93] ? t[127] : t[211];
  assign t[89] = ~(t[128]);
  assign t[8] = ~(t[18]);
  assign t[90] = t[93] ? t[129] : t[212];
  assign t[91] = t[120] ^ t[81];
  assign t[92] = t[123] ^ t[130];
  assign t[93] = ~(t[18]);
  assign t[94] = t[203] ^ t[131];
  assign t[95] = t[132] ^ t[58];
  assign t[96] = t[133] & t[134];
  assign t[97] = t[135] ? x[62] : x[61];
  assign t[98] = ~(t[136]);
  assign t[99] = ~(t[86]);
  assign t[9] = t[194] ^ t[19];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind87(x, y);
 input [116:0] x;
 output y;

 wire [249:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[98] ^ t[135]);
  assign t[101] = t[136] ^ t[137];
  assign t[102] = t[79] ? x[53] : x[52];
  assign t[103] = t[138] & t[139];
  assign t[104] = t[140] & t[126];
  assign t[105] = t[141] & t[142];
  assign t[106] = t[143];
  assign t[107] = ~t[144];
  assign t[108] = ~(t[69] ^ t[145]);
  assign t[109] = t[146] ^ t[147];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[146] ^ t[148];
  assign t[111] = t[149] ^ t[62];
  assign t[112] = t[90] ^ t[40];
  assign t[113] = t[34] ^ t[150];
  assign t[114] = t[151];
  assign t[115] = t[145] ^ t[70];
  assign t[116] = ~(t[152] & t[153]);
  assign t[117] = t[154] ^ t[212];
  assign t[118] = ~(t[208]);
  assign t[119] = t[155] & t[154];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[156] ? x[58] : x[57];
  assign t[121] = t[156] ? x[60] : x[59];
  assign t[122] = t[7] ? t[157] : t[213];
  assign t[123] = t[7] ? t[158] : t[214];
  assign t[124] = t[210] ^ t[159];
  assign t[125] = t[211] ^ t[160];
  assign t[126] = t[7] ? t[161] : t[215];
  assign t[127] = t[162] ? x[71] : x[70];
  assign t[128] = ~(t[111] ^ t[63]);
  assign t[129] = t[38] ^ t[134];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[162] ? x[73] : x[72];
  assign t[131] = ~(t[137]);
  assign t[132] = ~(t[149]);
  assign t[133] = ~(t[62]);
  assign t[134] = t[94] ? t[163] : t[216];
  assign t[135] = t[38] ^ t[149];
  assign t[136] = t[149] ^ t[60];
  assign t[137] = t[134] ^ t[62];
  assign t[138] = ~(t[164]);
  assign t[139] = ~(t[90]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[91]);
  assign t[141] = ~(t[103] ^ t[165]);
  assign t[142] = t[112] ^ t[164];
  assign t[143] = t[7] ? t[166] : t[217];
  assign t[144] = t[7] ? t[167] : t[218];
  assign t[145] = t[168] ^ t[169];
  assign t[146] = t[107] ^ t[114];
  assign t[147] = t[170];
  assign t[148] = t[145] ^ t[171];
  assign t[149] = t[94] ? t[172] : t[219];
  assign t[14] = ~(t[26]);
  assign t[150] = t[173] & t[174];
  assign t[151] = t[7] ? t[175] : t[220];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[176] | t[118]);
  assign t[154] = ~(t[221]);
  assign t[155] = ~(t[212]);
  assign t[156] = ~(t[49]);
  assign t[157] = t[213] ^ t[177];
  assign t[158] = t[214] ^ t[178];
  assign t[159] = t[27] ? x[93] : x[92];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[27] ? x[95] : x[94];
  assign t[161] = t[215] ^ t[179];
  assign t[162] = ~(t[49]);
  assign t[163] = t[216] ^ t[180];
  assign t[164] = t[126] ^ t[91];
  assign t[165] = t[67] ^ t[90];
  assign t[166] = t[217] ^ t[181];
  assign t[167] = t[218] ^ t[182];
  assign t[168] = t[183] & t[184];
  assign t[169] = t[185] & t[147];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[7] ? t[186] : t[222];
  assign t[171] = t[187] & t[188];
  assign t[172] = t[219] ^ t[189];
  assign t[173] = ~(t[190] ^ t[34]);
  assign t[174] = t[18] ^ t[86];
  assign t[175] = t[220] ^ t[191];
  assign t[176] = ~(t[202]);
  assign t[177] = t[156] ? x[100] : x[99];
  assign t[178] = t[156] ? x[102] : x[101];
  assign t[179] = t[27] ? x[104] : x[103];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[162] ? x[106] : x[105];
  assign t[181] = t[79] ? x[108] : x[107];
  assign t[182] = t[156] ? x[110] : x[109];
  assign t[183] = ~(t[192]);
  assign t[184] = ~(t[106]);
  assign t[185] = ~(t[107]);
  assign t[186] = t[222] ^ t[193];
  assign t[187] = ~(t[168] ^ t[194]);
  assign t[188] = t[195] ^ t[192];
  assign t[189] = t[162] ? x[112] : x[111];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[122] ^ t[32];
  assign t[191] = t[79] ? x[114] : x[113];
  assign t[192] = t[147] ^ t[107];
  assign t[193] = t[79] ? x[116] : x[115];
  assign t[194] = t[146] ^ t[106];
  assign t[195] = t[106] ^ t[114];
  assign t[196] = t[223] ^ x[4];
  assign t[197] = t[224] ^ x[9];
  assign t[198] = t[225] ^ x[12];
  assign t[199] = t[226] ^ x[15];
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[18];
  assign t[201] = t[228] ^ x[21];
  assign t[202] = t[229] ^ x[24];
  assign t[203] = t[230] ^ x[27];
  assign t[204] = t[231] ^ x[30];
  assign t[205] = t[232] ^ x[33];
  assign t[206] = t[233] ^ x[36];
  assign t[207] = t[234] ^ x[39];
  assign t[208] = t[235] ^ x[42];
  assign t[209] = t[236] ^ x[45];
  assign t[20] = ~(t[36] ^ t[37]);
  assign t[210] = t[237] ^ x[48];
  assign t[211] = t[238] ^ x[51];
  assign t[212] = t[239] ^ x[56];
  assign t[213] = t[240] ^ x[63];
  assign t[214] = t[241] ^ x[66];
  assign t[215] = t[242] ^ x[69];
  assign t[216] = t[243] ^ x[76];
  assign t[217] = t[244] ^ x[79];
  assign t[218] = t[245] ^ x[82];
  assign t[219] = t[246] ^ x[85];
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[247] ^ x[88];
  assign t[221] = t[248] ^ x[91];
  assign t[222] = t[249] ^ x[98];
  assign t[223] = (x[2] & x[3]);
  assign t[224] = (x[7] & x[8]);
  assign t[225] = (x[10] & x[11]);
  assign t[226] = (x[13] & x[14]);
  assign t[227] = (x[16] & x[17]);
  assign t[228] = (x[19] & x[20]);
  assign t[229] = (x[22] & x[23]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (x[25] & x[26]);
  assign t[231] = (x[28] & x[29]);
  assign t[232] = (x[31] & x[32]);
  assign t[233] = (x[34] & x[35]);
  assign t[234] = (x[37] & x[38]);
  assign t[235] = (x[40] & x[41]);
  assign t[236] = (x[43] & x[44]);
  assign t[237] = (x[46] & x[47]);
  assign t[238] = (x[49] & x[50]);
  assign t[239] = (x[54] & x[55]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (x[61] & x[62]);
  assign t[241] = (x[64] & x[65]);
  assign t[242] = (x[67] & x[68]);
  assign t[243] = (x[74] & x[75]);
  assign t[244] = (x[77] & x[78]);
  assign t[245] = (x[80] & x[81]);
  assign t[246] = (x[83] & x[84]);
  assign t[247] = (x[86] & x[87]);
  assign t[248] = (x[89] & x[90]);
  assign t[249] = (x[96] & x[97]);
  assign t[24] = ~(t[44] ^ t[10]);
  assign t[25] = ~(t[45] ^ t[46]);
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49]);
  assign t[28] = ~(t[197]);
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[199]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = t[199] ^ t[52];
  assign t[33] = t[200] ^ t[53];
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] & t[57];
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[62] ^ t[60];
  assign t[39] = t[63] ^ t[64];
  assign t[3] = t[7] ? t[8] : t[196];
  assign t[40] = t[7] ? t[65] : t[201];
  assign t[41] = t[66] ^ t[59];
  assign t[42] = t[67] ^ t[68];
  assign t[43] = t[69] ^ t[70];
  assign t[44] = ~(t[71] ^ t[72]);
  assign t[45] = t[21] ^ t[73];
  assign t[46] = ~(t[74] ^ t[75]);
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = t[202] | t[78];
  assign t[49] = ~(t[79]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[200]);
  assign t[51] = ~(t[80] & t[203]);
  assign t[52] = t[7] ? t[81] : t[204];
  assign t[53] = t[7] ? t[82] : t[205];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[85] & t[86];
  assign t[56] = ~(t[54] ^ t[87]);
  assign t[57] = t[88] ^ t[89];
  assign t[58] = t[90] ^ t[91];
  assign t[59] = t[92] & t[93];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[94] ? t[95] : t[206];
  assign t[61] = t[63] ^ t[96];
  assign t[62] = t[94] ? t[97] : t[207];
  assign t[63] = t[98] ^ t[99];
  assign t[64] = t[100] & t[101];
  assign t[65] = t[201] ^ t[102];
  assign t[66] = t[103] ^ t[104];
  assign t[67] = t[91] ^ t[40];
  assign t[68] = t[66] ^ t[105];
  assign t[69] = t[106] ^ t[107];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[108] & t[109];
  assign t[71] = t[110] ^ t[22];
  assign t[72] = t[111] ^ t[96];
  assign t[73] = t[112] ^ t[104];
  assign t[74] = t[33] ^ t[113];
  assign t[75] = t[114] ^ t[115];
  assign t[76] = ~(t[78] & t[116]);
  assign t[77] = ~(t[208] ^ t[117]);
  assign t[78] = ~(t[118] & t[119]);
  assign t[79] = ~(t[48]);
  assign t[7] = ~(t[14]);
  assign t[80] = ~(t[209]);
  assign t[81] = t[204] ^ t[120];
  assign t[82] = t[205] ^ t[121];
  assign t[83] = ~(t[89]);
  assign t[84] = ~(t[122]);
  assign t[85] = ~(t[32]);
  assign t[86] = t[209] ^ t[123];
  assign t[87] = t[18] ^ t[122];
  assign t[88] = t[122] ^ t[33];
  assign t[89] = t[86] ^ t[32];
  assign t[8] = t[196] ^ t[15];
  assign t[90] = t[7] ? t[124] : t[210];
  assign t[91] = t[7] ? t[125] : t[211];
  assign t[92] = ~(t[58] ^ t[66]);
  assign t[93] = t[67] ^ t[126];
  assign t[94] = ~(t[14]);
  assign t[95] = t[206] ^ t[127];
  assign t[96] = t[128] & t[129];
  assign t[97] = t[207] ^ t[130];
  assign t[98] = t[131] & t[132];
  assign t[99] = t[133] & t[134];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind88(x, y);
 input [116:0] x;
 output y;

 wire [260:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[137] ^ t[120];
  assign t[101] = t[138] & t[139];
  assign t[102] = t[7] ? t[140] : t[222];
  assign t[103] = t[141] ^ t[142];
  assign t[104] = t[41] ^ t[143];
  assign t[105] = t[144] ^ t[145];
  assign t[106] = t[7] ? t[146] : t[223];
  assign t[107] = ~(t[71] ^ t[100]);
  assign t[108] = t[65] ^ t[147];
  assign t[109] = t[148] & t[149];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = ~(t[150] & t[151]);
  assign t[111] = t[152] ^ t[224];
  assign t[112] = ~(t[216]);
  assign t[113] = t[153] & t[152];
  assign t[114] = t[99] ^ t[154];
  assign t[115] = t[155] ^ t[156];
  assign t[116] = t[157] & t[158];
  assign t[117] = t[156] ^ t[144];
  assign t[118] = t[159] ^ t[160];
  assign t[119] = t[106] ^ t[99];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[161] & t[147];
  assign t[121] = t[162] ? x[59] : x[58];
  assign t[122] = t[218] ^ t[163];
  assign t[123] = t[164] & t[165];
  assign t[124] = t[166] & t[87];
  assign t[125] = t[7] ? t[167] : t[225];
  assign t[126] = t[219] ^ t[168];
  assign t[127] = ~(t[130]);
  assign t[128] = ~(t[95]);
  assign t[129] = t[36] ^ t[95];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[97] ^ t[58];
  assign t[131] = t[78] ? x[64] : x[63];
  assign t[132] = t[95] ^ t[58];
  assign t[133] = t[7] ? t[169] : t[226];
  assign t[134] = t[7] ? t[170] : t[227];
  assign t[135] = t[220] ^ t[171];
  assign t[136] = t[221] ^ t[172];
  assign t[137] = t[173] & t[174];
  assign t[138] = ~(t[137] ^ t[175]);
  assign t[139] = t[119] ^ t[176];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[222] ^ t[177];
  assign t[141] = t[155] ^ t[144];
  assign t[142] = t[178] & t[179];
  assign t[143] = t[132] ^ t[62];
  assign t[144] = t[180] ? t[181] : t[228];
  assign t[145] = t[159] ^ t[116];
  assign t[146] = t[223] ^ t[182];
  assign t[147] = t[7] ? t[183] : t[229];
  assign t[148] = ~(t[123] ^ t[184]);
  assign t[149] = t[185] ^ t[186];
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[153] | t[152]);
  assign t[151] = ~(t[187] | t[112]);
  assign t[152] = ~(t[230]);
  assign t[153] = ~(t[224]);
  assign t[154] = t[100] ^ t[72];
  assign t[155] = t[180] ? t[188] : t[231];
  assign t[156] = t[180] ? t[189] : t[232];
  assign t[157] = ~(t[115] ^ t[159]);
  assign t[158] = t[117] ^ t[179];
  assign t[159] = t[190] ^ t[142];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[191] & t[192];
  assign t[161] = ~(t[98]);
  assign t[162] = ~(t[48]);
  assign t[163] = t[162] ? x[87] : x[86];
  assign t[164] = ~(t[186]);
  assign t[165] = ~(t[54]);
  assign t[166] = ~(t[55]);
  assign t[167] = t[225] ^ t[193];
  assign t[168] = t[162] ? x[89] : x[88];
  assign t[169] = t[226] ^ t[194];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[227] ^ t[195];
  assign t[171] = t[27] ? x[91] : x[90];
  assign t[172] = t[78] ? x[93] : x[92];
  assign t[173] = ~(t[176]);
  assign t[174] = ~(t[106]);
  assign t[175] = t[65] ^ t[106];
  assign t[176] = t[147] ^ t[98];
  assign t[177] = t[162] ? x[95] : x[94];
  assign t[178] = ~(t[156]);
  assign t[179] = t[180] ? t[196] : t[233];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = ~(t[14]);
  assign t[181] = t[228] ^ t[197];
  assign t[182] = t[27] ? x[100] : x[99];
  assign t[183] = t[229] ^ t[198];
  assign t[184] = t[73] ^ t[54];
  assign t[185] = t[54] ^ t[67];
  assign t[186] = t[87] ^ t[55];
  assign t[187] = ~(t[211]);
  assign t[188] = t[231] ^ t[199];
  assign t[189] = t[232] ^ t[200];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[201] & t[202];
  assign t[191] = ~(t[190] ^ t[203]);
  assign t[192] = t[141] ^ t[204];
  assign t[193] = t[162] ? x[102] : x[101];
  assign t[194] = t[78] ? x[104] : x[103];
  assign t[195] = t[78] ? x[106] : x[105];
  assign t[196] = t[233] ^ t[205];
  assign t[197] = t[206] ? x[108] : x[107];
  assign t[198] = t[27] ? x[110] : x[109];
  assign t[199] = t[206] ? x[112] : x[111];
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[206] ? x[114] : x[113];
  assign t[201] = ~(t[204]);
  assign t[202] = ~(t[155]);
  assign t[203] = t[117] ^ t[155];
  assign t[204] = t[179] ^ t[156];
  assign t[205] = t[206] ? x[116] : x[115];
  assign t[206] = ~(t[48]);
  assign t[207] = t[234] ^ x[4];
  assign t[208] = t[235] ^ x[9];
  assign t[209] = t[236] ^ x[12];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[15];
  assign t[211] = t[238] ^ x[18];
  assign t[212] = t[239] ^ x[21];
  assign t[213] = t[240] ^ x[24];
  assign t[214] = t[241] ^ x[27];
  assign t[215] = t[242] ^ x[30];
  assign t[216] = t[243] ^ x[33];
  assign t[217] = t[244] ^ x[36];
  assign t[218] = t[245] ^ x[39];
  assign t[219] = t[246] ^ x[42];
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[247] ^ x[45];
  assign t[221] = t[248] ^ x[48];
  assign t[222] = t[249] ^ x[51];
  assign t[223] = t[250] ^ x[54];
  assign t[224] = t[251] ^ x[57];
  assign t[225] = t[252] ^ x[62];
  assign t[226] = t[253] ^ x[67];
  assign t[227] = t[254] ^ x[70];
  assign t[228] = t[255] ^ x[73];
  assign t[229] = t[256] ^ x[76];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[79];
  assign t[231] = t[258] ^ x[82];
  assign t[232] = t[259] ^ x[85];
  assign t[233] = t[260] ^ x[98];
  assign t[234] = (x[2] & x[3]);
  assign t[235] = (x[7] & x[8]);
  assign t[236] = (x[10] & x[11]);
  assign t[237] = (x[13] & x[14]);
  assign t[238] = (x[16] & x[17]);
  assign t[239] = (x[19] & x[20]);
  assign t[23] = ~(t[32] ^ t[42]);
  assign t[240] = (x[22] & x[23]);
  assign t[241] = (x[25] & x[26]);
  assign t[242] = (x[28] & x[29]);
  assign t[243] = (x[31] & x[32]);
  assign t[244] = (x[34] & x[35]);
  assign t[245] = (x[37] & x[38]);
  assign t[246] = (x[40] & x[41]);
  assign t[247] = (x[43] & x[44]);
  assign t[248] = (x[46] & x[47]);
  assign t[249] = (x[49] & x[50]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (x[52] & x[53]);
  assign t[251] = (x[55] & x[56]);
  assign t[252] = (x[60] & x[61]);
  assign t[253] = (x[65] & x[66]);
  assign t[254] = (x[68] & x[69]);
  assign t[255] = (x[71] & x[72]);
  assign t[256] = (x[74] & x[75]);
  assign t[257] = (x[77] & x[78]);
  assign t[258] = (x[80] & x[81]);
  assign t[259] = (x[83] & x[84]);
  assign t[25] = ~(t[45] ^ t[21]);
  assign t[260] = (x[96] & x[97]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[208]);
  assign t[29] = ~(t[209]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[210]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = ~(t[51] ^ t[45]);
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] & t[57];
  assign t[36] = t[58] ^ t[38];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[61];
  assign t[39] = t[59] ^ t[62];
  assign t[3] = t[7] ? t[8] : t[207];
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] ^ t[68];
  assign t[43] = ~(t[69] ^ t[70]);
  assign t[44] = t[71] ^ t[72];
  assign t[45] = t[73] ^ t[74];
  assign t[46] = ~(t[75] & t[76]);
  assign t[47] = t[211] | t[77];
  assign t[48] = ~(t[78]);
  assign t[49] = ~(t[212]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[79] & t[213]);
  assign t[51] = ~(t[80] ^ t[81]);
  assign t[52] = t[82] ^ t[83];
  assign t[53] = ~(t[42] ^ t[21]);
  assign t[54] = t[7] ? t[84] : t[214];
  assign t[55] = t[210] ^ t[85];
  assign t[56] = ~(t[34] ^ t[86]);
  assign t[57] = t[73] ^ t[87];
  assign t[58] = ~t[88];
  assign t[59] = t[89] ^ t[64];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[90] & t[91];
  assign t[61] = t[7] ? t[92] : t[215];
  assign t[62] = t[93] & t[94];
  assign t[63] = t[95] ^ t[38];
  assign t[64] = t[96] & t[97];
  assign t[65] = t[98] ^ t[99];
  assign t[66] = t[100] ^ t[101];
  assign t[67] = t[212] ^ t[102];
  assign t[68] = t[86] ^ t[35];
  assign t[69] = t[103] ^ t[19];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[104] ^ t[105]);
  assign t[71] = t[106] ^ t[98];
  assign t[72] = t[107] & t[108];
  assign t[73] = t[55] ^ t[67];
  assign t[74] = t[86] ^ t[109];
  assign t[75] = ~(t[77] & t[110]);
  assign t[76] = ~(t[216] ^ t[111]);
  assign t[77] = ~(t[112] & t[113]);
  assign t[78] = ~(t[47]);
  assign t[79] = ~(t[217]);
  assign t[7] = ~(t[14]);
  assign t[80] = t[20] ^ t[114];
  assign t[81] = t[115] ^ t[116];
  assign t[82] = t[117] ^ t[118];
  assign t[83] = t[119] ^ t[120];
  assign t[84] = t[214] ^ t[121];
  assign t[85] = t[7] ? t[122] : t[218];
  assign t[86] = t[123] ^ t[124];
  assign t[87] = t[217] ^ t[125];
  assign t[88] = t[7] ? t[126] : t[219];
  assign t[89] = t[127] & t[128];
  assign t[8] = t[207] ^ t[15];
  assign t[90] = ~(t[89] ^ t[129]);
  assign t[91] = t[63] ^ t[130];
  assign t[92] = t[215] ^ t[131];
  assign t[93] = ~(t[132] ^ t[59]);
  assign t[94] = t[36] ^ t[97];
  assign t[95] = t[133];
  assign t[96] = ~(t[58]);
  assign t[97] = t[134];
  assign t[98] = t[7] ? t[135] : t[220];
  assign t[99] = t[7] ? t[136] : t[221];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind89(x, y);
 input [116:0] x;
 output y;

 wire [242:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[126] ^ t[59];
  assign t[101] = t[136] ? t[137] : t[207];
  assign t[102] = t[136] ? t[138] : t[208];
  assign t[103] = ~(t[68] ^ t[139]);
  assign t[104] = t[140] ^ t[141];
  assign t[105] = t[142] & t[143];
  assign t[106] = ~(t[105] ^ t[144]);
  assign t[107] = t[18] ^ t[145];
  assign t[108] = ~(t[146] & t[147]);
  assign t[109] = t[148] ^ t[209];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = ~(t[202]);
  assign t[111] = t[149] & t[148];
  assign t[112] = ~(t[49]);
  assign t[113] = t[112] ? x[70] : x[69];
  assign t[114] = t[203] ^ t[150];
  assign t[115] = t[112] ? x[72] : x[71];
  assign t[116] = t[101] ^ t[122];
  assign t[117] = t[151] & t[141];
  assign t[118] = t[32] ^ t[54];
  assign t[119] = t[152] & t[153];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[127] ^ t[154];
  assign t[121] = t[155] ^ t[89];
  assign t[122] = t[136] ? t[156] : t[210];
  assign t[123] = t[139] ^ t[69];
  assign t[124] = t[204] ^ t[157];
  assign t[125] = t[205] ^ t[158];
  assign t[126] = t[159] ^ t[160];
  assign t[127] = t[86] ^ t[99];
  assign t[128] = t[7] ? t[161] : t[211];
  assign t[129] = ~(t[155] ^ t[41]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[22] ^ t[95];
  assign t[131] = t[112] ? x[80] : x[79];
  assign t[132] = t[75] ? x[82] : x[81];
  assign t[133] = t[162];
  assign t[134] = t[7] ? t[163] : t[212];
  assign t[135] = t[206] ^ t[164];
  assign t[136] = ~(t[14]);
  assign t[137] = t[207] ^ t[165];
  assign t[138] = t[208] ^ t[166];
  assign t[139] = t[167] ^ t[117];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[102] ^ t[122];
  assign t[141] = t[136] ? t[168] : t[213];
  assign t[142] = ~(t[145]);
  assign t[143] = ~(t[32]);
  assign t[144] = t[45] ^ t[32];
  assign t[145] = t[35] ^ t[54];
  assign t[146] = ~(t[149] | t[148]);
  assign t[147] = ~(t[169] | t[110]);
  assign t[148] = ~(t[214]);
  assign t[149] = ~(t[209]);
  assign t[14] = ~(t[26]);
  assign t[150] = t[112] ? x[93] : x[92];
  assign t[151] = ~(t[102]);
  assign t[152] = ~(t[118] ^ t[70]);
  assign t[153] = t[45] ^ t[35];
  assign t[154] = t[126] ^ t[170];
  assign t[155] = t[133] ^ t[39];
  assign t[156] = t[210] ^ t[171];
  assign t[157] = t[27] ? x[95] : x[94];
  assign t[158] = t[27] ? x[97] : x[96];
  assign t[159] = t[172] & t[173];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[174] & t[128];
  assign t[161] = t[211] ^ t[175];
  assign t[162] = t[7] ? t[176] : t[215];
  assign t[163] = t[212] ^ t[177];
  assign t[164] = t[75] ? x[102] : x[101];
  assign t[165] = t[178] ? x[104] : x[103];
  assign t[166] = t[178] ? x[106] : x[105];
  assign t[167] = t[179] & t[180];
  assign t[168] = t[213] ^ t[181];
  assign t[169] = ~(t[196]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[182] & t[183];
  assign t[171] = t[178] ? x[108] : x[107];
  assign t[172] = ~(t[184]);
  assign t[173] = ~(t[85]);
  assign t[174] = ~(t[86]);
  assign t[175] = t[27] ? x[110] : x[109];
  assign t[176] = t[215] ^ t[185];
  assign t[177] = t[75] ? x[112] : x[111];
  assign t[178] = ~(t[49]);
  assign t[179] = ~(t[186]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = ~(t[101]);
  assign t[181] = t[178] ? x[114] : x[113];
  assign t[182] = ~(t[159] ^ t[187]);
  assign t[183] = t[188] ^ t[184];
  assign t[184] = t[128] ^ t[86];
  assign t[185] = t[75] ? x[116] : x[115];
  assign t[186] = t[141] ^ t[102];
  assign t[187] = t[127] ^ t[85];
  assign t[188] = t[85] ^ t[99];
  assign t[189] = t[216] ^ x[4];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[217] ^ x[9];
  assign t[191] = t[218] ^ x[12];
  assign t[192] = t[219] ^ x[15];
  assign t[193] = t[220] ^ x[18];
  assign t[194] = t[221] ^ x[21];
  assign t[195] = t[222] ^ x[24];
  assign t[196] = t[223] ^ x[27];
  assign t[197] = t[224] ^ x[30];
  assign t[198] = t[225] ^ x[33];
  assign t[199] = t[226] ^ x[36];
  assign t[19] = t[34] & t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[39];
  assign t[201] = t[228] ^ x[42];
  assign t[202] = t[229] ^ x[45];
  assign t[203] = t[230] ^ x[50];
  assign t[204] = t[231] ^ x[53];
  assign t[205] = t[232] ^ x[56];
  assign t[206] = t[233] ^ x[59];
  assign t[207] = t[234] ^ x[62];
  assign t[208] = t[235] ^ x[65];
  assign t[209] = t[236] ^ x[68];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[75];
  assign t[211] = t[238] ^ x[78];
  assign t[212] = t[239] ^ x[85];
  assign t[213] = t[240] ^ x[88];
  assign t[214] = t[241] ^ x[91];
  assign t[215] = t[242] ^ x[100];
  assign t[216] = (x[2] & x[3]);
  assign t[217] = (x[7] & x[8]);
  assign t[218] = (x[10] & x[11]);
  assign t[219] = (x[13] & x[14]);
  assign t[21] = ~(t[25] ^ t[38]);
  assign t[220] = (x[16] & x[17]);
  assign t[221] = (x[19] & x[20]);
  assign t[222] = (x[22] & x[23]);
  assign t[223] = (x[25] & x[26]);
  assign t[224] = (x[28] & x[29]);
  assign t[225] = (x[31] & x[32]);
  assign t[226] = (x[34] & x[35]);
  assign t[227] = (x[37] & x[38]);
  assign t[228] = (x[40] & x[41]);
  assign t[229] = (x[43] & x[44]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (x[48] & x[49]);
  assign t[231] = (x[51] & x[52]);
  assign t[232] = (x[54] & x[55]);
  assign t[233] = (x[57] & x[58]);
  assign t[234] = (x[60] & x[61]);
  assign t[235] = (x[63] & x[64]);
  assign t[236] = (x[66] & x[67]);
  assign t[237] = (x[73] & x[74]);
  assign t[238] = (x[76] & x[77]);
  assign t[239] = (x[83] & x[84]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (x[86] & x[87]);
  assign t[241] = (x[89] & x[90]);
  assign t[242] = (x[98] & x[99]);
  assign t[24] = ~(t[43] ^ t[44]);
  assign t[25] = t[45] ^ t[46];
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49]);
  assign t[28] = ~(t[190]);
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[192]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = t[7] ? t[52] : t[193];
  assign t[33] = t[194] ^ t[53];
  assign t[34] = ~(t[54]);
  assign t[35] = t[195] ^ t[55];
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[37] = t[58] ^ t[59];
  assign t[38] = t[40] ^ t[60];
  assign t[39] = ~t[61];
  assign t[3] = t[7] ? t[8] : t[189];
  assign t[40] = t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[12] ^ t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[54] ^ t[33];
  assign t[46] = t[70] ^ t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[196] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[194]);
  assign t[51] = ~(t[76] & t[197]);
  assign t[52] = t[193] ^ t[77];
  assign t[53] = t[7] ? t[78] : t[198];
  assign t[54] = t[192] ^ t[79];
  assign t[55] = t[7] ? t[80] : t[199];
  assign t[56] = t[81] ^ t[82];
  assign t[57] = ~(t[83] ^ t[84]);
  assign t[58] = t[85] ^ t[86];
  assign t[59] = t[87] & t[88];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[41] ^ t[89];
  assign t[61] = t[7] ? t[90] : t[200];
  assign t[62] = t[7] ? t[91] : t[201];
  assign t[63] = t[92] & t[93];
  assign t[64] = t[94] & t[95];
  assign t[65] = ~(t[63] ^ t[96]);
  assign t[66] = t[97] ^ t[98];
  assign t[67] = t[99] ^ t[100];
  assign t[68] = t[101] ^ t[102];
  assign t[69] = t[103] & t[104];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[105] ^ t[19];
  assign t[71] = t[106] & t[107];
  assign t[72] = ~(t[74] & t[108]);
  assign t[73] = ~(t[202] ^ t[109]);
  assign t[74] = ~(t[110] & t[111]);
  assign t[75] = ~(t[48]);
  assign t[76] = ~(t[195]);
  assign t[77] = t[112] ? x[47] : x[46];
  assign t[78] = t[198] ^ t[113];
  assign t[79] = t[7] ? t[114] : t[203];
  assign t[7] = ~(t[14]);
  assign t[80] = t[199] ^ t[115];
  assign t[81] = t[116] ^ t[117];
  assign t[82] = t[118] ^ t[119];
  assign t[83] = t[120] ^ t[121];
  assign t[84] = t[122] ^ t[123];
  assign t[85] = t[7] ? t[124] : t[204];
  assign t[86] = t[7] ? t[125] : t[205];
  assign t[87] = ~(t[58] ^ t[126]);
  assign t[88] = t[127] ^ t[128];
  assign t[89] = t[129] & t[130];
  assign t[8] = t[189] ^ t[15];
  assign t[90] = t[200] ^ t[131];
  assign t[91] = t[201] ^ t[132];
  assign t[92] = ~(t[98]);
  assign t[93] = ~(t[133]);
  assign t[94] = ~(t[39]);
  assign t[95] = t[134];
  assign t[96] = t[22] ^ t[133];
  assign t[97] = t[133] ^ t[40];
  assign t[98] = t[95] ^ t[39];
  assign t[99] = t[7] ? t[135] : t[206];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind90(x, y);
 input [116:0] x;
 output y;

 wire [249:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[137];
  assign t[101] = t[87] ^ t[22];
  assign t[102] = t[135] ? x[61] : x[60];
  assign t[103] = t[135] ? x[63] : x[62];
  assign t[104] = t[138] & t[139];
  assign t[105] = t[140] & t[71];
  assign t[106] = t[7] ? t[141] : t[214];
  assign t[107] = t[206] ^ t[142];
  assign t[108] = ~(t[143] & t[144]);
  assign t[109] = t[145] ^ t[215];
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = ~(t[207]);
  assign t[111] = t[146] & t[145];
  assign t[112] = t[147] ^ t[64];
  assign t[113] = ~(t[148] ^ t[38]);
  assign t[114] = t[149] ^ t[150];
  assign t[115] = t[42] ^ t[106];
  assign t[116] = t[69] ^ t[25];
  assign t[117] = t[209] ^ t[151];
  assign t[118] = t[210] ^ t[152];
  assign t[119] = t[26] ? t[153] : t[216];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[211] ^ t[154];
  assign t[121] = t[155] & t[156];
  assign t[122] = t[157] ^ t[53];
  assign t[123] = t[158] & t[159];
  assign t[124] = t[7] ? t[160] : t[217];
  assign t[125] = t[7] ? t[161] : t[218];
  assign t[126] = ~(t[14]);
  assign t[127] = t[212] ^ t[162];
  assign t[128] = t[197] ^ t[163];
  assign t[129] = t[126] ? t[164] : t[219];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[165] & t[166];
  assign t[131] = t[213] ^ t[167];
  assign t[132] = t[168] & t[169];
  assign t[133] = ~(t[170] ^ t[94]);
  assign t[134] = t[149] ^ t[90];
  assign t[135] = ~(t[171]);
  assign t[136] = t[100] ^ t[87];
  assign t[137] = t[26] ? t[172] : t[220];
  assign t[138] = ~(t[173]);
  assign t[139] = ~(t[42]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[43]);
  assign t[141] = t[214] ^ t[174];
  assign t[142] = t[135] ? x[86] : x[85];
  assign t[143] = ~(t[146] | t[145]);
  assign t[144] = ~(t[175] | t[110]);
  assign t[145] = ~(t[221]);
  assign t[146] = ~(t[215]);
  assign t[147] = t[86] ^ t[22];
  assign t[148] = t[176] ^ t[123];
  assign t[149] = t[128] ^ t[60];
  assign t[14] = ~(t[26]);
  assign t[150] = t[94] ^ t[177];
  assign t[151] = t[178] ? x[91] : x[90];
  assign t[152] = t[27] ? x[93] : x[92];
  assign t[153] = t[216] ^ t[179];
  assign t[154] = t[27] ? x[95] : x[94];
  assign t[155] = ~(t[104] ^ t[180]);
  assign t[156] = t[115] ^ t[173];
  assign t[157] = t[181] & t[182];
  assign t[158] = ~(t[176] ^ t[122]);
  assign t[159] = t[91] ^ t[83];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[217] ^ t[183];
  assign t[161] = t[218] ^ t[184];
  assign t[162] = t[185] ? x[97] : x[96];
  assign t[163] = t[126] ? t[186] : t[222];
  assign t[164] = t[219] ^ t[187];
  assign t[165] = ~(t[157] ^ t[188]);
  assign t[166] = t[52] ^ t[189];
  assign t[167] = t[185] ? x[102] : x[101];
  assign t[168] = ~(t[190]);
  assign t[169] = ~(t[88]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[88] ^ t[128];
  assign t[171] = ~(t[27]);
  assign t[172] = t[220] ^ t[191];
  assign t[173] = t[71] ^ t[43];
  assign t[174] = t[135] ? x[104] : x[103];
  assign t[175] = ~(t[203]);
  assign t[176] = t[80] ^ t[119];
  assign t[177] = t[192] & t[193];
  assign t[178] = ~(t[171]);
  assign t[179] = t[178] ? x[106] : x[105];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[70] ^ t[42];
  assign t[181] = ~(t[189]);
  assign t[182] = ~(t[80]);
  assign t[183] = t[135] ? x[108] : x[107];
  assign t[184] = t[135] ? x[110] : x[109];
  assign t[185] = ~(t[171]);
  assign t[186] = t[222] ^ t[194];
  assign t[187] = t[185] ? x[112] : x[111];
  assign t[188] = t[91] ^ t[80];
  assign t[189] = t[83] ^ t[119];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[90] ^ t[128];
  assign t[191] = t[135] ? x[114] : x[113];
  assign t[192] = ~(t[132] ^ t[195]);
  assign t[193] = t[57] ^ t[190];
  assign t[194] = t[185] ? x[116] : x[115];
  assign t[195] = t[149] ^ t[88];
  assign t[196] = t[223] ^ x[4];
  assign t[197] = t[224] ^ x[9];
  assign t[198] = t[225] ^ x[12];
  assign t[199] = t[226] ^ x[15];
  assign t[19] = ~(t[34] ^ t[35]);
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[18];
  assign t[201] = t[228] ^ x[21];
  assign t[202] = t[229] ^ x[24];
  assign t[203] = t[230] ^ x[27];
  assign t[204] = t[231] ^ x[30];
  assign t[205] = t[232] ^ x[33];
  assign t[206] = t[233] ^ x[36];
  assign t[207] = t[234] ^ x[39];
  assign t[208] = t[235] ^ x[42];
  assign t[209] = t[236] ^ x[45];
  assign t[20] = t[36] ^ t[35];
  assign t[210] = t[237] ^ x[48];
  assign t[211] = t[238] ^ x[51];
  assign t[212] = t[239] ^ x[54];
  assign t[213] = t[240] ^ x[57];
  assign t[214] = t[241] ^ x[66];
  assign t[215] = t[242] ^ x[69];
  assign t[216] = t[243] ^ x[72];
  assign t[217] = t[244] ^ x[75];
  assign t[218] = t[245] ^ x[78];
  assign t[219] = t[246] ^ x[81];
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = t[247] ^ x[84];
  assign t[221] = t[248] ^ x[89];
  assign t[222] = t[249] ^ x[100];
  assign t[223] = (x[2] & x[3]);
  assign t[224] = (x[7] & x[8]);
  assign t[225] = (x[10] & x[11]);
  assign t[226] = (x[13] & x[14]);
  assign t[227] = (x[16] & x[17]);
  assign t[228] = (x[19] & x[20]);
  assign t[229] = (x[22] & x[23]);
  assign t[22] = ~t[39];
  assign t[230] = (x[25] & x[26]);
  assign t[231] = (x[28] & x[29]);
  assign t[232] = (x[31] & x[32]);
  assign t[233] = (x[34] & x[35]);
  assign t[234] = (x[37] & x[38]);
  assign t[235] = (x[40] & x[41]);
  assign t[236] = (x[43] & x[44]);
  assign t[237] = (x[46] & x[47]);
  assign t[238] = (x[49] & x[50]);
  assign t[239] = (x[52] & x[53]);
  assign t[23] = t[40] ^ t[41];
  assign t[240] = (x[55] & x[56]);
  assign t[241] = (x[64] & x[65]);
  assign t[242] = (x[67] & x[68]);
  assign t[243] = (x[70] & x[71]);
  assign t[244] = (x[73] & x[74]);
  assign t[245] = (x[76] & x[77]);
  assign t[246] = (x[79] & x[80]);
  assign t[247] = (x[82] & x[83]);
  assign t[248] = (x[87] & x[88]);
  assign t[249] = (x[98] & x[99]);
  assign t[24] = t[42] ^ t[43];
  assign t[25] = t[44] & t[45];
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[197]);
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[199]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = ~(t[50] ^ t[51]);
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] ^ t[41];
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ t[13];
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[7] ? t[62] : t[200];
  assign t[3] = t[7] ? t[8] : t[196];
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65] & t[66];
  assign t[42] = t[7] ? t[67] : t[201];
  assign t[43] = t[7] ? t[68] : t[202];
  assign t[44] = ~(t[24] ^ t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[203] | t[74];
  assign t[48] = ~(t[204]);
  assign t[49] = ~(t[75] & t[205]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[76] ^ t[77];
  assign t[51] = ~(t[78] ^ t[79]);
  assign t[52] = t[80] ^ t[81];
  assign t[53] = t[82] & t[83];
  assign t[54] = t[70] ^ t[84];
  assign t[55] = t[81] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ^ t[60];
  assign t[58] = t[89] & t[90];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[205] ^ t[93];
  assign t[61] = t[94] ^ t[95];
  assign t[62] = t[200] ^ t[96];
  assign t[63] = t[97] & t[98];
  assign t[64] = t[99] & t[100];
  assign t[65] = ~(t[56] ^ t[40]);
  assign t[66] = t[101] ^ t[100];
  assign t[67] = t[201] ^ t[102];
  assign t[68] = t[202] ^ t[103];
  assign t[69] = t[104] ^ t[105];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[43] ^ t[106];
  assign t[71] = t[7] ? t[107] : t[206];
  assign t[72] = ~(t[74] & t[108]);
  assign t[73] = ~(t[207] ^ t[109]);
  assign t[74] = ~(t[110] & t[111]);
  assign t[75] = ~(t[208]);
  assign t[76] = t[12] ^ t[112];
  assign t[77] = ~(t[113] ^ t[114]);
  assign t[78] = t[115] ^ t[105];
  assign t[79] = t[106] ^ t[116];
  assign t[7] = ~(t[14]);
  assign t[80] = t[26] ? t[117] : t[209];
  assign t[81] = t[26] ? t[118] : t[210];
  assign t[82] = ~(t[119]);
  assign t[83] = t[26] ? t[120] : t[211];
  assign t[84] = t[69] ^ t[121];
  assign t[85] = t[122] ^ t[123];
  assign t[86] = t[124];
  assign t[87] = ~t[125];
  assign t[88] = t[126] ? t[127] : t[212];
  assign t[89] = ~(t[128]);
  assign t[8] = t[196] ^ t[15];
  assign t[90] = t[198] ^ t[129];
  assign t[91] = t[119] ^ t[81];
  assign t[92] = t[122] ^ t[130];
  assign t[93] = t[126] ? t[131] : t[213];
  assign t[94] = t[132] ^ t[58];
  assign t[95] = t[133] & t[134];
  assign t[96] = t[135] ? x[59] : x[58];
  assign t[97] = ~(t[136]);
  assign t[98] = ~(t[86]);
  assign t[99] = ~(t[87]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind91(x, y);
 input [116:0] x;
 output y;

 wire [249:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[136] ^ t[137];
  assign t[101] = t[79] ? x[53] : x[52];
  assign t[102] = t[138] & t[139];
  assign t[103] = t[140] & t[125];
  assign t[104] = t[141] & t[142];
  assign t[105] = t[7] ? t[143] : t[212];
  assign t[106] = t[7] ? t[144] : t[213];
  assign t[107] = ~(t[69] ^ t[145]);
  assign t[108] = t[146] ^ t[147];
  assign t[109] = t[146] ^ t[148];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[149] ^ t[62];
  assign t[111] = t[90] ^ t[40];
  assign t[112] = t[34] ^ t[150];
  assign t[113] = t[7] ? t[151] : t[214];
  assign t[114] = t[145] ^ t[70];
  assign t[115] = ~(t[152] & t[153]);
  assign t[116] = t[154] ^ t[215];
  assign t[117] = ~(t[206]);
  assign t[118] = t[155] & t[154];
  assign t[119] = t[27] ? x[67] : x[66];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[27] ? x[69] : x[68];
  assign t[121] = t[156];
  assign t[122] = t[26] ? t[157] : t[216];
  assign t[123] = t[208] ^ t[158];
  assign t[124] = t[209] ^ t[159];
  assign t[125] = t[26] ? t[160] : t[217];
  assign t[126] = ~(t[14]);
  assign t[127] = t[210] ^ t[161];
  assign t[128] = ~(t[110] ^ t[63]);
  assign t[129] = t[38] ^ t[134];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[211] ^ t[162];
  assign t[131] = ~(t[137]);
  assign t[132] = ~(t[149]);
  assign t[133] = ~(t[62]);
  assign t[134] = t[198] ^ t[163];
  assign t[135] = t[38] ^ t[149];
  assign t[136] = t[149] ^ t[60];
  assign t[137] = t[134] ^ t[62];
  assign t[138] = ~(t[164]);
  assign t[139] = ~(t[90]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[91]);
  assign t[141] = ~(t[102] ^ t[165]);
  assign t[142] = t[111] ^ t[164];
  assign t[143] = t[212] ^ t[166];
  assign t[144] = t[213] ^ t[167];
  assign t[145] = t[168] ^ t[169];
  assign t[146] = t[106] ^ t[113];
  assign t[147] = t[7] ? t[170] : t[218];
  assign t[148] = t[145] ^ t[171];
  assign t[149] = t[126] ? t[172] : t[219];
  assign t[14] = ~(t[26]);
  assign t[150] = t[173] & t[174];
  assign t[151] = t[214] ^ t[175];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[176] | t[117]);
  assign t[154] = ~(t[220]);
  assign t[155] = ~(t[215]);
  assign t[156] = t[7] ? t[177] : t[221];
  assign t[157] = t[216] ^ t[178];
  assign t[158] = t[179] ? x[89] : x[88];
  assign t[159] = t[179] ? x[91] : x[90];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[217] ^ t[180];
  assign t[161] = t[181] ? x[93] : x[92];
  assign t[162] = t[181] ? x[95] : x[94];
  assign t[163] = t[126] ? t[182] : t[222];
  assign t[164] = t[125] ^ t[91];
  assign t[165] = t[67] ^ t[90];
  assign t[166] = t[27] ? x[100] : x[99];
  assign t[167] = t[27] ? x[102] : x[101];
  assign t[168] = t[183] & t[184];
  assign t[169] = t[185] & t[147];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[218] ^ t[186];
  assign t[171] = t[187] & t[188];
  assign t[172] = t[219] ^ t[189];
  assign t[173] = ~(t[190] ^ t[34]);
  assign t[174] = t[18] ^ t[86];
  assign t[175] = t[27] ? x[104] : x[103];
  assign t[176] = ~(t[201]);
  assign t[177] = t[221] ^ t[191];
  assign t[178] = t[27] ? x[106] : x[105];
  assign t[179] = ~(t[49]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[79] ? x[108] : x[107];
  assign t[181] = ~(t[49]);
  assign t[182] = t[222] ^ t[192];
  assign t[183] = ~(t[193]);
  assign t[184] = ~(t[105]);
  assign t[185] = ~(t[106]);
  assign t[186] = t[27] ? x[110] : x[109];
  assign t[187] = ~(t[168] ^ t[194]);
  assign t[188] = t[195] ^ t[193];
  assign t[189] = t[181] ? x[112] : x[111];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[121] ^ t[32];
  assign t[191] = t[27] ? x[114] : x[113];
  assign t[192] = t[181] ? x[116] : x[115];
  assign t[193] = t[147] ^ t[106];
  assign t[194] = t[146] ^ t[105];
  assign t[195] = t[105] ^ t[113];
  assign t[196] = t[223] ^ x[4];
  assign t[197] = t[224] ^ x[9];
  assign t[198] = t[225] ^ x[12];
  assign t[199] = t[226] ^ x[15];
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[18];
  assign t[201] = t[228] ^ x[21];
  assign t[202] = t[229] ^ x[24];
  assign t[203] = t[230] ^ x[27];
  assign t[204] = t[231] ^ x[30];
  assign t[205] = t[232] ^ x[33];
  assign t[206] = t[233] ^ x[36];
  assign t[207] = t[234] ^ x[39];
  assign t[208] = t[235] ^ x[42];
  assign t[209] = t[236] ^ x[45];
  assign t[20] = ~(t[36] ^ t[37]);
  assign t[210] = t[237] ^ x[48];
  assign t[211] = t[238] ^ x[51];
  assign t[212] = t[239] ^ x[56];
  assign t[213] = t[240] ^ x[59];
  assign t[214] = t[241] ^ x[62];
  assign t[215] = t[242] ^ x[65];
  assign t[216] = t[243] ^ x[72];
  assign t[217] = t[244] ^ x[75];
  assign t[218] = t[245] ^ x[78];
  assign t[219] = t[246] ^ x[81];
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[247] ^ x[84];
  assign t[221] = t[248] ^ x[87];
  assign t[222] = t[249] ^ x[98];
  assign t[223] = (x[2] & x[3]);
  assign t[224] = (x[7] & x[8]);
  assign t[225] = (x[10] & x[11]);
  assign t[226] = (x[13] & x[14]);
  assign t[227] = (x[16] & x[17]);
  assign t[228] = (x[19] & x[20]);
  assign t[229] = (x[22] & x[23]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (x[25] & x[26]);
  assign t[231] = (x[28] & x[29]);
  assign t[232] = (x[31] & x[32]);
  assign t[233] = (x[34] & x[35]);
  assign t[234] = (x[37] & x[38]);
  assign t[235] = (x[40] & x[41]);
  assign t[236] = (x[43] & x[44]);
  assign t[237] = (x[46] & x[47]);
  assign t[238] = (x[49] & x[50]);
  assign t[239] = (x[54] & x[55]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (x[57] & x[58]);
  assign t[241] = (x[60] & x[61]);
  assign t[242] = (x[63] & x[64]);
  assign t[243] = (x[70] & x[71]);
  assign t[244] = (x[73] & x[74]);
  assign t[245] = (x[76] & x[77]);
  assign t[246] = (x[79] & x[80]);
  assign t[247] = (x[82] & x[83]);
  assign t[248] = (x[85] & x[86]);
  assign t[249] = (x[96] & x[97]);
  assign t[24] = ~(t[44] ^ t[10]);
  assign t[25] = ~(t[45] ^ t[46]);
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49]);
  assign t[28] = ~(t[197]);
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[199]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~t[52];
  assign t[33] = ~t[53];
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] & t[57];
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[62] ^ t[60];
  assign t[39] = t[63] ^ t[64];
  assign t[3] = t[7] ? t[8] : t[196];
  assign t[40] = t[26] ? t[65] : t[200];
  assign t[41] = t[66] ^ t[59];
  assign t[42] = t[67] ^ t[68];
  assign t[43] = t[69] ^ t[70];
  assign t[44] = ~(t[71] ^ t[72]);
  assign t[45] = t[21] ^ t[73];
  assign t[46] = ~(t[74] ^ t[75]);
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = t[201] | t[78];
  assign t[49] = ~(t[79]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[202]);
  assign t[51] = ~(t[80] & t[203]);
  assign t[52] = t[7] ? t[81] : t[204];
  assign t[53] = t[7] ? t[82] : t[205];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[85] & t[86];
  assign t[56] = ~(t[54] ^ t[87]);
  assign t[57] = t[88] ^ t[89];
  assign t[58] = t[90] ^ t[91];
  assign t[59] = t[92] & t[93];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[203] ^ t[94];
  assign t[61] = t[63] ^ t[95];
  assign t[62] = t[197] ^ t[96];
  assign t[63] = t[97] ^ t[98];
  assign t[64] = t[99] & t[100];
  assign t[65] = t[200] ^ t[101];
  assign t[66] = t[102] ^ t[103];
  assign t[67] = t[91] ^ t[40];
  assign t[68] = t[66] ^ t[104];
  assign t[69] = t[105] ^ t[106];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[107] & t[108];
  assign t[71] = t[109] ^ t[22];
  assign t[72] = t[110] ^ t[95];
  assign t[73] = t[111] ^ t[103];
  assign t[74] = t[33] ^ t[112];
  assign t[75] = t[113] ^ t[114];
  assign t[76] = ~(t[78] & t[115]);
  assign t[77] = ~(t[206] ^ t[116]);
  assign t[78] = ~(t[117] & t[118]);
  assign t[79] = ~(t[48]);
  assign t[7] = ~(t[14]);
  assign t[80] = ~(t[207]);
  assign t[81] = t[204] ^ t[119];
  assign t[82] = t[205] ^ t[120];
  assign t[83] = ~(t[89]);
  assign t[84] = ~(t[121]);
  assign t[85] = ~(t[32]);
  assign t[86] = t[122];
  assign t[87] = t[18] ^ t[121];
  assign t[88] = t[121] ^ t[33];
  assign t[89] = t[86] ^ t[32];
  assign t[8] = t[196] ^ t[15];
  assign t[90] = t[26] ? t[123] : t[208];
  assign t[91] = t[26] ? t[124] : t[209];
  assign t[92] = ~(t[58] ^ t[66]);
  assign t[93] = t[67] ^ t[125];
  assign t[94] = t[126] ? t[127] : t[210];
  assign t[95] = t[128] & t[129];
  assign t[96] = t[126] ? t[130] : t[211];
  assign t[97] = t[131] & t[132];
  assign t[98] = t[133] & t[134];
  assign t[99] = ~(t[97] ^ t[135]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind92(x, y);
 input [116:0] x;
 output y;

 wire [260:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[30] ? x[50] : x[49];
  assign t[101] = ~(t[136] ^ t[64]);
  assign t[102] = t[39] ^ t[105];
  assign t[103] = t[66] ? t[137] : t[222];
  assign t[104] = ~(t[63]);
  assign t[105] = t[66] ? t[138] : t[223];
  assign t[106] = t[7] ? t[139] : t[224];
  assign t[107] = t[7] ? t[140] : t[225];
  assign t[108] = t[141] ^ t[125];
  assign t[109] = t[142] & t[143];
  assign t[10] = t[19] ^ t[20];
  assign t[110] = t[66] ? t[144] : t[226];
  assign t[111] = t[145] ^ t[146];
  assign t[112] = t[44] ^ t[147];
  assign t[113] = t[148] ^ t[149];
  assign t[114] = t[7] ? t[150] : t[227];
  assign t[115] = ~(t[77] ^ t[108]);
  assign t[116] = t[71] ^ t[151];
  assign t[117] = t[152] & t[153];
  assign t[118] = ~(t[208]);
  assign t[119] = t[107] ^ t[154];
  assign t[11] = ~(t[21] ^ t[22]);
  assign t[120] = t[155] ^ t[156];
  assign t[121] = t[157] & t[158];
  assign t[122] = t[156] ^ t[148];
  assign t[123] = t[159] ^ t[160];
  assign t[124] = t[114] ^ t[107];
  assign t[125] = t[161] & t[151];
  assign t[126] = t[220] ^ t[162];
  assign t[127] = t[221] ^ t[163];
  assign t[128] = t[164] & t[165];
  assign t[129] = t[166] & t[94];
  assign t[12] = ~(t[23] ^ t[24]);
  assign t[130] = t[7] ? t[167] : t[228];
  assign t[131] = t[30] ? x[73] : x[72];
  assign t[132] = ~(t[135]);
  assign t[133] = ~(t[103]);
  assign t[134] = t[39] ^ t[103];
  assign t[135] = t[105] ^ t[63];
  assign t[136] = t[103] ^ t[63];
  assign t[137] = t[222] ^ t[168];
  assign t[138] = t[223] ^ t[169];
  assign t[139] = t[224] ^ t[170];
  assign t[13] = ~(t[25] ^ t[26]);
  assign t[140] = t[225] ^ t[171];
  assign t[141] = t[172] & t[173];
  assign t[142] = ~(t[141] ^ t[174]);
  assign t[143] = t[124] ^ t[175];
  assign t[144] = t[226] ^ t[176];
  assign t[145] = t[155] ^ t[148];
  assign t[146] = t[177] & t[178];
  assign t[147] = t[136] ^ t[68];
  assign t[148] = t[216] ^ t[179];
  assign t[149] = t[159] ^ t[121];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[227] ^ t[180];
  assign t[151] = t[7] ? t[181] : t[229];
  assign t[152] = ~(t[128] ^ t[182]);
  assign t[153] = t[183] ^ t[184];
  assign t[154] = t[108] ^ t[78];
  assign t[155] = t[185] ? t[186] : t[230];
  assign t[156] = t[210] ^ t[187];
  assign t[157] = ~(t[120] ^ t[159]);
  assign t[158] = t[122] ^ t[178];
  assign t[159] = t[188] ^ t[146];
  assign t[15] = t[208] | t[29];
  assign t[160] = t[189] & t[190];
  assign t[161] = ~(t[106]);
  assign t[162] = t[30] ? x[81] : x[80];
  assign t[163] = t[30] ? x[83] : x[82];
  assign t[164] = ~(t[184]);
  assign t[165] = ~(t[59]);
  assign t[166] = ~(t[60]);
  assign t[167] = t[228] ^ t[191];
  assign t[168] = t[30] ? x[85] : x[84];
  assign t[169] = t[30] ? x[87] : x[86];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[192] ? x[89] : x[88];
  assign t[171] = t[85] ? x[91] : x[90];
  assign t[172] = ~(t[175]);
  assign t[173] = ~(t[114]);
  assign t[174] = t[71] ^ t[114];
  assign t[175] = t[151] ^ t[106];
  assign t[176] = t[30] ? x[93] : x[92];
  assign t[177] = ~(t[156]);
  assign t[178] = t[211] ^ t[193];
  assign t[179] = t[185] ? t[194] : t[231];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[192] ? x[98] : x[97];
  assign t[181] = t[229] ^ t[195];
  assign t[182] = t[79] ^ t[59];
  assign t[183] = t[59] ^ t[73];
  assign t[184] = t[94] ^ t[60];
  assign t[185] = ~(t[99]);
  assign t[186] = t[230] ^ t[196];
  assign t[187] = t[185] ? t[197] : t[232];
  assign t[188] = t[198] & t[199];
  assign t[189] = ~(t[188] ^ t[200]);
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[145] ^ t[201];
  assign t[191] = t[30] ? x[103] : x[102];
  assign t[192] = ~(t[53]);
  assign t[193] = t[185] ? t[202] : t[233];
  assign t[194] = t[231] ^ t[203];
  assign t[195] = t[85] ? x[108] : x[107];
  assign t[196] = t[204] ? x[110] : x[109];
  assign t[197] = t[232] ^ t[205];
  assign t[198] = ~(t[201]);
  assign t[199] = ~(t[155]);
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = t[122] ^ t[155];
  assign t[201] = t[178] ^ t[156];
  assign t[202] = t[233] ^ t[206];
  assign t[203] = t[204] ? x[112] : x[111];
  assign t[204] = ~(t[53]);
  assign t[205] = t[204] ? x[114] : x[113];
  assign t[206] = t[204] ? x[116] : x[115];
  assign t[207] = t[234] ^ x[4];
  assign t[208] = t[235] ^ x[7];
  assign t[209] = t[236] ^ x[12];
  assign t[20] = t[37] ^ t[38];
  assign t[210] = t[237] ^ x[15];
  assign t[211] = t[238] ^ x[18];
  assign t[212] = t[239] ^ x[21];
  assign t[213] = t[240] ^ x[24];
  assign t[214] = t[241] ^ x[27];
  assign t[215] = t[242] ^ x[30];
  assign t[216] = t[243] ^ x[33];
  assign t[217] = t[244] ^ x[36];
  assign t[218] = t[245] ^ x[39];
  assign t[219] = t[246] ^ x[42];
  assign t[21] = t[39] ^ t[40];
  assign t[220] = t[247] ^ x[45];
  assign t[221] = t[248] ^ x[48];
  assign t[222] = t[249] ^ x[53];
  assign t[223] = t[250] ^ x[56];
  assign t[224] = t[251] ^ x[59];
  assign t[225] = t[252] ^ x[62];
  assign t[226] = t[253] ^ x[65];
  assign t[227] = t[254] ^ x[68];
  assign t[228] = t[255] ^ x[71];
  assign t[229] = t[256] ^ x[76];
  assign t[22] = t[41] ^ t[42];
  assign t[230] = t[257] ^ x[79];
  assign t[231] = t[258] ^ x[96];
  assign t[232] = t[259] ^ x[101];
  assign t[233] = t[260] ^ x[106];
  assign t[234] = (x[2] & x[3]);
  assign t[235] = (x[5] & x[6]);
  assign t[236] = (x[10] & x[11]);
  assign t[237] = (x[13] & x[14]);
  assign t[238] = (x[16] & x[17]);
  assign t[239] = (x[19] & x[20]);
  assign t[23] = t[43] ^ t[44];
  assign t[240] = (x[22] & x[23]);
  assign t[241] = (x[25] & x[26]);
  assign t[242] = (x[28] & x[29]);
  assign t[243] = (x[31] & x[32]);
  assign t[244] = (x[34] & x[35]);
  assign t[245] = (x[37] & x[38]);
  assign t[246] = (x[40] & x[41]);
  assign t[247] = (x[43] & x[44]);
  assign t[248] = (x[46] & x[47]);
  assign t[249] = (x[51] & x[52]);
  assign t[24] = ~(t[35] ^ t[45]);
  assign t[250] = (x[54] & x[55]);
  assign t[251] = (x[57] & x[58]);
  assign t[252] = (x[60] & x[61]);
  assign t[253] = (x[63] & x[64]);
  assign t[254] = (x[66] & x[67]);
  assign t[255] = (x[69] & x[70]);
  assign t[256] = (x[74] & x[75]);
  assign t[257] = (x[77] & x[78]);
  assign t[258] = (x[94] & x[95]);
  assign t[259] = (x[99] & x[100]);
  assign t[25] = t[46] ^ t[47];
  assign t[260] = (x[104] & x[105]);
  assign t[26] = ~(t[48] ^ t[22]);
  assign t[27] = ~(t[29] & t[49]);
  assign t[28] = ~(t[209] ^ t[50]);
  assign t[29] = ~(t[51] & t[52]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[53]);
  assign t[31] = ~(t[210]);
  assign t[32] = ~(t[211]);
  assign t[33] = ~(t[212]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = ~(t[56] ^ t[48]);
  assign t[36] = ~(t[57] ^ t[58]);
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[61] & t[62];
  assign t[39] = t[63] ^ t[41];
  assign t[3] = t[7] ? t[8] : t[207];
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[66] ? t[67] : t[213];
  assign t[42] = t[64] ^ t[68];
  assign t[43] = t[69] ^ t[70];
  assign t[44] = t[71] ^ t[72];
  assign t[45] = t[73] ^ t[74];
  assign t[46] = ~(t[75] ^ t[76]);
  assign t[47] = t[77] ^ t[78];
  assign t[48] = t[79] ^ t[80];
  assign t[49] = ~(t[81] & t[82]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[83] ^ t[214];
  assign t[51] = ~(t[209]);
  assign t[52] = t[84] & t[83];
  assign t[53] = ~(t[85]);
  assign t[54] = ~(t[215]);
  assign t[55] = ~(t[86] & t[216]);
  assign t[56] = ~(t[87] ^ t[88]);
  assign t[57] = t[89] ^ t[90];
  assign t[58] = ~(t[45] ^ t[22]);
  assign t[59] = t[91];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = ~t[92];
  assign t[61] = ~(t[37] ^ t[93]);
  assign t[62] = t[79] ^ t[94];
  assign t[63] = t[66] ? t[95] : t[217];
  assign t[64] = t[96] ^ t[70];
  assign t[65] = t[97] & t[98];
  assign t[66] = ~(t[99]);
  assign t[67] = t[213] ^ t[100];
  assign t[68] = t[101] & t[102];
  assign t[69] = t[103] ^ t[41];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[104] & t[105];
  assign t[71] = t[106] ^ t[107];
  assign t[72] = t[108] ^ t[109];
  assign t[73] = ~t[110];
  assign t[74] = t[93] ^ t[38];
  assign t[75] = t[111] ^ t[20];
  assign t[76] = ~(t[112] ^ t[113]);
  assign t[77] = t[114] ^ t[106];
  assign t[78] = t[115] & t[116];
  assign t[79] = t[60] ^ t[73];
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = t[93] ^ t[117];
  assign t[81] = ~(t[84] | t[83]);
  assign t[82] = ~(t[118] | t[51]);
  assign t[83] = ~(t[218]);
  assign t[84] = ~(t[214]);
  assign t[85] = ~(t[15]);
  assign t[86] = ~(t[219]);
  assign t[87] = t[21] ^ t[119];
  assign t[88] = t[120] ^ t[121];
  assign t[89] = t[122] ^ t[123];
  assign t[8] = t[207] ^ t[16];
  assign t[90] = t[124] ^ t[125];
  assign t[91] = t[66] ? t[126] : t[220];
  assign t[92] = t[66] ? t[127] : t[221];
  assign t[93] = t[128] ^ t[129];
  assign t[94] = t[130];
  assign t[95] = t[217] ^ t[131];
  assign t[96] = t[132] & t[133];
  assign t[97] = ~(t[96] ^ t[134]);
  assign t[98] = t[69] ^ t[135];
  assign t[99] = ~(t[7]);
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind93(x, y);
 input [116:0] x;
 output y;

 wire [242:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[190] ^ t[135];
  assign t[101] = ~(t[67] ^ t[136]);
  assign t[102] = t[137] ^ t[138];
  assign t[103] = t[139] & t[140];
  assign t[104] = ~(t[103] ^ t[141]);
  assign t[105] = t[18] ^ t[142];
  assign t[106] = ~(t[143] & t[144]);
  assign t[107] = t[145] ^ t[209];
  assign t[108] = ~(t[201]);
  assign t[109] = t[146] & t[145];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[129] ? x[72] : x[71];
  assign t[111] = t[129] ? x[74] : x[73];
  assign t[112] = t[203] ^ t[147];
  assign t[113] = t[129] ? x[76] : x[75];
  assign t[114] = t[99] ^ t[120];
  assign t[115] = t[148] & t[138];
  assign t[116] = t[32] ^ t[53];
  assign t[117] = t[149] & t[150];
  assign t[118] = t[125] ^ t[151];
  assign t[119] = t[152] ^ t[87];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[197] ^ t[153];
  assign t[121] = t[136] ^ t[68];
  assign t[122] = t[204] ^ t[154];
  assign t[123] = t[205] ^ t[155];
  assign t[124] = t[156] ^ t[157];
  assign t[125] = t[84] ^ t[97];
  assign t[126] = t[26] ? t[158] : t[210];
  assign t[127] = ~(t[152] ^ t[41]);
  assign t[128] = t[22] ^ t[93];
  assign t[129] = ~(t[159]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[7] ? t[160] : t[211];
  assign t[131] = t[206] ^ t[161];
  assign t[132] = t[207] ^ t[162];
  assign t[133] = ~(t[14]);
  assign t[134] = t[208] ^ t[163];
  assign t[135] = t[133] ? t[164] : t[212];
  assign t[136] = t[165] ^ t[115];
  assign t[137] = t[100] ^ t[120];
  assign t[138] = t[191] ^ t[166];
  assign t[139] = ~(t[142]);
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = ~(t[32]);
  assign t[141] = t[45] ^ t[32];
  assign t[142] = t[35] ^ t[53];
  assign t[143] = ~(t[146] | t[145]);
  assign t[144] = ~(t[167] | t[108]);
  assign t[145] = ~(t[213]);
  assign t[146] = ~(t[209]);
  assign t[147] = t[129] ? x[90] : x[89];
  assign t[148] = ~(t[100]);
  assign t[149] = ~(t[116] ^ t[69]);
  assign t[14] = ~(t[26]);
  assign t[150] = t[45] ^ t[35];
  assign t[151] = t[124] ^ t[168];
  assign t[152] = t[130] ^ t[39];
  assign t[153] = t[133] ? t[169] : t[214];
  assign t[154] = t[170] ? x[95] : x[94];
  assign t[155] = t[170] ? x[97] : x[96];
  assign t[156] = t[171] & t[172];
  assign t[157] = t[173] & t[126];
  assign t[158] = t[210] ^ t[174];
  assign t[159] = ~(t[27]);
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[211] ^ t[175];
  assign t[161] = t[129] ? x[99] : x[98];
  assign t[162] = t[27] ? x[101] : x[100];
  assign t[163] = t[176] ? x[103] : x[102];
  assign t[164] = t[212] ^ t[177];
  assign t[165] = t[178] & t[179];
  assign t[166] = t[133] ? t[180] : t[215];
  assign t[167] = ~(t[195]);
  assign t[168] = t[181] & t[182];
  assign t[169] = t[214] ^ t[183];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = ~(t[159]);
  assign t[171] = ~(t[184]);
  assign t[172] = ~(t[83]);
  assign t[173] = ~(t[84]);
  assign t[174] = t[27] ? x[108] : x[107];
  assign t[175] = t[129] ? x[110] : x[109];
  assign t[176] = ~(t[159]);
  assign t[177] = t[176] ? x[112] : x[111];
  assign t[178] = ~(t[185]);
  assign t[179] = ~(t[99]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[215] ^ t[186];
  assign t[181] = ~(t[156] ^ t[187]);
  assign t[182] = t[188] ^ t[184];
  assign t[183] = t[176] ? x[114] : x[113];
  assign t[184] = t[126] ^ t[84];
  assign t[185] = t[138] ^ t[100];
  assign t[186] = t[176] ? x[116] : x[115];
  assign t[187] = t[125] ^ t[83];
  assign t[188] = t[83] ^ t[97];
  assign t[189] = t[216] ^ x[4];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[217] ^ x[9];
  assign t[191] = t[218] ^ x[12];
  assign t[192] = t[219] ^ x[15];
  assign t[193] = t[220] ^ x[18];
  assign t[194] = t[221] ^ x[21];
  assign t[195] = t[222] ^ x[24];
  assign t[196] = t[223] ^ x[27];
  assign t[197] = t[224] ^ x[30];
  assign t[198] = t[225] ^ x[33];
  assign t[199] = t[226] ^ x[36];
  assign t[19] = t[34] & t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[39];
  assign t[201] = t[228] ^ x[42];
  assign t[202] = t[229] ^ x[45];
  assign t[203] = t[230] ^ x[48];
  assign t[204] = t[231] ^ x[51];
  assign t[205] = t[232] ^ x[54];
  assign t[206] = t[233] ^ x[61];
  assign t[207] = t[234] ^ x[64];
  assign t[208] = t[235] ^ x[67];
  assign t[209] = t[236] ^ x[70];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[79];
  assign t[211] = t[238] ^ x[82];
  assign t[212] = t[239] ^ x[85];
  assign t[213] = t[240] ^ x[88];
  assign t[214] = t[241] ^ x[93];
  assign t[215] = t[242] ^ x[106];
  assign t[216] = (x[2] & x[3]);
  assign t[217] = (x[7] & x[8]);
  assign t[218] = (x[10] & x[11]);
  assign t[219] = (x[13] & x[14]);
  assign t[21] = ~(t[25] ^ t[38]);
  assign t[220] = (x[16] & x[17]);
  assign t[221] = (x[19] & x[20]);
  assign t[222] = (x[22] & x[23]);
  assign t[223] = (x[25] & x[26]);
  assign t[224] = (x[28] & x[29]);
  assign t[225] = (x[31] & x[32]);
  assign t[226] = (x[34] & x[35]);
  assign t[227] = (x[37] & x[38]);
  assign t[228] = (x[40] & x[41]);
  assign t[229] = (x[43] & x[44]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (x[46] & x[47]);
  assign t[231] = (x[49] & x[50]);
  assign t[232] = (x[52] & x[53]);
  assign t[233] = (x[59] & x[60]);
  assign t[234] = (x[62] & x[63]);
  assign t[235] = (x[65] & x[66]);
  assign t[236] = (x[68] & x[69]);
  assign t[237] = (x[77] & x[78]);
  assign t[238] = (x[80] & x[81]);
  assign t[239] = (x[83] & x[84]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (x[86] & x[87]);
  assign t[241] = (x[91] & x[92]);
  assign t[242] = (x[104] & x[105]);
  assign t[24] = ~(t[43] ^ t[44]);
  assign t[25] = t[45] ^ t[46];
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[190]);
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[192]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[51];
  assign t[33] = ~t[52];
  assign t[34] = ~(t[53]);
  assign t[35] = t[54];
  assign t[36] = ~(t[55] ^ t[56]);
  assign t[37] = t[57] ^ t[58];
  assign t[38] = t[40] ^ t[59];
  assign t[39] = t[7] ? t[60] : t[193];
  assign t[3] = t[7] ? t[8] : t[189];
  assign t[40] = t[7] ? t[61] : t[194];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] & t[65];
  assign t[43] = t[12] ^ t[66];
  assign t[44] = t[67] ^ t[68];
  assign t[45] = t[53] ^ t[33];
  assign t[46] = t[69] ^ t[70];
  assign t[47] = ~(t[71] & t[72]);
  assign t[48] = t[195] | t[73];
  assign t[49] = ~(t[196]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[74] & t[197]);
  assign t[51] = t[7] ? t[75] : t[198];
  assign t[52] = t[7] ? t[76] : t[199];
  assign t[53] = ~t[77];
  assign t[54] = t[26] ? t[78] : t[200];
  assign t[55] = t[79] ^ t[80];
  assign t[56] = ~(t[81] ^ t[82]);
  assign t[57] = t[83] ^ t[84];
  assign t[58] = t[85] & t[86];
  assign t[59] = t[41] ^ t[87];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[193] ^ t[88];
  assign t[61] = t[194] ^ t[89];
  assign t[62] = t[90] & t[91];
  assign t[63] = t[92] & t[93];
  assign t[64] = ~(t[62] ^ t[94]);
  assign t[65] = t[95] ^ t[96];
  assign t[66] = t[97] ^ t[98];
  assign t[67] = t[99] ^ t[100];
  assign t[68] = t[101] & t[102];
  assign t[69] = t[103] ^ t[19];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[104] & t[105];
  assign t[71] = ~(t[73] & t[106]);
  assign t[72] = ~(t[201] ^ t[107]);
  assign t[73] = ~(t[108] & t[109]);
  assign t[74] = ~(t[202]);
  assign t[75] = t[198] ^ t[110];
  assign t[76] = t[199] ^ t[111];
  assign t[77] = t[7] ? t[112] : t[203];
  assign t[78] = t[200] ^ t[113];
  assign t[79] = t[114] ^ t[115];
  assign t[7] = ~(t[14]);
  assign t[80] = t[116] ^ t[117];
  assign t[81] = t[118] ^ t[119];
  assign t[82] = t[120] ^ t[121];
  assign t[83] = t[26] ? t[122] : t[204];
  assign t[84] = t[26] ? t[123] : t[205];
  assign t[85] = ~(t[57] ^ t[124]);
  assign t[86] = t[125] ^ t[126];
  assign t[87] = t[127] & t[128];
  assign t[88] = t[129] ? x[56] : x[55];
  assign t[89] = t[129] ? x[58] : x[57];
  assign t[8] = t[189] ^ t[15];
  assign t[90] = ~(t[96]);
  assign t[91] = ~(t[130]);
  assign t[92] = ~(t[39]);
  assign t[93] = t[7] ? t[131] : t[206];
  assign t[94] = t[22] ^ t[130];
  assign t[95] = t[130] ^ t[40];
  assign t[96] = t[93] ^ t[39];
  assign t[97] = t[26] ? t[132] : t[207];
  assign t[98] = t[124] ^ t[58];
  assign t[99] = t[133] ? t[134] : t[208];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind94(x, y);
 input [116:0] x;
 output y;

 wire [249:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[7] ? t[136] : t[213];
  assign t[101] = t[87] ^ t[22];
  assign t[102] = t[137] ? x[61] : x[60];
  assign t[103] = t[137] ? x[63] : x[62];
  assign t[104] = t[138] & t[139];
  assign t[105] = t[140] & t[71];
  assign t[106] = t[7] ? t[141] : t[214];
  assign t[107] = t[206] ^ t[142];
  assign t[108] = ~(t[143] & t[144]);
  assign t[109] = t[145] ^ t[215];
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = ~(t[207]);
  assign t[111] = t[146] & t[145];
  assign t[112] = t[147] ^ t[64];
  assign t[113] = ~(t[148] ^ t[38]);
  assign t[114] = t[149] ^ t[150];
  assign t[115] = t[42] ^ t[106];
  assign t[116] = t[69] ^ t[25];
  assign t[117] = t[209] ^ t[151];
  assign t[118] = t[152] ? t[153] : t[216];
  assign t[119] = t[200] ^ t[154];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[26] ? t[155] : t[217];
  assign t[121] = t[156] & t[157];
  assign t[122] = t[158] ^ t[53];
  assign t[123] = t[159] & t[160];
  assign t[124] = t[210] ^ t[161];
  assign t[125] = t[211] ^ t[162];
  assign t[126] = t[26] ? t[163] : t[218];
  assign t[127] = t[164];
  assign t[128] = t[26] ? t[165] : t[219];
  assign t[129] = t[166] & t[167];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[212] ^ t[168];
  assign t[131] = t[169] & t[170];
  assign t[132] = ~(t[171] ^ t[94]);
  assign t[133] = t[149] ^ t[90];
  assign t[134] = ~(t[27]);
  assign t[135] = t[100] ^ t[87];
  assign t[136] = t[213] ^ t[172];
  assign t[137] = ~(t[134]);
  assign t[138] = ~(t[173]);
  assign t[139] = ~(t[42]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[43]);
  assign t[141] = t[214] ^ t[174];
  assign t[142] = t[137] ? x[83] : x[82];
  assign t[143] = ~(t[146] | t[145]);
  assign t[144] = ~(t[175] | t[110]);
  assign t[145] = ~(t[220]);
  assign t[146] = ~(t[215]);
  assign t[147] = t[86] ^ t[22];
  assign t[148] = t[176] ^ t[123];
  assign t[149] = t[127] ^ t[60];
  assign t[14] = ~(t[26]);
  assign t[150] = t[94] ^ t[177];
  assign t[151] = t[96] ? x[88] : x[87];
  assign t[152] = ~(t[14]);
  assign t[153] = t[216] ^ t[178];
  assign t[154] = t[26] ? t[179] : t[221];
  assign t[155] = t[217] ^ t[180];
  assign t[156] = ~(t[104] ^ t[181]);
  assign t[157] = t[115] ^ t[173];
  assign t[158] = t[182] & t[183];
  assign t[159] = ~(t[176] ^ t[122]);
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[91] ^ t[83];
  assign t[161] = t[96] ? x[93] : x[92];
  assign t[162] = t[96] ? x[95] : x[94];
  assign t[163] = t[218] ^ t[184];
  assign t[164] = t[26] ? t[185] : t[222];
  assign t[165] = t[219] ^ t[186];
  assign t[166] = ~(t[158] ^ t[187]);
  assign t[167] = t[52] ^ t[188];
  assign t[168] = t[27] ? x[100] : x[99];
  assign t[169] = ~(t[189]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = ~(t[88]);
  assign t[171] = t[88] ^ t[127];
  assign t[172] = t[96] ? x[102] : x[101];
  assign t[173] = t[71] ^ t[43];
  assign t[174] = t[137] ? x[104] : x[103];
  assign t[175] = ~(t[203]);
  assign t[176] = t[80] ^ t[119];
  assign t[177] = t[190] & t[191];
  assign t[178] = t[192] ? x[106] : x[105];
  assign t[179] = t[221] ^ t[193];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[27] ? x[108] : x[107];
  assign t[181] = t[70] ^ t[42];
  assign t[182] = ~(t[188]);
  assign t[183] = ~(t[80]);
  assign t[184] = t[27] ? x[110] : x[109];
  assign t[185] = t[222] ^ t[194];
  assign t[186] = t[192] ? x[112] : x[111];
  assign t[187] = t[91] ^ t[80];
  assign t[188] = t[83] ^ t[119];
  assign t[189] = t[90] ^ t[127];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = ~(t[131] ^ t[195]);
  assign t[191] = t[57] ^ t[189];
  assign t[192] = ~(t[134]);
  assign t[193] = t[96] ? x[114] : x[113];
  assign t[194] = t[192] ? x[116] : x[115];
  assign t[195] = t[149] ^ t[88];
  assign t[196] = t[223] ^ x[4];
  assign t[197] = t[224] ^ x[9];
  assign t[198] = t[225] ^ x[12];
  assign t[199] = t[226] ^ x[15];
  assign t[19] = ~(t[34] ^ t[35]);
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[18];
  assign t[201] = t[228] ^ x[21];
  assign t[202] = t[229] ^ x[24];
  assign t[203] = t[230] ^ x[27];
  assign t[204] = t[231] ^ x[30];
  assign t[205] = t[232] ^ x[33];
  assign t[206] = t[233] ^ x[38];
  assign t[207] = t[234] ^ x[41];
  assign t[208] = t[235] ^ x[44];
  assign t[209] = t[236] ^ x[47];
  assign t[20] = t[36] ^ t[35];
  assign t[210] = t[237] ^ x[50];
  assign t[211] = t[238] ^ x[53];
  assign t[212] = t[239] ^ x[56];
  assign t[213] = t[240] ^ x[59];
  assign t[214] = t[241] ^ x[66];
  assign t[215] = t[242] ^ x[69];
  assign t[216] = t[243] ^ x[72];
  assign t[217] = t[244] ^ x[75];
  assign t[218] = t[245] ^ x[78];
  assign t[219] = t[246] ^ x[81];
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = t[247] ^ x[86];
  assign t[221] = t[248] ^ x[91];
  assign t[222] = t[249] ^ x[98];
  assign t[223] = (x[2] & x[3]);
  assign t[224] = (x[7] & x[8]);
  assign t[225] = (x[10] & x[11]);
  assign t[226] = (x[13] & x[14]);
  assign t[227] = (x[16] & x[17]);
  assign t[228] = (x[19] & x[20]);
  assign t[229] = (x[22] & x[23]);
  assign t[22] = t[7] ? t[39] : t[197];
  assign t[230] = (x[25] & x[26]);
  assign t[231] = (x[28] & x[29]);
  assign t[232] = (x[31] & x[32]);
  assign t[233] = (x[36] & x[37]);
  assign t[234] = (x[39] & x[40]);
  assign t[235] = (x[42] & x[43]);
  assign t[236] = (x[45] & x[46]);
  assign t[237] = (x[48] & x[49]);
  assign t[238] = (x[51] & x[52]);
  assign t[239] = (x[54] & x[55]);
  assign t[23] = t[40] ^ t[41];
  assign t[240] = (x[57] & x[58]);
  assign t[241] = (x[64] & x[65]);
  assign t[242] = (x[67] & x[68]);
  assign t[243] = (x[70] & x[71]);
  assign t[244] = (x[73] & x[74]);
  assign t[245] = (x[76] & x[77]);
  assign t[246] = (x[79] & x[80]);
  assign t[247] = (x[84] & x[85]);
  assign t[248] = (x[89] & x[90]);
  assign t[249] = (x[96] & x[97]);
  assign t[24] = t[42] ^ t[43];
  assign t[25] = t[44] & t[45];
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[198]);
  assign t[29] = ~(t[199]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[200]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = ~(t[50] ^ t[51]);
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] ^ t[41];
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ t[13];
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[197] ^ t[62];
  assign t[3] = t[7] ? t[8] : t[196];
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65] & t[66];
  assign t[42] = t[7] ? t[67] : t[201];
  assign t[43] = t[7] ? t[68] : t[202];
  assign t[44] = ~(t[24] ^ t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[203] | t[74];
  assign t[48] = ~(t[204]);
  assign t[49] = ~(t[75] & t[205]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[76] ^ t[77];
  assign t[51] = ~(t[78] ^ t[79]);
  assign t[52] = t[80] ^ t[81];
  assign t[53] = t[82] & t[83];
  assign t[54] = t[70] ^ t[84];
  assign t[55] = t[81] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ^ t[60];
  assign t[58] = t[89] & t[90];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[93];
  assign t[61] = t[94] ^ t[95];
  assign t[62] = t[96] ? x[35] : x[34];
  assign t[63] = t[97] & t[98];
  assign t[64] = t[99] & t[100];
  assign t[65] = ~(t[56] ^ t[40]);
  assign t[66] = t[101] ^ t[100];
  assign t[67] = t[201] ^ t[102];
  assign t[68] = t[202] ^ t[103];
  assign t[69] = t[104] ^ t[105];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[43] ^ t[106];
  assign t[71] = t[7] ? t[107] : t[206];
  assign t[72] = ~(t[74] & t[108]);
  assign t[73] = ~(t[207] ^ t[109]);
  assign t[74] = ~(t[110] & t[111]);
  assign t[75] = ~(t[208]);
  assign t[76] = t[12] ^ t[112];
  assign t[77] = ~(t[113] ^ t[114]);
  assign t[78] = t[115] ^ t[105];
  assign t[79] = t[106] ^ t[116];
  assign t[7] = ~(t[14]);
  assign t[80] = t[26] ? t[117] : t[209];
  assign t[81] = t[204] ^ t[118];
  assign t[82] = ~(t[119]);
  assign t[83] = t[208] ^ t[120];
  assign t[84] = t[69] ^ t[121];
  assign t[85] = t[122] ^ t[123];
  assign t[86] = t[7] ? t[124] : t[210];
  assign t[87] = t[7] ? t[125] : t[211];
  assign t[88] = ~t[126];
  assign t[89] = ~(t[127]);
  assign t[8] = t[196] ^ t[15];
  assign t[90] = t[128];
  assign t[91] = t[119] ^ t[81];
  assign t[92] = t[122] ^ t[129];
  assign t[93] = t[26] ? t[130] : t[212];
  assign t[94] = t[131] ^ t[58];
  assign t[95] = t[132] & t[133];
  assign t[96] = ~(t[134]);
  assign t[97] = ~(t[135]);
  assign t[98] = ~(t[86]);
  assign t[99] = ~(t[87]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind95(x, y);
 input [116:0] x;
 output y;

 wire [249:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[205] ^ t[135];
  assign t[101] = t[136] & t[137];
  assign t[102] = t[138] & t[123];
  assign t[103] = t[139] & t[140];
  assign t[104] = t[7] ? t[141] : t[212];
  assign t[105] = t[7] ? t[142] : t[213];
  assign t[106] = ~(t[68] ^ t[143]);
  assign t[107] = t[144] ^ t[145];
  assign t[108] = t[144] ^ t[146];
  assign t[109] = t[147] ^ t[61];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[88] ^ t[40];
  assign t[111] = t[34] ^ t[148];
  assign t[112] = t[7] ? t[149] : t[214];
  assign t[113] = t[143] ^ t[69];
  assign t[114] = ~(t[150] & t[151]);
  assign t[115] = t[152] ^ t[215];
  assign t[116] = ~(t[206]);
  assign t[117] = t[153] & t[152];
  assign t[118] = ~(t[154]);
  assign t[119] = t[7] ? t[155] : t[216];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[208] ^ t[156];
  assign t[121] = t[209] ^ t[157];
  assign t[122] = t[26] ? t[158] : t[217];
  assign t[123] = t[207] ^ t[159];
  assign t[124] = t[210] ^ t[160];
  assign t[125] = ~(t[109] ^ t[62]);
  assign t[126] = t[38] ^ t[131];
  assign t[127] = t[211] ^ t[161];
  assign t[128] = ~(t[134]);
  assign t[129] = ~(t[147]);
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = ~(t[61]);
  assign t[131] = t[162];
  assign t[132] = t[38] ^ t[147];
  assign t[133] = t[147] ^ t[59];
  assign t[134] = t[131] ^ t[61];
  assign t[135] = t[163] ? x[75] : x[74];
  assign t[136] = ~(t[164]);
  assign t[137] = ~(t[88]);
  assign t[138] = ~(t[89]);
  assign t[139] = ~(t[101] ^ t[165]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[110] ^ t[164];
  assign t[141] = t[212] ^ t[166];
  assign t[142] = t[213] ^ t[167];
  assign t[143] = t[168] ^ t[169];
  assign t[144] = t[105] ^ t[112];
  assign t[145] = t[7] ? t[170] : t[218];
  assign t[146] = t[143] ^ t[171];
  assign t[147] = ~t[172];
  assign t[148] = t[173] & t[174];
  assign t[149] = t[214] ^ t[175];
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[153] | t[152]);
  assign t[151] = ~(t[176] | t[116]);
  assign t[152] = ~(t[219]);
  assign t[153] = ~(t[215]);
  assign t[154] = ~(t[27]);
  assign t[155] = t[216] ^ t[177];
  assign t[156] = t[118] ? x[83] : x[82];
  assign t[157] = t[118] ? x[85] : x[84];
  assign t[158] = t[217] ^ t[178];
  assign t[159] = t[26] ? t[179] : t[220];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[27] ? x[90] : x[89];
  assign t[161] = t[163] ? x[92] : x[91];
  assign t[162] = t[26] ? t[180] : t[221];
  assign t[163] = ~(t[154]);
  assign t[164] = t[123] ^ t[89];
  assign t[165] = t[66] ^ t[88];
  assign t[166] = t[181] ? x[97] : x[96];
  assign t[167] = t[181] ? x[99] : x[98];
  assign t[168] = t[182] & t[183];
  assign t[169] = t[184] & t[145];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[218] ^ t[185];
  assign t[171] = t[186] & t[187];
  assign t[172] = t[26] ? t[188] : t[222];
  assign t[173] = ~(t[189] ^ t[34]);
  assign t[174] = t[18] ^ t[84];
  assign t[175] = t[181] ? x[104] : x[103];
  assign t[176] = ~(t[203]);
  assign t[177] = t[118] ? x[106] : x[105];
  assign t[178] = t[118] ? x[108] : x[107];
  assign t[179] = t[220] ^ t[190];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[221] ^ t[191];
  assign t[181] = ~(t[154]);
  assign t[182] = ~(t[192]);
  assign t[183] = ~(t[104]);
  assign t[184] = ~(t[105]);
  assign t[185] = t[181] ? x[110] : x[109];
  assign t[186] = ~(t[168] ^ t[193]);
  assign t[187] = t[194] ^ t[192];
  assign t[188] = t[222] ^ t[195];
  assign t[189] = t[119] ^ t[32];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[27] ? x[112] : x[111];
  assign t[191] = t[163] ? x[114] : x[113];
  assign t[192] = t[145] ^ t[105];
  assign t[193] = t[144] ^ t[104];
  assign t[194] = t[104] ^ t[112];
  assign t[195] = t[27] ? x[116] : x[115];
  assign t[196] = t[223] ^ x[4];
  assign t[197] = t[224] ^ x[9];
  assign t[198] = t[225] ^ x[12];
  assign t[199] = t[226] ^ x[15];
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[18];
  assign t[201] = t[228] ^ x[21];
  assign t[202] = t[229] ^ x[24];
  assign t[203] = t[230] ^ x[27];
  assign t[204] = t[231] ^ x[30];
  assign t[205] = t[232] ^ x[33];
  assign t[206] = t[233] ^ x[36];
  assign t[207] = t[234] ^ x[39];
  assign t[208] = t[235] ^ x[46];
  assign t[209] = t[236] ^ x[49];
  assign t[20] = ~(t[36] ^ t[37]);
  assign t[210] = t[237] ^ x[52];
  assign t[211] = t[238] ^ x[55];
  assign t[212] = t[239] ^ x[58];
  assign t[213] = t[240] ^ x[61];
  assign t[214] = t[241] ^ x[64];
  assign t[215] = t[242] ^ x[67];
  assign t[216] = t[243] ^ x[70];
  assign t[217] = t[244] ^ x[73];
  assign t[218] = t[245] ^ x[78];
  assign t[219] = t[246] ^ x[81];
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[247] ^ x[88];
  assign t[221] = t[248] ^ x[95];
  assign t[222] = t[249] ^ x[102];
  assign t[223] = (x[2] & x[3]);
  assign t[224] = (x[7] & x[8]);
  assign t[225] = (x[10] & x[11]);
  assign t[226] = (x[13] & x[14]);
  assign t[227] = (x[16] & x[17]);
  assign t[228] = (x[19] & x[20]);
  assign t[229] = (x[22] & x[23]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (x[25] & x[26]);
  assign t[231] = (x[28] & x[29]);
  assign t[232] = (x[31] & x[32]);
  assign t[233] = (x[34] & x[35]);
  assign t[234] = (x[37] & x[38]);
  assign t[235] = (x[44] & x[45]);
  assign t[236] = (x[47] & x[48]);
  assign t[237] = (x[50] & x[51]);
  assign t[238] = (x[53] & x[54]);
  assign t[239] = (x[56] & x[57]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (x[59] & x[60]);
  assign t[241] = (x[62] & x[63]);
  assign t[242] = (x[65] & x[66]);
  assign t[243] = (x[68] & x[69]);
  assign t[244] = (x[71] & x[72]);
  assign t[245] = (x[76] & x[77]);
  assign t[246] = (x[79] & x[80]);
  assign t[247] = (x[86] & x[87]);
  assign t[248] = (x[93] & x[94]);
  assign t[249] = (x[100] & x[101]);
  assign t[24] = ~(t[44] ^ t[10]);
  assign t[25] = ~(t[45] ^ t[46]);
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[197]);
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[199]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[7] ? t[51] : t[200];
  assign t[33] = t[7] ? t[52] : t[201];
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[55] & t[56];
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[61] ^ t[59];
  assign t[39] = t[62] ^ t[63];
  assign t[3] = t[7] ? t[8] : t[196];
  assign t[40] = t[202] ^ t[64];
  assign t[41] = t[65] ^ t[58];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = ~(t[70] ^ t[71]);
  assign t[45] = t[21] ^ t[72];
  assign t[46] = ~(t[73] ^ t[74]);
  assign t[47] = ~(t[75] & t[76]);
  assign t[48] = t[203] | t[77];
  assign t[49] = ~(t[202]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[78] & t[204]);
  assign t[51] = t[200] ^ t[79];
  assign t[52] = t[201] ^ t[80];
  assign t[53] = t[81] & t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = ~(t[53] ^ t[85]);
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ^ t[89];
  assign t[58] = t[90] & t[91];
  assign t[59] = t[92];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[62] ^ t[93];
  assign t[61] = t[94];
  assign t[62] = t[95] ^ t[96];
  assign t[63] = t[97] & t[98];
  assign t[64] = t[99] ? t[100] : t[205];
  assign t[65] = t[101] ^ t[102];
  assign t[66] = t[89] ^ t[40];
  assign t[67] = t[65] ^ t[103];
  assign t[68] = t[104] ^ t[105];
  assign t[69] = t[106] & t[107];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[108] ^ t[22];
  assign t[71] = t[109] ^ t[93];
  assign t[72] = t[110] ^ t[102];
  assign t[73] = t[33] ^ t[111];
  assign t[74] = t[112] ^ t[113];
  assign t[75] = ~(t[77] & t[114]);
  assign t[76] = ~(t[206] ^ t[115]);
  assign t[77] = ~(t[116] & t[117]);
  assign t[78] = ~(t[207]);
  assign t[79] = t[118] ? x[41] : x[40];
  assign t[7] = ~(t[14]);
  assign t[80] = t[118] ? x[43] : x[42];
  assign t[81] = ~(t[87]);
  assign t[82] = ~(t[119]);
  assign t[83] = ~(t[32]);
  assign t[84] = t[7] ? t[120] : t[208];
  assign t[85] = t[18] ^ t[119];
  assign t[86] = t[119] ^ t[33];
  assign t[87] = t[84] ^ t[32];
  assign t[88] = t[26] ? t[121] : t[209];
  assign t[89] = t[199] ^ t[122];
  assign t[8] = t[196] ^ t[15];
  assign t[90] = ~(t[57] ^ t[65]);
  assign t[91] = t[66] ^ t[123];
  assign t[92] = t[26] ? t[124] : t[210];
  assign t[93] = t[125] & t[126];
  assign t[94] = t[26] ? t[127] : t[211];
  assign t[95] = t[128] & t[129];
  assign t[96] = t[130] & t[131];
  assign t[97] = ~(t[95] ^ t[132]);
  assign t[98] = t[133] ^ t[134];
  assign t[99] = ~(t[14]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind96(x, y);
 input [116:0] x;
 output y;

 wire [260:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[137] ^ t[120];
  assign t[101] = t[138] & t[139];
  assign t[102] = t[218] ^ t[140];
  assign t[103] = t[141] ^ t[142];
  assign t[104] = t[41] ^ t[143];
  assign t[105] = t[144] ^ t[145];
  assign t[106] = t[26] ? t[146] : t[224];
  assign t[107] = ~(t[71] ^ t[100]);
  assign t[108] = t[65] ^ t[147];
  assign t[109] = t[148] & t[149];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = ~(t[150] & t[151]);
  assign t[111] = t[152] ^ t[225];
  assign t[112] = ~(t[219]);
  assign t[113] = t[153] & t[152];
  assign t[114] = t[99] ^ t[154];
  assign t[115] = t[155] ^ t[156];
  assign t[116] = t[157] & t[158];
  assign t[117] = t[156] ^ t[144];
  assign t[118] = t[159] ^ t[160];
  assign t[119] = t[106] ^ t[99];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[161] & t[147];
  assign t[121] = t[27] ? x[64] : x[63];
  assign t[122] = t[27] ? x[66] : x[65];
  assign t[123] = t[162] & t[163];
  assign t[124] = t[164] & t[87];
  assign t[125] = t[221] ^ t[165];
  assign t[126] = t[131] ? x[68] : x[67];
  assign t[127] = ~(t[130]);
  assign t[128] = ~(t[95]);
  assign t[129] = t[36] ^ t[95];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[97] ^ t[58];
  assign t[131] = ~(t[48]);
  assign t[132] = t[95] ^ t[58];
  assign t[133] = t[222] ^ t[166];
  assign t[134] = t[223] ^ t[167];
  assign t[135] = t[26] ? t[168] : t[226];
  assign t[136] = t[169] ? t[170] : t[227];
  assign t[137] = t[171] & t[172];
  assign t[138] = ~(t[137] ^ t[173]);
  assign t[139] = t[119] ^ t[174];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[27] ? x[76] : x[75];
  assign t[141] = t[155] ^ t[144];
  assign t[142] = t[175] & t[176];
  assign t[143] = t[132] ^ t[62];
  assign t[144] = t[177];
  assign t[145] = t[159] ^ t[116];
  assign t[146] = t[224] ^ t[178];
  assign t[147] = t[220] ^ t[179];
  assign t[148] = ~(t[123] ^ t[180]);
  assign t[149] = t[181] ^ t[182];
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[153] | t[152]);
  assign t[151] = ~(t[183] | t[112]);
  assign t[152] = ~(t[228]);
  assign t[153] = ~(t[225]);
  assign t[154] = t[100] ^ t[72];
  assign t[155] = ~t[184];
  assign t[156] = t[185];
  assign t[157] = ~(t[115] ^ t[159]);
  assign t[158] = t[117] ^ t[176];
  assign t[159] = t[186] ^ t[142];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[187] & t[188];
  assign t[161] = ~(t[98]);
  assign t[162] = ~(t[182]);
  assign t[163] = ~(t[54]);
  assign t[164] = ~(t[55]);
  assign t[165] = t[27] ? x[81] : x[80];
  assign t[166] = t[131] ? x[83] : x[82];
  assign t[167] = t[131] ? x[85] : x[84];
  assign t[168] = t[226] ^ t[189];
  assign t[169] = ~(t[14]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[227] ^ t[190];
  assign t[171] = ~(t[174]);
  assign t[172] = ~(t[106]);
  assign t[173] = t[65] ^ t[106];
  assign t[174] = t[147] ^ t[98];
  assign t[175] = ~(t[156]);
  assign t[176] = t[191];
  assign t[177] = t[26] ? t[192] : t[229];
  assign t[178] = t[27] ? x[90] : x[89];
  assign t[179] = t[26] ? t[193] : t[230];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[73] ^ t[54];
  assign t[181] = t[54] ^ t[67];
  assign t[182] = t[87] ^ t[55];
  assign t[183] = ~(t[212]);
  assign t[184] = t[26] ? t[194] : t[231];
  assign t[185] = t[26] ? t[195] : t[232];
  assign t[186] = t[196] & t[197];
  assign t[187] = ~(t[186] ^ t[198]);
  assign t[188] = t[141] ^ t[199];
  assign t[189] = t[27] ? x[101] : x[100];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[200] ? x[103] : x[102];
  assign t[191] = t[26] ? t[201] : t[233];
  assign t[192] = t[229] ^ t[202];
  assign t[193] = t[230] ^ t[203];
  assign t[194] = t[231] ^ t[204];
  assign t[195] = t[232] ^ t[205];
  assign t[196] = ~(t[199]);
  assign t[197] = ~(t[155]);
  assign t[198] = t[117] ^ t[155];
  assign t[199] = t[176] ^ t[156];
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = ~(t[48]);
  assign t[201] = t[233] ^ t[206];
  assign t[202] = t[78] ? x[108] : x[107];
  assign t[203] = t[78] ? x[110] : x[109];
  assign t[204] = t[78] ? x[112] : x[111];
  assign t[205] = t[200] ? x[114] : x[113];
  assign t[206] = t[200] ? x[116] : x[115];
  assign t[207] = t[234] ^ x[4];
  assign t[208] = t[235] ^ x[9];
  assign t[209] = t[236] ^ x[12];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[15];
  assign t[211] = t[238] ^ x[18];
  assign t[212] = t[239] ^ x[21];
  assign t[213] = t[240] ^ x[24];
  assign t[214] = t[241] ^ x[27];
  assign t[215] = t[242] ^ x[30];
  assign t[216] = t[243] ^ x[33];
  assign t[217] = t[244] ^ x[36];
  assign t[218] = t[245] ^ x[39];
  assign t[219] = t[246] ^ x[42];
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[247] ^ x[45];
  assign t[221] = t[248] ^ x[48];
  assign t[222] = t[249] ^ x[53];
  assign t[223] = t[250] ^ x[56];
  assign t[224] = t[251] ^ x[59];
  assign t[225] = t[252] ^ x[62];
  assign t[226] = t[253] ^ x[71];
  assign t[227] = t[254] ^ x[74];
  assign t[228] = t[255] ^ x[79];
  assign t[229] = t[256] ^ x[88];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[93];
  assign t[231] = t[258] ^ x[96];
  assign t[232] = t[259] ^ x[99];
  assign t[233] = t[260] ^ x[106];
  assign t[234] = (x[2] & x[3]);
  assign t[235] = (x[7] & x[8]);
  assign t[236] = (x[10] & x[11]);
  assign t[237] = (x[13] & x[14]);
  assign t[238] = (x[16] & x[17]);
  assign t[239] = (x[19] & x[20]);
  assign t[23] = ~(t[32] ^ t[42]);
  assign t[240] = (x[22] & x[23]);
  assign t[241] = (x[25] & x[26]);
  assign t[242] = (x[28] & x[29]);
  assign t[243] = (x[31] & x[32]);
  assign t[244] = (x[34] & x[35]);
  assign t[245] = (x[37] & x[38]);
  assign t[246] = (x[40] & x[41]);
  assign t[247] = (x[43] & x[44]);
  assign t[248] = (x[46] & x[47]);
  assign t[249] = (x[51] & x[52]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (x[54] & x[55]);
  assign t[251] = (x[57] & x[58]);
  assign t[252] = (x[60] & x[61]);
  assign t[253] = (x[69] & x[70]);
  assign t[254] = (x[72] & x[73]);
  assign t[255] = (x[77] & x[78]);
  assign t[256] = (x[86] & x[87]);
  assign t[257] = (x[91] & x[92]);
  assign t[258] = (x[94] & x[95]);
  assign t[259] = (x[97] & x[98]);
  assign t[25] = ~(t[45] ^ t[21]);
  assign t[260] = (x[104] & x[105]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[208]);
  assign t[29] = ~(t[209]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[210]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = ~(t[51] ^ t[45]);
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] & t[57];
  assign t[36] = t[58] ^ t[38];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[7] ? t[61] : t[211];
  assign t[39] = t[59] ^ t[62];
  assign t[3] = t[7] ? t[8] : t[207];
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] ^ t[68];
  assign t[43] = ~(t[69] ^ t[70]);
  assign t[44] = t[71] ^ t[72];
  assign t[45] = t[73] ^ t[74];
  assign t[46] = ~(t[75] & t[76]);
  assign t[47] = t[212] | t[77];
  assign t[48] = ~(t[78]);
  assign t[49] = ~(t[213]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[79] & t[214]);
  assign t[51] = ~(t[80] ^ t[81]);
  assign t[52] = t[82] ^ t[83];
  assign t[53] = ~(t[42] ^ t[21]);
  assign t[54] = t[7] ? t[84] : t[215];
  assign t[55] = t[7] ? t[85] : t[216];
  assign t[56] = ~(t[34] ^ t[86]);
  assign t[57] = t[73] ^ t[87];
  assign t[58] = t[7] ? t[88] : t[217];
  assign t[59] = t[89] ^ t[64];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[90] & t[91];
  assign t[61] = t[211] ^ t[92];
  assign t[62] = t[93] & t[94];
  assign t[63] = t[95] ^ t[38];
  assign t[64] = t[96] & t[97];
  assign t[65] = t[98] ^ t[99];
  assign t[66] = t[100] ^ t[101];
  assign t[67] = t[7] ? t[102] : t[218];
  assign t[68] = t[86] ^ t[35];
  assign t[69] = t[103] ^ t[19];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[104] ^ t[105]);
  assign t[71] = t[106] ^ t[98];
  assign t[72] = t[107] & t[108];
  assign t[73] = t[55] ^ t[67];
  assign t[74] = t[86] ^ t[109];
  assign t[75] = ~(t[77] & t[110]);
  assign t[76] = ~(t[219] ^ t[111]);
  assign t[77] = ~(t[112] & t[113]);
  assign t[78] = ~(t[47]);
  assign t[79] = ~(t[220]);
  assign t[7] = ~(t[14]);
  assign t[80] = t[20] ^ t[114];
  assign t[81] = t[115] ^ t[116];
  assign t[82] = t[117] ^ t[118];
  assign t[83] = t[119] ^ t[120];
  assign t[84] = t[215] ^ t[121];
  assign t[85] = t[216] ^ t[122];
  assign t[86] = t[123] ^ t[124];
  assign t[87] = t[7] ? t[125] : t[221];
  assign t[88] = t[217] ^ t[126];
  assign t[89] = t[127] & t[128];
  assign t[8] = t[207] ^ t[15];
  assign t[90] = ~(t[89] ^ t[129]);
  assign t[91] = t[63] ^ t[130];
  assign t[92] = t[131] ? x[50] : x[49];
  assign t[93] = ~(t[132] ^ t[59]);
  assign t[94] = t[36] ^ t[97];
  assign t[95] = t[7] ? t[133] : t[222];
  assign t[96] = ~(t[58]);
  assign t[97] = t[7] ? t[134] : t[223];
  assign t[98] = t[210] ^ t[135];
  assign t[99] = t[213] ^ t[136];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind97(x, y);
 input [116:0] x;
 output y;

 wire [242:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[132];
  assign t[101] = ~(t[67] ^ t[133]);
  assign t[102] = t[134] ^ t[135];
  assign t[103] = t[136] & t[137];
  assign t[104] = ~(t[103] ^ t[138]);
  assign t[105] = t[18] ^ t[139];
  assign t[106] = ~(t[140] & t[141]);
  assign t[107] = t[142] ^ t[206];
  assign t[108] = ~(t[202]);
  assign t[109] = t[143] & t[142];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = ~(t[144]);
  assign t[111] = t[110] ? x[69] : x[68];
  assign t[112] = t[99] ^ t[118];
  assign t[113] = t[145] & t[135];
  assign t[114] = t[32] ^ t[53];
  assign t[115] = t[146] & t[147];
  assign t[116] = t[123] ^ t[148];
  assign t[117] = t[149] ^ t[87];
  assign t[118] = t[150];
  assign t[119] = t[133] ^ t[68];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[204] ^ t[151];
  assign t[121] = t[26] ? t[152] : t[207];
  assign t[122] = t[153] ^ t[154];
  assign t[123] = t[84] ^ t[97];
  assign t[124] = t[203] ^ t[155];
  assign t[125] = ~(t[149] ^ t[41]);
  assign t[126] = t[22] ^ t[93];
  assign t[127] = ~(t[144]);
  assign t[128] = t[7] ? t[156] : t[208];
  assign t[129] = t[205] ^ t[157];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ? t[159] : t[209];
  assign t[131] = t[26] ? t[160] : t[210];
  assign t[132] = t[26] ? t[161] : t[211];
  assign t[133] = t[162] ^ t[113];
  assign t[134] = t[100] ^ t[118];
  assign t[135] = t[163];
  assign t[136] = ~(t[139]);
  assign t[137] = ~(t[32]);
  assign t[138] = t[45] ^ t[32];
  assign t[139] = t[35] ^ t[53];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = ~(t[143] | t[142]);
  assign t[141] = ~(t[164] | t[108]);
  assign t[142] = ~(t[212]);
  assign t[143] = ~(t[206]);
  assign t[144] = ~(t[27]);
  assign t[145] = ~(t[100]);
  assign t[146] = ~(t[114] ^ t[69]);
  assign t[147] = t[45] ^ t[35];
  assign t[148] = t[122] ^ t[165];
  assign t[149] = t[128] ^ t[39];
  assign t[14] = ~(t[26]);
  assign t[150] = t[26] ? t[166] : t[213];
  assign t[151] = t[110] ? x[92] : x[91];
  assign t[152] = t[207] ^ t[167];
  assign t[153] = t[168] & t[169];
  assign t[154] = t[170] & t[124];
  assign t[155] = t[26] ? t[171] : t[214];
  assign t[156] = t[208] ^ t[172];
  assign t[157] = t[127] ? x[97] : x[96];
  assign t[158] = ~(t[14]);
  assign t[159] = t[209] ^ t[173];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[210] ^ t[174];
  assign t[161] = t[211] ^ t[175];
  assign t[162] = t[176] & t[177];
  assign t[163] = t[26] ? t[178] : t[215];
  assign t[164] = ~(t[198]);
  assign t[165] = t[179] & t[180];
  assign t[166] = t[213] ^ t[181];
  assign t[167] = t[110] ? x[102] : x[101];
  assign t[168] = ~(t[182]);
  assign t[169] = ~(t[83]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = ~(t[84]);
  assign t[171] = t[214] ^ t[183];
  assign t[172] = t[127] ? x[104] : x[103];
  assign t[173] = t[184] ? x[106] : x[105];
  assign t[174] = t[27] ? x[108] : x[107];
  assign t[175] = t[184] ? x[110] : x[109];
  assign t[176] = ~(t[185]);
  assign t[177] = ~(t[99]);
  assign t[178] = t[215] ^ t[186];
  assign t[179] = ~(t[153] ^ t[187]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[188] ^ t[182];
  assign t[181] = t[27] ? x[112] : x[111];
  assign t[182] = t[124] ^ t[84];
  assign t[183] = t[27] ? x[114] : x[113];
  assign t[184] = ~(t[144]);
  assign t[185] = t[135] ^ t[100];
  assign t[186] = t[184] ? x[116] : x[115];
  assign t[187] = t[123] ^ t[83];
  assign t[188] = t[83] ^ t[97];
  assign t[189] = t[216] ^ x[4];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[217] ^ x[9];
  assign t[191] = t[218] ^ x[12];
  assign t[192] = t[219] ^ x[15];
  assign t[193] = t[220] ^ x[18];
  assign t[194] = t[221] ^ x[21];
  assign t[195] = t[222] ^ x[24];
  assign t[196] = t[223] ^ x[27];
  assign t[197] = t[224] ^ x[30];
  assign t[198] = t[225] ^ x[33];
  assign t[199] = t[226] ^ x[36];
  assign t[19] = t[34] & t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[39];
  assign t[201] = t[228] ^ x[42];
  assign t[202] = t[229] ^ x[45];
  assign t[203] = t[230] ^ x[48];
  assign t[204] = t[231] ^ x[57];
  assign t[205] = t[232] ^ x[64];
  assign t[206] = t[233] ^ x[67];
  assign t[207] = t[234] ^ x[72];
  assign t[208] = t[235] ^ x[75];
  assign t[209] = t[236] ^ x[78];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[81];
  assign t[211] = t[238] ^ x[84];
  assign t[212] = t[239] ^ x[87];
  assign t[213] = t[240] ^ x[90];
  assign t[214] = t[241] ^ x[95];
  assign t[215] = t[242] ^ x[100];
  assign t[216] = (x[2] & x[3]);
  assign t[217] = (x[7] & x[8]);
  assign t[218] = (x[10] & x[11]);
  assign t[219] = (x[13] & x[14]);
  assign t[21] = ~(t[25] ^ t[38]);
  assign t[220] = (x[16] & x[17]);
  assign t[221] = (x[19] & x[20]);
  assign t[222] = (x[22] & x[23]);
  assign t[223] = (x[25] & x[26]);
  assign t[224] = (x[28] & x[29]);
  assign t[225] = (x[31] & x[32]);
  assign t[226] = (x[34] & x[35]);
  assign t[227] = (x[37] & x[38]);
  assign t[228] = (x[40] & x[41]);
  assign t[229] = (x[43] & x[44]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (x[46] & x[47]);
  assign t[231] = (x[55] & x[56]);
  assign t[232] = (x[62] & x[63]);
  assign t[233] = (x[65] & x[66]);
  assign t[234] = (x[70] & x[71]);
  assign t[235] = (x[73] & x[74]);
  assign t[236] = (x[76] & x[77]);
  assign t[237] = (x[79] & x[80]);
  assign t[238] = (x[82] & x[83]);
  assign t[239] = (x[85] & x[86]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (x[88] & x[89]);
  assign t[241] = (x[93] & x[94]);
  assign t[242] = (x[98] & x[99]);
  assign t[24] = ~(t[43] ^ t[44]);
  assign t[25] = t[45] ^ t[46];
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[190]);
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[192]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[7] ? t[51] : t[193];
  assign t[33] = t[7] ? t[52] : t[194];
  assign t[34] = ~(t[53]);
  assign t[35] = t[7] ? t[54] : t[195];
  assign t[36] = ~(t[55] ^ t[56]);
  assign t[37] = t[57] ^ t[58];
  assign t[38] = t[40] ^ t[59];
  assign t[39] = t[7] ? t[60] : t[196];
  assign t[3] = t[7] ? t[8] : t[189];
  assign t[40] = t[7] ? t[61] : t[197];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] & t[65];
  assign t[43] = t[12] ^ t[66];
  assign t[44] = t[67] ^ t[68];
  assign t[45] = t[53] ^ t[33];
  assign t[46] = t[69] ^ t[70];
  assign t[47] = ~(t[71] & t[72]);
  assign t[48] = t[198] | t[73];
  assign t[49] = ~(t[199]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[74] & t[200]);
  assign t[51] = t[193] ^ t[75];
  assign t[52] = t[194] ^ t[76];
  assign t[53] = t[7] ? t[77] : t[201];
  assign t[54] = t[195] ^ t[78];
  assign t[55] = t[79] ^ t[80];
  assign t[56] = ~(t[81] ^ t[82]);
  assign t[57] = t[83] ^ t[84];
  assign t[58] = t[85] & t[86];
  assign t[59] = t[41] ^ t[87];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[196] ^ t[88];
  assign t[61] = t[197] ^ t[89];
  assign t[62] = t[90] & t[91];
  assign t[63] = t[92] & t[93];
  assign t[64] = ~(t[62] ^ t[94]);
  assign t[65] = t[95] ^ t[96];
  assign t[66] = t[97] ^ t[98];
  assign t[67] = t[99] ^ t[100];
  assign t[68] = t[101] & t[102];
  assign t[69] = t[103] ^ t[19];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[104] & t[105];
  assign t[71] = ~(t[73] & t[106]);
  assign t[72] = ~(t[202] ^ t[107]);
  assign t[73] = ~(t[108] & t[109]);
  assign t[74] = ~(t[203]);
  assign t[75] = t[110] ? x[50] : x[49];
  assign t[76] = t[110] ? x[52] : x[51];
  assign t[77] = t[201] ^ t[111];
  assign t[78] = t[110] ? x[54] : x[53];
  assign t[79] = t[112] ^ t[113];
  assign t[7] = ~(t[14]);
  assign t[80] = t[114] ^ t[115];
  assign t[81] = t[116] ^ t[117];
  assign t[82] = t[118] ^ t[119];
  assign t[83] = t[26] ? t[120] : t[204];
  assign t[84] = t[192] ^ t[121];
  assign t[85] = ~(t[57] ^ t[122]);
  assign t[86] = t[123] ^ t[124];
  assign t[87] = t[125] & t[126];
  assign t[88] = t[127] ? x[59] : x[58];
  assign t[89] = t[127] ? x[61] : x[60];
  assign t[8] = t[189] ^ t[15];
  assign t[90] = ~(t[96]);
  assign t[91] = ~(t[128]);
  assign t[92] = ~(t[39]);
  assign t[93] = t[7] ? t[129] : t[205];
  assign t[94] = t[22] ^ t[128];
  assign t[95] = t[128] ^ t[40];
  assign t[96] = t[93] ^ t[39];
  assign t[97] = t[199] ^ t[130];
  assign t[98] = t[122] ^ t[58];
  assign t[99] = ~t[131];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind98(x, y);
 input [116:0] x;
 output y;

 wire [225:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[136] ? x[64] : x[63];
  assign t[101] = ~(t[107]);
  assign t[102] = ~(t[84]);
  assign t[103] = ~(t[40]);
  assign t[104] = t[7] ? t[137] : t[191];
  assign t[105] = t[22] ^ t[84];
  assign t[106] = t[84] ^ t[41];
  assign t[107] = t[104] ^ t[40];
  assign t[108] = t[79] ? x[69] : x[68];
  assign t[109] = ~(t[138]);
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = ~(t[123]);
  assign t[111] = ~(t[124]);
  assign t[112] = t[175] ^ t[139];
  assign t[113] = t[124] ^ t[24];
  assign t[114] = ~(t[140] & t[141]);
  assign t[115] = t[142] ^ t[192];
  assign t[116] = ~(t[185]);
  assign t[117] = t[143] & t[142];
  assign t[118] = t[187] ^ t[144];
  assign t[119] = t[89] ? t[145] : t[193];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[188] ^ t[146];
  assign t[121] = t[189] ^ t[147];
  assign t[122] = t[148] & t[149];
  assign t[123] = t[7] ? t[150] : t[194];
  assign t[124] = t[174] ^ t[151];
  assign t[125] = t[152] ? x[80] : x[79];
  assign t[126] = t[153] & t[154];
  assign t[127] = ~(t[155] ^ t[91]);
  assign t[128] = t[156] ^ t[83];
  assign t[129] = t[79] ? x[82] : x[81];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[27] ? x[84] : x[83];
  assign t[131] = ~(t[157]);
  assign t[132] = ~(t[36]);
  assign t[133] = ~(t[37]);
  assign t[134] = t[26] ? t[158] : t[195];
  assign t[135] = t[190] ^ t[159];
  assign t[136] = ~(t[49]);
  assign t[137] = t[191] ^ t[160];
  assign t[138] = t[112] ^ t[124];
  assign t[139] = t[7] ? t[161] : t[196];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[143] | t[142]);
  assign t[141] = ~(t[162] | t[116]);
  assign t[142] = ~(t[197]);
  assign t[143] = ~(t[192]);
  assign t[144] = t[152] ? x[95] : x[94];
  assign t[145] = t[193] ^ t[163];
  assign t[146] = t[152] ? x[97] : x[96];
  assign t[147] = t[136] ? x[99] : x[98];
  assign t[148] = ~(t[95] ^ t[164]);
  assign t[149] = t[165] ^ t[157];
  assign t[14] = ~(t[26]);
  assign t[150] = t[194] ^ t[166];
  assign t[151] = t[26] ? t[167] : t[198];
  assign t[152] = ~(t[49]);
  assign t[153] = ~(t[168]);
  assign t[154] = ~(t[81]);
  assign t[155] = t[81] ^ t[119];
  assign t[156] = t[119] ^ t[58];
  assign t[157] = t[64] ^ t[37];
  assign t[158] = t[195] ^ t[169];
  assign t[159] = t[136] ? x[104] : x[103];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[136] ? x[106] : x[105];
  assign t[161] = t[196] ^ t[170];
  assign t[162] = ~(t[180]);
  assign t[163] = t[152] ? x[108] : x[107];
  assign t[164] = t[63] ^ t[36];
  assign t[165] = t[36] ^ t[97];
  assign t[166] = t[79] ? x[110] : x[109];
  assign t[167] = t[198] ^ t[171];
  assign t[168] = t[83] ^ t[119];
  assign t[169] = t[79] ? x[112] : x[111];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[27] ? x[114] : x[113];
  assign t[171] = t[27] ? x[116] : x[115];
  assign t[172] = t[199] ^ x[4];
  assign t[173] = t[200] ^ x[9];
  assign t[174] = t[201] ^ x[12];
  assign t[175] = t[202] ^ x[15];
  assign t[176] = t[203] ^ x[18];
  assign t[177] = t[204] ^ x[21];
  assign t[178] = t[205] ^ x[24];
  assign t[179] = t[206] ^ x[27];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[207] ^ x[30];
  assign t[181] = t[208] ^ x[33];
  assign t[182] = t[209] ^ x[36];
  assign t[183] = t[210] ^ x[39];
  assign t[184] = t[211] ^ x[42];
  assign t[185] = t[212] ^ x[45];
  assign t[186] = t[213] ^ x[48];
  assign t[187] = t[214] ^ x[51];
  assign t[188] = t[215] ^ x[54];
  assign t[189] = t[216] ^ x[57];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[217] ^ x[60];
  assign t[191] = t[218] ^ x[67];
  assign t[192] = t[219] ^ x[72];
  assign t[193] = t[220] ^ x[75];
  assign t[194] = t[221] ^ x[78];
  assign t[195] = t[222] ^ x[87];
  assign t[196] = t[223] ^ x[90];
  assign t[197] = t[224] ^ x[93];
  assign t[198] = t[225] ^ x[102];
  assign t[199] = (x[2] & x[3]);
  assign t[19] = ~(t[34] ^ t[35]);
  assign t[1] = ~(t[4]);
  assign t[200] = (x[7] & x[8]);
  assign t[201] = (x[10] & x[11]);
  assign t[202] = (x[13] & x[14]);
  assign t[203] = (x[16] & x[17]);
  assign t[204] = (x[19] & x[20]);
  assign t[205] = (x[22] & x[23]);
  assign t[206] = (x[25] & x[26]);
  assign t[207] = (x[28] & x[29]);
  assign t[208] = (x[31] & x[32]);
  assign t[209] = (x[34] & x[35]);
  assign t[20] = t[36] ^ t[37];
  assign t[210] = (x[37] & x[38]);
  assign t[211] = (x[40] & x[41]);
  assign t[212] = (x[43] & x[44]);
  assign t[213] = (x[46] & x[47]);
  assign t[214] = (x[49] & x[50]);
  assign t[215] = (x[52] & x[53]);
  assign t[216] = (x[55] & x[56]);
  assign t[217] = (x[58] & x[59]);
  assign t[218] = (x[65] & x[66]);
  assign t[219] = (x[70] & x[71]);
  assign t[21] = t[38] & t[39];
  assign t[220] = (x[73] & x[74]);
  assign t[221] = (x[76] & x[77]);
  assign t[222] = (x[85] & x[86]);
  assign t[223] = (x[88] & x[89]);
  assign t[224] = (x[91] & x[92]);
  assign t[225] = (x[100] & x[101]);
  assign t[22] = t[40] ^ t[41];
  assign t[23] = t[42] ^ t[43];
  assign t[24] = t[173] ^ t[44];
  assign t[25] = t[45] ^ t[46];
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49]);
  assign t[28] = ~(t[174]);
  assign t[29] = ~(t[175]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[176]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = t[52] ^ t[53];
  assign t[33] = t[54] ^ t[55];
  assign t[34] = t[56] ^ t[57];
  assign t[35] = t[58] ^ t[59];
  assign t[36] = ~t[60];
  assign t[37] = t[61];
  assign t[38] = ~(t[20] ^ t[62]);
  assign t[39] = t[63] ^ t[64];
  assign t[3] = t[7] ? t[8] : t[172];
  assign t[40] = t[7] ? t[65] : t[177];
  assign t[41] = t[7] ? t[66] : t[178];
  assign t[42] = t[67] ^ t[68];
  assign t[43] = t[69] & t[70];
  assign t[44] = t[7] ? t[71] : t[179];
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] & t[75];
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = t[180] | t[78];
  assign t[49] = ~(t[79]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[181]);
  assign t[51] = ~(t[80] & t[173]);
  assign t[52] = t[81] ^ t[58];
  assign t[53] = t[82] & t[83];
  assign t[54] = t[84] ^ t[40];
  assign t[55] = t[85] & t[86];
  assign t[56] = t[63] ^ t[87];
  assign t[57] = t[88] ^ t[46];
  assign t[58] = t[89] ? t[90] : t[182];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[26] ? t[93] : t[183];
  assign t[61] = t[26] ? t[94] : t[184];
  assign t[62] = t[95] ^ t[96];
  assign t[63] = t[37] ^ t[97];
  assign t[64] = t[98];
  assign t[65] = t[177] ^ t[99];
  assign t[66] = t[178] ^ t[100];
  assign t[67] = t[101] & t[102];
  assign t[68] = t[103] & t[104];
  assign t[69] = ~(t[67] ^ t[105]);
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[106] ^ t[107];
  assign t[71] = t[179] ^ t[108];
  assign t[72] = t[109] & t[110];
  assign t[73] = t[111] & t[112];
  assign t[74] = ~(t[88] ^ t[45]);
  assign t[75] = t[113] ^ t[112];
  assign t[76] = ~(t[78] & t[114]);
  assign t[77] = ~(t[185] ^ t[115]);
  assign t[78] = ~(t[116] & t[117]);
  assign t[79] = ~(t[48]);
  assign t[7] = ~(t[14]);
  assign t[80] = ~(t[186]);
  assign t[81] = t[89] ? t[118] : t[187];
  assign t[82] = ~(t[119]);
  assign t[83] = t[89] ? t[120] : t[188];
  assign t[84] = t[7] ? t[121] : t[189];
  assign t[85] = ~(t[54] ^ t[42]);
  assign t[86] = t[22] ^ t[104];
  assign t[87] = t[62] ^ t[122];
  assign t[88] = t[123] ^ t[124];
  assign t[89] = ~(t[14]);
  assign t[8] = t[172] ^ t[15];
  assign t[90] = t[182] ^ t[125];
  assign t[91] = t[126] ^ t[53];
  assign t[92] = t[127] & t[128];
  assign t[93] = t[183] ^ t[129];
  assign t[94] = t[184] ^ t[130];
  assign t[95] = t[131] & t[132];
  assign t[96] = t[133] & t[64];
  assign t[97] = ~t[134];
  assign t[98] = t[26] ? t[135] : t[190];
  assign t[99] = t[136] ? x[62] : x[61];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind99(x, y);
 input [116:0] x;
 output y;

 wire [234:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[133] & t[134];
  assign t[101] = ~(t[113] ^ t[67]);
  assign t[102] = t[135] ^ t[39];
  assign t[103] = t[136] ? x[65] : x[64];
  assign t[104] = t[136] ? x[67] : x[66];
  assign t[105] = t[137] & t[138];
  assign t[106] = t[193] ^ t[139];
  assign t[107] = ~(t[140] & t[141]);
  assign t[108] = t[142] ^ t[201];
  assign t[109] = ~(t[194]);
  assign t[10] = ~(t[18] ^ t[19]);
  assign t[110] = t[143] & t[142];
  assign t[111] = t[196] ^ t[144];
  assign t[112] = ~(t[44]);
  assign t[113] = t[36] ^ t[62];
  assign t[114] = t[145] ? t[146] : t[202];
  assign t[115] = t[117] ^ t[147];
  assign t[116] = t[145] ? t[148] : t[203];
  assign t[117] = t[149] ^ t[150];
  assign t[118] = t[151] & t[152];
  assign t[119] = t[197] ^ t[153];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[7] ? t[154] : t[204];
  assign t[121] = t[198] ^ t[155];
  assign t[122] = ~(t[156] ^ t[65]);
  assign t[123] = t[40] ^ t[89];
  assign t[124] = t[77] ? x[81] : x[80];
  assign t[125] = t[77] ? x[83] : x[82];
  assign t[126] = t[199] ^ t[157];
  assign t[127] = t[136] ? x[85] : x[84];
  assign t[128] = t[200] ^ t[158];
  assign t[129] = ~(t[132]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = ~(t[87]);
  assign t[131] = t[40] ^ t[87];
  assign t[132] = t[89] ^ t[64];
  assign t[133] = ~(t[159]);
  assign t[134] = ~(t[36]);
  assign t[135] = t[62] ^ t[37];
  assign t[136] = ~(t[49]);
  assign t[137] = ~(t[160]);
  assign t[138] = ~(t[43]);
  assign t[139] = t[136] ? x[87] : x[86];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[143] | t[142]);
  assign t[141] = ~(t[161] | t[109]);
  assign t[142] = ~(t[205]);
  assign t[143] = ~(t[201]);
  assign t[144] = t[136] ? x[92] : x[91];
  assign t[145] = ~(t[14]);
  assign t[146] = t[202] ^ t[162];
  assign t[147] = t[163] & t[164];
  assign t[148] = t[203] ^ t[165];
  assign t[149] = t[166] & t[167];
  assign t[14] = ~(t[26]);
  assign t[150] = t[168] & t[169];
  assign t[151] = ~(t[149] ^ t[170]);
  assign t[152] = t[171] ^ t[172];
  assign t[153] = t[77] ? x[94] : x[93];
  assign t[154] = t[204] ^ t[173];
  assign t[155] = t[77] ? x[96] : x[95];
  assign t[156] = t[87] ^ t[64];
  assign t[157] = t[27] ? x[98] : x[97];
  assign t[158] = t[27] ? x[100] : x[99];
  assign t[159] = t[39] ^ t[62];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[73] ^ t[44];
  assign t[161] = ~(t[187]);
  assign t[162] = t[174] ? x[102] : x[101];
  assign t[163] = ~(t[175] ^ t[117]);
  assign t[164] = t[85] ^ t[169];
  assign t[165] = t[174] ? x[104] : x[103];
  assign t[166] = ~(t[172]);
  assign t[167] = ~(t[176]);
  assign t[168] = ~(t[116]);
  assign t[169] = t[145] ? t[177] : t[206];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[85] ^ t[176];
  assign t[171] = t[176] ^ t[114];
  assign t[172] = t[169] ^ t[116];
  assign t[173] = t[27] ? x[109] : x[108];
  assign t[174] = ~(t[49]);
  assign t[175] = t[176] ^ t[116];
  assign t[176] = t[145] ? t[178] : t[207];
  assign t[177] = t[206] ^ t[179];
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[174] ? x[114] : x[113];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[174] ? x[116] : x[115];
  assign t[181] = t[208] ^ x[4];
  assign t[182] = t[209] ^ x[9];
  assign t[183] = t[210] ^ x[12];
  assign t[184] = t[211] ^ x[15];
  assign t[185] = t[212] ^ x[18];
  assign t[186] = t[213] ^ x[21];
  assign t[187] = t[214] ^ x[24];
  assign t[188] = t[215] ^ x[27];
  assign t[189] = t[216] ^ x[30];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[217] ^ x[33];
  assign t[191] = t[218] ^ x[36];
  assign t[192] = t[219] ^ x[39];
  assign t[193] = t[220] ^ x[42];
  assign t[194] = t[221] ^ x[45];
  assign t[195] = t[222] ^ x[48];
  assign t[196] = t[223] ^ x[51];
  assign t[197] = t[224] ^ x[54];
  assign t[198] = t[225] ^ x[57];
  assign t[199] = t[226] ^ x[60];
  assign t[19] = ~(t[34] ^ t[35]);
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[63];
  assign t[201] = t[228] ^ x[70];
  assign t[202] = t[229] ^ x[73];
  assign t[203] = t[230] ^ x[76];
  assign t[204] = t[231] ^ x[79];
  assign t[205] = t[232] ^ x[90];
  assign t[206] = t[233] ^ x[107];
  assign t[207] = t[234] ^ x[112];
  assign t[208] = (x[2] & x[3]);
  assign t[209] = (x[7] & x[8]);
  assign t[20] = t[36] ^ t[37];
  assign t[210] = (x[10] & x[11]);
  assign t[211] = (x[13] & x[14]);
  assign t[212] = (x[16] & x[17]);
  assign t[213] = (x[19] & x[20]);
  assign t[214] = (x[22] & x[23]);
  assign t[215] = (x[25] & x[26]);
  assign t[216] = (x[28] & x[29]);
  assign t[217] = (x[31] & x[32]);
  assign t[218] = (x[34] & x[35]);
  assign t[219] = (x[37] & x[38]);
  assign t[21] = t[38] & t[39];
  assign t[220] = (x[40] & x[41]);
  assign t[221] = (x[43] & x[44]);
  assign t[222] = (x[46] & x[47]);
  assign t[223] = (x[49] & x[50]);
  assign t[224] = (x[52] & x[53]);
  assign t[225] = (x[55] & x[56]);
  assign t[226] = (x[58] & x[59]);
  assign t[227] = (x[61] & x[62]);
  assign t[228] = (x[68] & x[69]);
  assign t[229] = (x[71] & x[72]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (x[74] & x[75]);
  assign t[231] = (x[77] & x[78]);
  assign t[232] = (x[88] & x[89]);
  assign t[233] = (x[105] & x[106]);
  assign t[234] = (x[110] & x[111]);
  assign t[23] = t[37] ^ t[42];
  assign t[24] = t[43] ^ t[44];
  assign t[25] = t[45] & t[46];
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49]);
  assign t[28] = ~(t[182]);
  assign t[29] = ~(t[183]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[184]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = t[52] ^ t[53];
  assign t[33] = ~(t[54] ^ t[55]);
  assign t[34] = t[56] ^ t[57];
  assign t[35] = t[58] ^ t[59];
  assign t[36] = ~t[60];
  assign t[37] = ~t[61];
  assign t[38] = ~(t[62]);
  assign t[39] = t[63];
  assign t[3] = t[7] ? t[8] : t[181];
  assign t[40] = t[64] ^ t[58];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] ^ t[68];
  assign t[43] = t[7] ? t[69] : t[185];
  assign t[44] = t[7] ? t[70] : t[186];
  assign t[45] = ~(t[24] ^ t[71]);
  assign t[46] = t[72] ^ t[73];
  assign t[47] = ~(t[74] & t[75]);
  assign t[48] = t[187] | t[76];
  assign t[49] = ~(t[77]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[188]);
  assign t[51] = ~(t[78] & t[189]);
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] ^ t[82];
  assign t[54] = ~(t[83] ^ t[84]);
  assign t[55] = t[85] ^ t[86];
  assign t[56] = t[87] ^ t[58];
  assign t[57] = t[88] & t[89];
  assign t[58] = t[189] ^ t[90];
  assign t[59] = t[65] ^ t[91];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[26] ? t[92] : t[190];
  assign t[61] = t[26] ? t[93] : t[191];
  assign t[62] = t[94];
  assign t[63] = t[26] ? t[95] : t[192];
  assign t[64] = t[182] ^ t[96];
  assign t[65] = t[97] ^ t[57];
  assign t[66] = t[98] & t[99];
  assign t[67] = t[100] ^ t[21];
  assign t[68] = t[101] & t[102];
  assign t[69] = t[185] ^ t[103];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[186] ^ t[104];
  assign t[71] = t[105] ^ t[82];
  assign t[72] = t[44] ^ t[79];
  assign t[73] = t[7] ? t[106] : t[193];
  assign t[74] = ~(t[76] & t[107]);
  assign t[75] = ~(t[194] ^ t[108]);
  assign t[76] = ~(t[109] & t[110]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[195]);
  assign t[79] = t[7] ? t[111] : t[196];
  assign t[7] = ~(t[14]);
  assign t[80] = t[71] ^ t[25];
  assign t[81] = t[43] ^ t[79];
  assign t[82] = t[112] & t[73];
  assign t[83] = t[113] ^ t[68];
  assign t[84] = t[114] ^ t[115];
  assign t[85] = t[116] ^ t[114];
  assign t[86] = t[117] ^ t[118];
  assign t[87] = t[7] ? t[119] : t[197];
  assign t[88] = ~(t[64]);
  assign t[89] = t[183] ^ t[120];
  assign t[8] = t[181] ^ t[15];
  assign t[90] = t[7] ? t[121] : t[198];
  assign t[91] = t[122] & t[123];
  assign t[92] = t[190] ^ t[124];
  assign t[93] = t[191] ^ t[125];
  assign t[94] = t[26] ? t[126] : t[199];
  assign t[95] = t[192] ^ t[127];
  assign t[96] = t[26] ? t[128] : t[200];
  assign t[97] = t[129] & t[130];
  assign t[98] = ~(t[97] ^ t[131]);
  assign t[99] = t[56] ^ t[132];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind100(x, y);
 input [116:0] x;
 output y;

 wire [245:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[132] ^ t[133];
  assign t[101] = t[134] ^ t[38];
  assign t[102] = t[201] ^ t[135];
  assign t[103] = t[121] ^ t[64];
  assign t[104] = ~(t[136] & t[137]);
  assign t[105] = t[138] ^ t[207];
  assign t[106] = ~(t[204]);
  assign t[107] = t[139] & t[138];
  assign t[108] = t[37] ^ t[56];
  assign t[109] = t[77] ? x[59] : x[58];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[75] ? x[61] : x[60];
  assign t[111] = ~(t[140]);
  assign t[112] = ~(t[134]);
  assign t[113] = ~(t[89]);
  assign t[114] = t[141];
  assign t[115] = t[134] ^ t[89];
  assign t[116] = t[26] ? t[142] : t[208];
  assign t[117] = ~(t[85] ^ t[143]);
  assign t[118] = t[101] ^ t[140];
  assign t[119] = t[206] ^ t[144];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[26] ? t[145] : t[209];
  assign t[121] = t[146] ^ t[147];
  assign t[122] = t[92] ^ t[102];
  assign t[123] = t[195] ^ t[148];
  assign t[124] = t[121] ^ t[149];
  assign t[125] = t[150] ? t[151] : t[210];
  assign t[126] = t[150] ? t[152] : t[211];
  assign t[127] = ~(t[96] ^ t[132]);
  assign t[128] = t[99] ^ t[153];
  assign t[129] = ~(t[52] ^ t[154]);
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[20] ^ t[108];
  assign t[131] = t[150] ? t[155] : t[212];
  assign t[132] = t[156] ^ t[157];
  assign t[133] = t[158] & t[159];
  assign t[134] = ~t[160];
  assign t[135] = t[7] ? t[161] : t[213];
  assign t[136] = ~(t[139] | t[138]);
  assign t[137] = ~(t[162] | t[106]);
  assign t[138] = ~(t[214]);
  assign t[139] = ~(t[207]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[114] ^ t[89];
  assign t[141] = t[26] ? t[163] : t[215];
  assign t[142] = t[208] ^ t[164];
  assign t[143] = t[61] ^ t[134];
  assign t[144] = t[75] ? x[87] : x[86];
  assign t[145] = t[209] ^ t[165];
  assign t[146] = t[166] & t[167];
  assign t[147] = t[168] & t[123];
  assign t[148] = t[7] ? t[169] : t[216];
  assign t[149] = t[170] & t[171];
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[14]);
  assign t[151] = t[210] ^ t[172];
  assign t[152] = t[211] ^ t[173];
  assign t[153] = t[150] ? t[174] : t[217];
  assign t[154] = t[67] ^ t[35];
  assign t[155] = t[212] ^ t[175];
  assign t[156] = t[176] & t[177];
  assign t[157] = t[178] & t[153];
  assign t[158] = ~(t[156] ^ t[179]);
  assign t[159] = t[180] ^ t[181];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[26] ? t[182] : t[218];
  assign t[161] = t[213] ^ t[183];
  assign t[162] = ~(t[199]);
  assign t[163] = t[215] ^ t[184];
  assign t[164] = t[27] ? x[98] : x[97];
  assign t[165] = t[27] ? x[100] : x[99];
  assign t[166] = ~(t[185]);
  assign t[167] = ~(t[91]);
  assign t[168] = ~(t[92]);
  assign t[169] = t[216] ^ t[186];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = ~(t[146] ^ t[187]);
  assign t[171] = t[188] ^ t[185];
  assign t[172] = t[189] ? x[102] : x[101];
  assign t[173] = t[189] ? x[104] : x[103];
  assign t[174] = t[217] ^ t[190];
  assign t[175] = t[189] ? x[106] : x[105];
  assign t[176] = ~(t[181]);
  assign t[177] = ~(t[125]);
  assign t[178] = ~(t[126]);
  assign t[179] = t[99] ^ t[125];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[125] ^ t[131];
  assign t[181] = t[153] ^ t[126];
  assign t[182] = t[218] ^ t[191];
  assign t[183] = t[75] ? x[108] : x[107];
  assign t[184] = t[77] ? x[110] : x[109];
  assign t[185] = t[123] ^ t[92];
  assign t[186] = t[27] ? x[112] : x[111];
  assign t[187] = t[122] ^ t[91];
  assign t[188] = t[91] ^ t[102];
  assign t[189] = ~(t[48]);
  assign t[18] = t[7] ? t[32] : t[193];
  assign t[190] = t[189] ? x[114] : x[113];
  assign t[191] = t[75] ? x[116] : x[115];
  assign t[192] = t[219] ^ x[4];
  assign t[193] = t[220] ^ x[9];
  assign t[194] = t[221] ^ x[12];
  assign t[195] = t[222] ^ x[15];
  assign t[196] = t[223] ^ x[18];
  assign t[197] = t[224] ^ x[21];
  assign t[198] = t[225] ^ x[24];
  assign t[199] = t[226] ^ x[27];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[30];
  assign t[201] = t[228] ^ x[33];
  assign t[202] = t[229] ^ x[38];
  assign t[203] = t[230] ^ x[41];
  assign t[204] = t[231] ^ x[44];
  assign t[205] = t[232] ^ x[47];
  assign t[206] = t[233] ^ x[54];
  assign t[207] = t[234] ^ x[57];
  assign t[208] = t[235] ^ x[64];
  assign t[209] = t[236] ^ x[67];
  assign t[20] = t[35] ^ t[18];
  assign t[210] = t[237] ^ x[70];
  assign t[211] = t[238] ^ x[73];
  assign t[212] = t[239] ^ x[76];
  assign t[213] = t[240] ^ x[79];
  assign t[214] = t[241] ^ x[82];
  assign t[215] = t[242] ^ x[85];
  assign t[216] = t[243] ^ x[90];
  assign t[217] = t[244] ^ x[93];
  assign t[218] = t[245] ^ x[96];
  assign t[219] = (x[2] & x[3]);
  assign t[21] = t[36] & t[37];
  assign t[220] = (x[7] & x[8]);
  assign t[221] = (x[10] & x[11]);
  assign t[222] = (x[13] & x[14]);
  assign t[223] = (x[16] & x[17]);
  assign t[224] = (x[19] & x[20]);
  assign t[225] = (x[22] & x[23]);
  assign t[226] = (x[25] & x[26]);
  assign t[227] = (x[28] & x[29]);
  assign t[228] = (x[31] & x[32]);
  assign t[229] = (x[36] & x[37]);
  assign t[22] = t[38] ^ t[39];
  assign t[230] = (x[39] & x[40]);
  assign t[231] = (x[42] & x[43]);
  assign t[232] = (x[45] & x[46]);
  assign t[233] = (x[52] & x[53]);
  assign t[234] = (x[55] & x[56]);
  assign t[235] = (x[62] & x[63]);
  assign t[236] = (x[65] & x[66]);
  assign t[237] = (x[68] & x[69]);
  assign t[238] = (x[71] & x[72]);
  assign t[239] = (x[74] & x[75]);
  assign t[23] = t[40] ^ t[41];
  assign t[240] = (x[77] & x[78]);
  assign t[241] = (x[80] & x[81]);
  assign t[242] = (x[83] & x[84]);
  assign t[243] = (x[88] & x[89]);
  assign t[244] = (x[91] & x[92]);
  assign t[245] = (x[94] & x[95]);
  assign t[24] = ~(t[42] ^ t[43]);
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[194]);
  assign t[29] = ~(t[195]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = ~(t[196]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[193] ^ t[51];
  assign t[33] = t[52] ^ t[21];
  assign t[34] = t[53] & t[54];
  assign t[35] = t[7] ? t[55] : t[197];
  assign t[36] = ~(t[56]);
  assign t[37] = t[7] ? t[57] : t[198];
  assign t[38] = ~t[58];
  assign t[39] = t[59] ^ t[60];
  assign t[3] = t[7] ? t[8] : t[192];
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = ~(t[65] ^ t[66]);
  assign t[43] = t[67] ^ t[68];
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[10] ^ t[71]);
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[199] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[200]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[76] & t[201]);
  assign t[51] = t[77] ? x[35] : x[34];
  assign t[52] = t[78] & t[79];
  assign t[53] = ~(t[80] ^ t[33]);
  assign t[54] = t[67] ^ t[37];
  assign t[55] = t[197] ^ t[81];
  assign t[56] = t[7] ? t[82] : t[202];
  assign t[57] = t[198] ^ t[83];
  assign t[58] = t[26] ? t[84] : t[203];
  assign t[59] = t[85] ^ t[86];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[87] & t[88];
  assign t[61] = t[89] ^ t[38];
  assign t[62] = t[59] ^ t[90];
  assign t[63] = t[91] ^ t[92];
  assign t[64] = t[93] & t[94];
  assign t[65] = t[95] ^ t[22];
  assign t[66] = t[96] ^ t[97];
  assign t[67] = t[56] ^ t[18];
  assign t[68] = t[33] ^ t[98];
  assign t[69] = t[99] ^ t[100];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[101] ^ t[86];
  assign t[71] = t[102] ^ t[103];
  assign t[72] = ~(t[74] & t[104]);
  assign t[73] = ~(t[204] ^ t[105]);
  assign t[74] = ~(t[106] & t[107]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[205]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[108]);
  assign t[79] = ~(t[35]);
  assign t[7] = ~(t[14]);
  assign t[80] = t[35] ^ t[56];
  assign t[81] = t[77] ? x[49] : x[48];
  assign t[82] = t[202] ^ t[109];
  assign t[83] = t[77] ? x[51] : x[50];
  assign t[84] = t[203] ^ t[110];
  assign t[85] = t[111] & t[112];
  assign t[86] = t[113] & t[114];
  assign t[87] = ~(t[115] ^ t[59]);
  assign t[88] = t[61] ^ t[114];
  assign t[89] = t[116];
  assign t[8] = t[192] ^ t[15];
  assign t[90] = t[117] & t[118];
  assign t[91] = t[7] ? t[119] : t[206];
  assign t[92] = t[194] ^ t[120];
  assign t[93] = ~(t[63] ^ t[121]);
  assign t[94] = t[122] ^ t[123];
  assign t[95] = t[122] ^ t[124];
  assign t[96] = t[125] ^ t[126];
  assign t[97] = t[127] & t[128];
  assign t[98] = t[129] & t[130];
  assign t[99] = t[126] ^ t[131];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind101(x, y);
 input [116:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[128]);
  assign t[101] = ~(t[130]);
  assign t[102] = ~(t[65]);
  assign t[103] = t[7] ? t[131] : t[190];
  assign t[104] = t[130] ^ t[65];
  assign t[105] = ~(t[132] & t[133]);
  assign t[106] = t[134] ^ t[191];
  assign t[107] = ~(t[185]);
  assign t[108] = t[135] & t[134];
  assign t[109] = t[27] ? x[72] : x[71];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[187] ^ t[136];
  assign t[111] = t[137] ? x[74] : x[73];
  assign t[112] = t[137] ? x[76] : x[75];
  assign t[113] = t[27] ? x[78] : x[77];
  assign t[114] = ~t[138];
  assign t[115] = t[26] ? t[139] : t[192];
  assign t[116] = t[140] ^ t[19];
  assign t[117] = t[141] & t[142];
  assign t[118] = t[143] & t[144];
  assign t[119] = ~(t[14]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[188] ^ t[145];
  assign t[121] = t[189] ^ t[146];
  assign t[122] = t[147] ^ t[148];
  assign t[123] = t[93] ^ t[149];
  assign t[124] = t[119] ? t[150] : t[193];
  assign t[125] = t[99] ? x[86] : x[85];
  assign t[126] = t[42] ^ t[130];
  assign t[127] = t[130] ^ t[24];
  assign t[128] = t[103] ^ t[65];
  assign t[129] = ~(t[27]);
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[7] ? t[151] : t[194];
  assign t[131] = t[190] ^ t[152];
  assign t[132] = ~(t[135] | t[134]);
  assign t[133] = ~(t[153] | t[107]);
  assign t[134] = ~(t[195]);
  assign t[135] = ~(t[191]);
  assign t[136] = t[137] ? x[94] : x[93];
  assign t[137] = ~(t[129]);
  assign t[138] = t[26] ? t[154] : t[196];
  assign t[139] = t[192] ^ t[155];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[156] & t[157];
  assign t[141] = ~(t[140] ^ t[158]);
  assign t[142] = t[18] ^ t[159];
  assign t[143] = ~(t[160] ^ t[38]);
  assign t[144] = t[20] ^ t[85];
  assign t[145] = t[161] ? x[99] : x[98];
  assign t[146] = t[161] ? x[101] : x[100];
  assign t[147] = t[162] & t[163];
  assign t[148] = t[164] & t[124];
  assign t[149] = t[119] ? t[165] : t[197];
  assign t[14] = ~(t[26]);
  assign t[150] = t[193] ^ t[166];
  assign t[151] = t[194] ^ t[167];
  assign t[152] = t[99] ? x[106] : x[105];
  assign t[153] = ~(t[178]);
  assign t[154] = t[196] ^ t[168];
  assign t[155] = t[99] ? x[108] : x[107];
  assign t[156] = ~(t[159]);
  assign t[157] = ~(t[32]);
  assign t[158] = t[89] ^ t[32];
  assign t[159] = t[35] ^ t[53];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[114] ^ t[36];
  assign t[161] = ~(t[129]);
  assign t[162] = ~(t[169]);
  assign t[163] = ~(t[92]);
  assign t[164] = ~(t[93]);
  assign t[165] = t[197] ^ t[170];
  assign t[166] = t[161] ? x[110] : x[109];
  assign t[167] = t[99] ? x[112] : x[111];
  assign t[168] = t[27] ? x[114] : x[113];
  assign t[169] = t[124] ^ t[93];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[161] ? x[116] : x[115];
  assign t[171] = t[198] ^ x[4];
  assign t[172] = t[199] ^ x[9];
  assign t[173] = t[200] ^ x[12];
  assign t[174] = t[201] ^ x[15];
  assign t[175] = t[202] ^ x[18];
  assign t[176] = t[203] ^ x[21];
  assign t[177] = t[204] ^ x[24];
  assign t[178] = t[205] ^ x[27];
  assign t[179] = t[206] ^ x[30];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[207] ^ x[33];
  assign t[181] = t[208] ^ x[36];
  assign t[182] = t[209] ^ x[39];
  assign t[183] = t[210] ^ x[42];
  assign t[184] = t[211] ^ x[45];
  assign t[185] = t[212] ^ x[50];
  assign t[186] = t[213] ^ x[53];
  assign t[187] = t[214] ^ x[58];
  assign t[188] = t[215] ^ x[61];
  assign t[189] = t[216] ^ x[64];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[217] ^ x[67];
  assign t[191] = t[218] ^ x[70];
  assign t[192] = t[219] ^ x[81];
  assign t[193] = t[220] ^ x[84];
  assign t[194] = t[221] ^ x[89];
  assign t[195] = t[222] ^ x[92];
  assign t[196] = t[223] ^ x[97];
  assign t[197] = t[224] ^ x[104];
  assign t[198] = (x[2] & x[3]);
  assign t[199] = (x[7] & x[8]);
  assign t[19] = t[34] & t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[10] & x[11]);
  assign t[201] = (x[13] & x[14]);
  assign t[202] = (x[16] & x[17]);
  assign t[203] = (x[19] & x[20]);
  assign t[204] = (x[22] & x[23]);
  assign t[205] = (x[25] & x[26]);
  assign t[206] = (x[28] & x[29]);
  assign t[207] = (x[31] & x[32]);
  assign t[208] = (x[34] & x[35]);
  assign t[209] = (x[37] & x[38]);
  assign t[20] = t[36] ^ t[37];
  assign t[210] = (x[40] & x[41]);
  assign t[211] = (x[43] & x[44]);
  assign t[212] = (x[48] & x[49]);
  assign t[213] = (x[51] & x[52]);
  assign t[214] = (x[56] & x[57]);
  assign t[215] = (x[59] & x[60]);
  assign t[216] = (x[62] & x[63]);
  assign t[217] = (x[65] & x[66]);
  assign t[218] = (x[68] & x[69]);
  assign t[219] = (x[79] & x[80]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = (x[82] & x[83]);
  assign t[221] = (x[87] & x[88]);
  assign t[222] = (x[90] & x[91]);
  assign t[223] = (x[95] & x[96]);
  assign t[224] = (x[102] & x[103]);
  assign t[22] = ~(t[40] ^ t[41]);
  assign t[23] = t[42] ^ t[43];
  assign t[24] = t[7] ? t[44] : t[172];
  assign t[25] = t[45] ^ t[46];
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[173]);
  assign t[29] = ~(t[174]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[175]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[7] ? t[51] : t[176];
  assign t[33] = t[177] ^ t[52];
  assign t[34] = ~(t[53]);
  assign t[35] = t[174] ^ t[54];
  assign t[36] = t[55];
  assign t[37] = ~t[56];
  assign t[38] = t[57] ^ t[58];
  assign t[39] = t[59] & t[60];
  assign t[3] = t[7] ? t[8] : t[171];
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] ^ t[24];
  assign t[43] = t[45] ^ t[66];
  assign t[44] = t[172] ^ t[67];
  assign t[45] = t[68] ^ t[69];
  assign t[46] = t[70] & t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[178] | t[74];
  assign t[49] = ~(t[179]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[75] & t[177]);
  assign t[51] = t[176] ^ t[76];
  assign t[52] = t[7] ? t[77] : t[180];
  assign t[53] = t[173] ^ t[78];
  assign t[54] = t[7] ? t[79] : t[181];
  assign t[55] = t[26] ? t[80] : t[182];
  assign t[56] = t[26] ? t[81] : t[183];
  assign t[57] = t[82] & t[83];
  assign t[58] = t[84] & t[85];
  assign t[59] = ~(t[57] ^ t[86]);
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[87] ^ t[88];
  assign t[61] = t[89] ^ t[90];
  assign t[62] = t[37] ^ t[91];
  assign t[63] = t[92] ^ t[93];
  assign t[64] = t[94] & t[95];
  assign t[65] = t[7] ? t[96] : t[184];
  assign t[66] = t[97] & t[98];
  assign t[67] = t[99] ? x[47] : x[46];
  assign t[68] = t[100] & t[101];
  assign t[69] = t[102] & t[103];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[104] ^ t[45]);
  assign t[71] = t[42] ^ t[103];
  assign t[72] = ~(t[74] & t[105]);
  assign t[73] = ~(t[185] ^ t[106]);
  assign t[74] = ~(t[107] & t[108]);
  assign t[75] = ~(t[186]);
  assign t[76] = t[27] ? x[55] : x[54];
  assign t[77] = t[180] ^ t[109];
  assign t[78] = t[26] ? t[110] : t[187];
  assign t[79] = t[181] ^ t[111];
  assign t[7] = ~(t[14]);
  assign t[80] = t[182] ^ t[112];
  assign t[81] = t[183] ^ t[113];
  assign t[82] = ~(t[88]);
  assign t[83] = ~(t[114]);
  assign t[84] = ~(t[36]);
  assign t[85] = t[115];
  assign t[86] = t[20] ^ t[114];
  assign t[87] = t[114] ^ t[37];
  assign t[88] = t[85] ^ t[36];
  assign t[89] = t[53] ^ t[33];
  assign t[8] = t[171] ^ t[15];
  assign t[90] = t[116] ^ t[117];
  assign t[91] = t[38] ^ t[118];
  assign t[92] = t[119] ? t[120] : t[188];
  assign t[93] = t[119] ? t[121] : t[189];
  assign t[94] = ~(t[63] ^ t[122]);
  assign t[95] = t[123] ^ t[124];
  assign t[96] = t[184] ^ t[125];
  assign t[97] = ~(t[68] ^ t[126]);
  assign t[98] = t[127] ^ t[128];
  assign t[99] = ~(t[129]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind102(x, y);
 input [116:0] x;
 output y;

 wire [225:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[7]);
  assign t[101] = t[134] ? x[68] : x[67];
  assign t[102] = t[134] ? x[70] : x[69];
  assign t[103] = t[135] & t[136];
  assign t[104] = t[137] & t[70];
  assign t[105] = t[65] ? t[138] : t[193];
  assign t[106] = t[185] ^ t[139];
  assign t[107] = t[186] ^ t[140];
  assign t[108] = t[187] ^ t[141];
  assign t[109] = ~(t[115]);
  assign t[10] = ~(t[19] ^ t[20]);
  assign t[110] = ~(t[91]);
  assign t[111] = ~(t[43]);
  assign t[112] = t[189] ^ t[142];
  assign t[113] = t[23] ^ t[91];
  assign t[114] = t[91] ^ t[44];
  assign t[115] = t[112] ^ t[43];
  assign t[116] = t[86] ? x[75] : x[74];
  assign t[117] = ~(t[143]);
  assign t[118] = ~(t[128]);
  assign t[119] = ~(t[129]);
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[144];
  assign t[121] = t[129] ^ t[25];
  assign t[122] = ~(t[173]);
  assign t[123] = t[190] ^ t[145];
  assign t[124] = t[96] ? t[146] : t[194];
  assign t[125] = t[191] ^ t[147];
  assign t[126] = t[192] ^ t[148];
  assign t[127] = t[149] & t[150];
  assign t[128] = t[151];
  assign t[129] = ~t[152];
  assign t[12] = t[23] ^ t[24];
  assign t[130] = t[153] ? x[80] : x[79];
  assign t[131] = t[154] & t[155];
  assign t[132] = ~(t[156] ^ t[98]);
  assign t[133] = t[157] ^ t[90];
  assign t[134] = ~(t[54]);
  assign t[135] = ~(t[158]);
  assign t[136] = ~(t[39]);
  assign t[137] = ~(t[40]);
  assign t[138] = t[193] ^ t[159];
  assign t[139] = t[134] ? x[82] : x[81];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[30] ? x[84] : x[83];
  assign t[141] = t[30] ? x[86] : x[85];
  assign t[142] = t[65] ? t[160] : t[195];
  assign t[143] = t[120] ^ t[129];
  assign t[144] = t[65] ? t[161] : t[196];
  assign t[145] = t[153] ? x[94] : x[93];
  assign t[146] = t[194] ^ t[162];
  assign t[147] = t[153] ? x[96] : x[95];
  assign t[148] = t[30] ? x[98] : x[97];
  assign t[149] = ~(t[103] ^ t[163]);
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[164] ^ t[158];
  assign t[151] = t[65] ? t[165] : t[197];
  assign t[152] = t[65] ? t[166] : t[198];
  assign t[153] = ~(t[54]);
  assign t[154] = ~(t[167]);
  assign t[155] = ~(t[88]);
  assign t[156] = t[88] ^ t[124];
  assign t[157] = t[124] ^ t[63];
  assign t[158] = t[70] ^ t[40];
  assign t[159] = t[86] ? x[106] : x[105];
  assign t[15] = t[173] | t[29];
  assign t[160] = t[195] ^ t[168];
  assign t[161] = t[196] ^ t[169];
  assign t[162] = t[153] ? x[108] : x[107];
  assign t[163] = t[69] ^ t[39];
  assign t[164] = t[39] ^ t[105];
  assign t[165] = t[197] ^ t[170];
  assign t[166] = t[198] ^ t[171];
  assign t[167] = t[90] ^ t[124];
  assign t[168] = t[30] ? x[110] : x[109];
  assign t[169] = t[86] ? x[112] : x[111];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[86] ? x[114] : x[113];
  assign t[171] = t[30] ? x[116] : x[115];
  assign t[172] = t[199] ^ x[4];
  assign t[173] = t[200] ^ x[7];
  assign t[174] = t[201] ^ x[12];
  assign t[175] = t[202] ^ x[15];
  assign t[176] = t[203] ^ x[18];
  assign t[177] = t[204] ^ x[21];
  assign t[178] = t[205] ^ x[24];
  assign t[179] = t[206] ^ x[27];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[207] ^ x[30];
  assign t[181] = t[208] ^ x[33];
  assign t[182] = t[209] ^ x[36];
  assign t[183] = t[210] ^ x[39];
  assign t[184] = t[211] ^ x[42];
  assign t[185] = t[212] ^ x[45];
  assign t[186] = t[213] ^ x[48];
  assign t[187] = t[214] ^ x[51];
  assign t[188] = t[215] ^ x[54];
  assign t[189] = t[216] ^ x[57];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[217] ^ x[60];
  assign t[191] = t[218] ^ x[63];
  assign t[192] = t[219] ^ x[66];
  assign t[193] = t[220] ^ x[73];
  assign t[194] = t[221] ^ x[78];
  assign t[195] = t[222] ^ x[89];
  assign t[196] = t[223] ^ x[92];
  assign t[197] = t[224] ^ x[101];
  assign t[198] = t[225] ^ x[104];
  assign t[199] = (x[2] & x[3]);
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[5] & x[6]);
  assign t[201] = (x[10] & x[11]);
  assign t[202] = (x[13] & x[14]);
  assign t[203] = (x[16] & x[17]);
  assign t[204] = (x[19] & x[20]);
  assign t[205] = (x[22] & x[23]);
  assign t[206] = (x[25] & x[26]);
  assign t[207] = (x[28] & x[29]);
  assign t[208] = (x[31] & x[32]);
  assign t[209] = (x[34] & x[35]);
  assign t[20] = ~(t[37] ^ t[38]);
  assign t[210] = (x[37] & x[38]);
  assign t[211] = (x[40] & x[41]);
  assign t[212] = (x[43] & x[44]);
  assign t[213] = (x[46] & x[47]);
  assign t[214] = (x[49] & x[50]);
  assign t[215] = (x[52] & x[53]);
  assign t[216] = (x[55] & x[56]);
  assign t[217] = (x[58] & x[59]);
  assign t[218] = (x[61] & x[62]);
  assign t[219] = (x[64] & x[65]);
  assign t[21] = t[39] ^ t[40];
  assign t[220] = (x[71] & x[72]);
  assign t[221] = (x[76] & x[77]);
  assign t[222] = (x[87] & x[88]);
  assign t[223] = (x[90] & x[91]);
  assign t[224] = (x[99] & x[100]);
  assign t[225] = (x[102] & x[103]);
  assign t[22] = t[41] & t[42];
  assign t[23] = t[43] ^ t[44];
  assign t[24] = t[45] ^ t[46];
  assign t[25] = t[47];
  assign t[26] = t[48] ^ t[49];
  assign t[27] = ~(t[29] & t[50]);
  assign t[28] = ~(t[174] ^ t[51]);
  assign t[29] = ~(t[52] & t[53]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[54]);
  assign t[31] = ~(t[175]);
  assign t[32] = ~(t[176]);
  assign t[33] = ~(t[177]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = t[57] ^ t[58];
  assign t[36] = t[59] ^ t[60];
  assign t[37] = t[61] ^ t[62];
  assign t[38] = t[63] ^ t[64];
  assign t[39] = t[65] ? t[66] : t[178];
  assign t[3] = t[7] ? t[8] : t[172];
  assign t[40] = t[65] ? t[67] : t[179];
  assign t[41] = ~(t[21] ^ t[68]);
  assign t[42] = t[69] ^ t[70];
  assign t[43] = t[177] ^ t[71];
  assign t[44] = t[180] ^ t[72];
  assign t[45] = t[73] ^ t[74];
  assign t[46] = t[75] & t[76];
  assign t[47] = t[65] ? t[77] : t[181];
  assign t[48] = t[78] ^ t[79];
  assign t[49] = t[80] & t[81];
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[82] & t[83]);
  assign t[51] = t[84] ^ t[182];
  assign t[52] = ~(t[174]);
  assign t[53] = t[85] & t[84];
  assign t[54] = ~(t[86]);
  assign t[55] = ~(t[180]);
  assign t[56] = ~(t[87] & t[183]);
  assign t[57] = t[88] ^ t[63];
  assign t[58] = t[89] & t[90];
  assign t[59] = t[91] ^ t[43];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[92] & t[93];
  assign t[61] = t[69] ^ t[94];
  assign t[62] = t[95] ^ t[49];
  assign t[63] = t[96] ? t[97] : t[184];
  assign t[64] = t[98] ^ t[99];
  assign t[65] = ~(t[100]);
  assign t[66] = t[178] ^ t[101];
  assign t[67] = t[179] ^ t[102];
  assign t[68] = t[103] ^ t[104];
  assign t[69] = t[40] ^ t[105];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[65] ? t[106] : t[185];
  assign t[71] = t[65] ? t[107] : t[186];
  assign t[72] = t[65] ? t[108] : t[187];
  assign t[73] = t[109] & t[110];
  assign t[74] = t[111] & t[112];
  assign t[75] = ~(t[73] ^ t[113]);
  assign t[76] = t[114] ^ t[115];
  assign t[77] = t[181] ^ t[116];
  assign t[78] = t[117] & t[118];
  assign t[79] = t[119] & t[120];
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[95] ^ t[48]);
  assign t[81] = t[121] ^ t[120];
  assign t[82] = ~(t[85] | t[84]);
  assign t[83] = ~(t[122] | t[52]);
  assign t[84] = ~(t[188]);
  assign t[85] = ~(t[182]);
  assign t[86] = ~(t[15]);
  assign t[87] = ~(t[189]);
  assign t[88] = t[96] ? t[123] : t[190];
  assign t[89] = ~(t[124]);
  assign t[8] = t[172] ^ t[16];
  assign t[90] = t[96] ? t[125] : t[191];
  assign t[91] = t[65] ? t[126] : t[192];
  assign t[92] = ~(t[59] ^ t[45]);
  assign t[93] = t[23] ^ t[112];
  assign t[94] = t[68] ^ t[127];
  assign t[95] = t[128] ^ t[129];
  assign t[96] = ~(t[100]);
  assign t[97] = t[184] ^ t[130];
  assign t[98] = t[131] ^ t[58];
  assign t[99] = t[132] & t[133];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind103(x, y);
 input [116:0] x;
 output y;

 wire [234:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[194] ^ t[128];
  assign t[101] = t[127] ? x[63] : x[62];
  assign t[102] = t[64] ? t[129] : t[199];
  assign t[103] = t[130] & t[131];
  assign t[104] = ~(t[103] ^ t[132]);
  assign t[105] = t[60] ^ t[133];
  assign t[106] = t[134] & t[135];
  assign t[107] = ~(t[116] ^ t[72]);
  assign t[108] = t[136] ^ t[42];
  assign t[109] = t[137] ? x[68] : x[67];
  assign t[10] = ~(t[19] ^ t[20]);
  assign t[110] = t[195] ^ t[138];
  assign t[111] = t[139] & t[140];
  assign t[112] = t[64] ? t[141] : t[200];
  assign t[113] = ~(t[182]);
  assign t[114] = t[64] ? t[142] : t[201];
  assign t[115] = ~(t[47]);
  assign t[116] = t[39] ^ t[67];
  assign t[117] = t[143] ? t[144] : t[202];
  assign t[118] = t[120] ^ t[145];
  assign t[119] = t[143] ? t[146] : t[203];
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[147] ^ t[148];
  assign t[121] = t[149] & t[150];
  assign t[122] = t[64] ? t[151] : t[204];
  assign t[123] = t[64] ? t[152] : t[205];
  assign t[124] = t[198] ^ t[153];
  assign t[125] = ~(t[154] ^ t[70]);
  assign t[126] = t[43] ^ t[94];
  assign t[127] = ~(t[155]);
  assign t[128] = t[127] ? x[88] : x[87];
  assign t[129] = t[199] ^ t[156];
  assign t[12] = t[23] ^ t[24];
  assign t[130] = ~(t[133]);
  assign t[131] = ~(t[92]);
  assign t[132] = t[43] ^ t[92];
  assign t[133] = t[94] ^ t[69];
  assign t[134] = ~(t[157]);
  assign t[135] = ~(t[39]);
  assign t[136] = t[67] ^ t[40];
  assign t[137] = ~(t[155]);
  assign t[138] = t[137] ? x[90] : x[89];
  assign t[139] = ~(t[158]);
  assign t[13] = t[25] ^ t[26];
  assign t[140] = ~(t[46]);
  assign t[141] = t[200] ^ t[159];
  assign t[142] = t[201] ^ t[160];
  assign t[143] = ~(t[97]);
  assign t[144] = t[202] ^ t[161];
  assign t[145] = t[162] & t[163];
  assign t[146] = t[203] ^ t[164];
  assign t[147] = t[165] & t[166];
  assign t[148] = t[167] & t[168];
  assign t[149] = ~(t[147] ^ t[169]);
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[170] ^ t[171];
  assign t[151] = t[204] ^ t[172];
  assign t[152] = t[205] ^ t[173];
  assign t[153] = t[30] ? x[92] : x[91];
  assign t[154] = t[92] ^ t[69];
  assign t[155] = ~(t[30]);
  assign t[156] = t[137] ? x[94] : x[93];
  assign t[157] = t[42] ^ t[67];
  assign t[158] = t[78] ^ t[47];
  assign t[159] = t[137] ? x[96] : x[95];
  assign t[15] = t[182] | t[29];
  assign t[160] = t[137] ? x[98] : x[97];
  assign t[161] = t[174] ? x[100] : x[99];
  assign t[162] = ~(t[175] ^ t[120]);
  assign t[163] = t[90] ^ t[168];
  assign t[164] = t[174] ? x[102] : x[101];
  assign t[165] = ~(t[171]);
  assign t[166] = ~(t[176]);
  assign t[167] = ~(t[119]);
  assign t[168] = t[143] ? t[177] : t[206];
  assign t[169] = t[90] ^ t[176];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[176] ^ t[117];
  assign t[171] = t[168] ^ t[119];
  assign t[172] = t[30] ? x[107] : x[106];
  assign t[173] = t[30] ? x[109] : x[108];
  assign t[174] = ~(t[155]);
  assign t[175] = t[176] ^ t[119];
  assign t[176] = t[143] ? t[178] : t[207];
  assign t[177] = t[206] ^ t[179];
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[174] ? x[114] : x[113];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[174] ? x[116] : x[115];
  assign t[181] = t[208] ^ x[4];
  assign t[182] = t[209] ^ x[7];
  assign t[183] = t[210] ^ x[12];
  assign t[184] = t[211] ^ x[15];
  assign t[185] = t[212] ^ x[18];
  assign t[186] = t[213] ^ x[21];
  assign t[187] = t[214] ^ x[24];
  assign t[188] = t[215] ^ x[27];
  assign t[189] = t[216] ^ x[30];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[217] ^ x[33];
  assign t[191] = t[218] ^ x[36];
  assign t[192] = t[219] ^ x[39];
  assign t[193] = t[220] ^ x[42];
  assign t[194] = t[221] ^ x[45];
  assign t[195] = t[222] ^ x[48];
  assign t[196] = t[223] ^ x[51];
  assign t[197] = t[224] ^ x[54];
  assign t[198] = t[225] ^ x[57];
  assign t[199] = t[226] ^ x[66];
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[71];
  assign t[201] = t[228] ^ x[74];
  assign t[202] = t[229] ^ x[77];
  assign t[203] = t[230] ^ x[80];
  assign t[204] = t[231] ^ x[83];
  assign t[205] = t[232] ^ x[86];
  assign t[206] = t[233] ^ x[105];
  assign t[207] = t[234] ^ x[112];
  assign t[208] = (x[2] & x[3]);
  assign t[209] = (x[5] & x[6]);
  assign t[20] = ~(t[37] ^ t[38]);
  assign t[210] = (x[10] & x[11]);
  assign t[211] = (x[13] & x[14]);
  assign t[212] = (x[16] & x[17]);
  assign t[213] = (x[19] & x[20]);
  assign t[214] = (x[22] & x[23]);
  assign t[215] = (x[25] & x[26]);
  assign t[216] = (x[28] & x[29]);
  assign t[217] = (x[31] & x[32]);
  assign t[218] = (x[34] & x[35]);
  assign t[219] = (x[37] & x[38]);
  assign t[21] = t[39] ^ t[40];
  assign t[220] = (x[40] & x[41]);
  assign t[221] = (x[43] & x[44]);
  assign t[222] = (x[46] & x[47]);
  assign t[223] = (x[49] & x[50]);
  assign t[224] = (x[52] & x[53]);
  assign t[225] = (x[55] & x[56]);
  assign t[226] = (x[64] & x[65]);
  assign t[227] = (x[69] & x[70]);
  assign t[228] = (x[72] & x[73]);
  assign t[229] = (x[75] & x[76]);
  assign t[22] = t[41] & t[42];
  assign t[230] = (x[78] & x[79]);
  assign t[231] = (x[81] & x[82]);
  assign t[232] = (x[84] & x[85]);
  assign t[233] = (x[103] & x[104]);
  assign t[234] = (x[110] & x[111]);
  assign t[23] = t[43] ^ t[44];
  assign t[24] = t[40] ^ t[45];
  assign t[25] = t[46] ^ t[47];
  assign t[26] = t[48] & t[49];
  assign t[27] = ~(t[29] & t[50]);
  assign t[28] = ~(t[183] ^ t[51]);
  assign t[29] = ~(t[52] & t[53]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[15]);
  assign t[31] = ~(t[184]);
  assign t[32] = ~(t[185]);
  assign t[33] = ~(t[186]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = t[56] ^ t[57];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[62] ^ t[63];
  assign t[39] = t[64] ? t[65] : t[187];
  assign t[3] = t[7] ? t[8] : t[181];
  assign t[40] = t[64] ? t[66] : t[188];
  assign t[41] = ~(t[67]);
  assign t[42] = t[64] ? t[68] : t[189];
  assign t[43] = t[69] ^ t[62];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[64] ? t[74] : t[190];
  assign t[47] = t[186] ^ t[75];
  assign t[48] = ~(t[25] ^ t[76]);
  assign t[49] = t[77] ^ t[78];
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[79] & t[80]);
  assign t[51] = t[81] ^ t[191];
  assign t[52] = ~(t[183]);
  assign t[53] = t[82] & t[81];
  assign t[54] = ~(t[192]);
  assign t[55] = ~(t[83] & t[193]);
  assign t[56] = t[84] ^ t[85];
  assign t[57] = t[86] ^ t[87];
  assign t[58] = ~(t[88] ^ t[89]);
  assign t[59] = t[90] ^ t[91];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[92] ^ t[62];
  assign t[61] = t[93] & t[94];
  assign t[62] = t[95];
  assign t[63] = t[70] ^ t[96];
  assign t[64] = ~(t[97]);
  assign t[65] = t[187] ^ t[98];
  assign t[66] = t[188] ^ t[99];
  assign t[67] = t[64] ? t[100] : t[194];
  assign t[68] = t[189] ^ t[101];
  assign t[69] = ~t[102];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[103] ^ t[61];
  assign t[71] = t[104] & t[105];
  assign t[72] = t[106] ^ t[22];
  assign t[73] = t[107] & t[108];
  assign t[74] = t[190] ^ t[109];
  assign t[75] = t[64] ? t[110] : t[195];
  assign t[76] = t[111] ^ t[87];
  assign t[77] = t[47] ^ t[84];
  assign t[78] = t[196] ^ t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[113] | t[52]);
  assign t[81] = ~(t[197]);
  assign t[82] = ~(t[191]);
  assign t[83] = ~(t[196]);
  assign t[84] = t[192] ^ t[114];
  assign t[85] = t[76] ^ t[26];
  assign t[86] = t[46] ^ t[84];
  assign t[87] = t[115] & t[78];
  assign t[88] = t[116] ^ t[73];
  assign t[89] = t[117] ^ t[118];
  assign t[8] = t[181] ^ t[16];
  assign t[90] = t[119] ^ t[117];
  assign t[91] = t[120] ^ t[121];
  assign t[92] = t[122];
  assign t[93] = ~(t[69]);
  assign t[94] = t[123];
  assign t[95] = t[64] ? t[124] : t[198];
  assign t[96] = t[125] & t[126];
  assign t[97] = ~(t[7]);
  assign t[98] = t[127] ? x[59] : x[58];
  assign t[99] = t[30] ? x[61] : x[60];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind104(x, y);
 input [116:0] x;
 output y;

 wire [245:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~t[125];
  assign t[101] = ~(t[69] ^ t[126]);
  assign t[102] = t[127] ^ t[128];
  assign t[103] = t[127] ^ t[129];
  assign t[104] = t[130] ^ t[131];
  assign t[105] = t[132] & t[133];
  assign t[106] = t[134] & t[135];
  assign t[107] = t[131] ^ t[136];
  assign t[108] = t[137] ^ t[138];
  assign t[109] = t[139] ^ t[41];
  assign t[10] = t[19] ^ t[20];
  assign t[110] = t[140];
  assign t[111] = t[126] ^ t[70];
  assign t[112] = ~(t[193]);
  assign t[113] = t[40] ^ t[62];
  assign t[114] = t[207] ^ t[141];
  assign t[115] = t[30] ? x[62] : x[61];
  assign t[116] = ~(t[142]);
  assign t[117] = ~(t[139]);
  assign t[118] = ~(t[97]);
  assign t[119] = t[56] ? t[143] : t[209];
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[139] ^ t[97];
  assign t[121] = t[208] ^ t[144];
  assign t[122] = ~(t[93] ^ t[145]);
  assign t[123] = t[109] ^ t[142];
  assign t[124] = t[56] ? t[146] : t[210];
  assign t[125] = t[56] ? t[147] : t[211];
  assign t[126] = t[148] ^ t[149];
  assign t[127] = t[100] ^ t[110];
  assign t[128] = t[150];
  assign t[129] = t[126] ^ t[151];
  assign t[12] = ~(t[23] ^ t[24]);
  assign t[130] = t[152] ? t[153] : t[212];
  assign t[131] = t[152] ? t[154] : t[213];
  assign t[132] = ~(t[104] ^ t[137]);
  assign t[133] = t[107] ^ t[155];
  assign t[134] = ~(t[58] ^ t[156]);
  assign t[135] = t[21] ^ t[113];
  assign t[136] = t[152] ? t[157] : t[214];
  assign t[137] = t[158] ^ t[159];
  assign t[138] = t[160] & t[161];
  assign t[139] = t[56] ? t[162] : t[215];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[56] ? t[163] : t[216];
  assign t[141] = t[30] ? x[88] : x[87];
  assign t[142] = t[119] ^ t[97];
  assign t[143] = t[209] ^ t[164];
  assign t[144] = t[165] ? x[90] : x[89];
  assign t[145] = t[67] ^ t[139];
  assign t[146] = t[210] ^ t[166];
  assign t[147] = t[211] ^ t[167];
  assign t[148] = t[168] & t[169];
  assign t[149] = t[170] & t[128];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[56] ? t[171] : t[217];
  assign t[151] = t[172] & t[173];
  assign t[152] = ~(t[84]);
  assign t[153] = t[212] ^ t[174];
  assign t[154] = t[213] ^ t[175];
  assign t[155] = t[152] ? t[176] : t[218];
  assign t[156] = t[73] ^ t[38];
  assign t[157] = t[214] ^ t[177];
  assign t[158] = t[178] & t[179];
  assign t[159] = t[180] & t[155];
  assign t[15] = t[193] | t[29];
  assign t[160] = ~(t[158] ^ t[181]);
  assign t[161] = t[182] ^ t[183];
  assign t[162] = t[215] ^ t[184];
  assign t[163] = t[216] ^ t[185];
  assign t[164] = t[165] ? x[98] : x[97];
  assign t[165] = ~(t[53]);
  assign t[166] = t[82] ? x[100] : x[99];
  assign t[167] = t[30] ? x[102] : x[101];
  assign t[168] = ~(t[186]);
  assign t[169] = ~(t[99]);
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = ~(t[100]);
  assign t[171] = t[217] ^ t[187];
  assign t[172] = ~(t[148] ^ t[188]);
  assign t[173] = t[189] ^ t[186];
  assign t[174] = t[190] ? x[104] : x[103];
  assign t[175] = t[190] ? x[106] : x[105];
  assign t[176] = t[218] ^ t[191];
  assign t[177] = t[190] ? x[108] : x[107];
  assign t[178] = ~(t[183]);
  assign t[179] = ~(t[130]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = ~(t[131]);
  assign t[181] = t[107] ^ t[130];
  assign t[182] = t[130] ^ t[136];
  assign t[183] = t[155] ^ t[131];
  assign t[184] = t[165] ? x[110] : x[109];
  assign t[185] = t[82] ? x[112] : x[111];
  assign t[186] = t[128] ^ t[100];
  assign t[187] = t[82] ? x[114] : x[113];
  assign t[188] = t[127] ^ t[99];
  assign t[189] = t[99] ^ t[110];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = ~(t[53]);
  assign t[191] = t[190] ? x[116] : x[115];
  assign t[192] = t[219] ^ x[4];
  assign t[193] = t[220] ^ x[7];
  assign t[194] = t[221] ^ x[12];
  assign t[195] = t[222] ^ x[15];
  assign t[196] = t[223] ^ x[18];
  assign t[197] = t[224] ^ x[21];
  assign t[198] = t[225] ^ x[24];
  assign t[199] = t[226] ^ x[27];
  assign t[19] = t[194] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[30];
  assign t[201] = t[228] ^ x[33];
  assign t[202] = t[229] ^ x[36];
  assign t[203] = t[230] ^ x[39];
  assign t[204] = t[231] ^ x[42];
  assign t[205] = t[232] ^ x[45];
  assign t[206] = t[233] ^ x[48];
  assign t[207] = t[234] ^ x[55];
  assign t[208] = t[235] ^ x[60];
  assign t[209] = t[236] ^ x[65];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[68];
  assign t[211] = t[238] ^ x[71];
  assign t[212] = t[239] ^ x[74];
  assign t[213] = t[240] ^ x[77];
  assign t[214] = t[241] ^ x[80];
  assign t[215] = t[242] ^ x[83];
  assign t[216] = t[243] ^ x[86];
  assign t[217] = t[244] ^ x[93];
  assign t[218] = t[245] ^ x[96];
  assign t[219] = (x[2] & x[3]);
  assign t[21] = t[38] ^ t[19];
  assign t[220] = (x[5] & x[6]);
  assign t[221] = (x[10] & x[11]);
  assign t[222] = (x[13] & x[14]);
  assign t[223] = (x[16] & x[17]);
  assign t[224] = (x[19] & x[20]);
  assign t[225] = (x[22] & x[23]);
  assign t[226] = (x[25] & x[26]);
  assign t[227] = (x[28] & x[29]);
  assign t[228] = (x[31] & x[32]);
  assign t[229] = (x[34] & x[35]);
  assign t[22] = t[39] & t[40];
  assign t[230] = (x[37] & x[38]);
  assign t[231] = (x[40] & x[41]);
  assign t[232] = (x[43] & x[44]);
  assign t[233] = (x[46] & x[47]);
  assign t[234] = (x[53] & x[54]);
  assign t[235] = (x[58] & x[59]);
  assign t[236] = (x[63] & x[64]);
  assign t[237] = (x[66] & x[67]);
  assign t[238] = (x[69] & x[70]);
  assign t[239] = (x[72] & x[73]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (x[75] & x[76]);
  assign t[241] = (x[78] & x[79]);
  assign t[242] = (x[81] & x[82]);
  assign t[243] = (x[84] & x[85]);
  assign t[244] = (x[91] & x[92]);
  assign t[245] = (x[94] & x[95]);
  assign t[24] = t[43] ^ t[44];
  assign t[25] = ~(t[45] ^ t[46]);
  assign t[26] = ~(t[47] ^ t[48]);
  assign t[27] = ~(t[29] & t[49]);
  assign t[28] = ~(t[195] ^ t[50]);
  assign t[29] = ~(t[51] & t[52]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = ~(t[53]);
  assign t[31] = ~(t[196]);
  assign t[32] = ~(t[197]);
  assign t[33] = ~(t[198]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = t[56] ? t[57] : t[199];
  assign t[36] = t[58] ^ t[22];
  assign t[37] = t[59] & t[60];
  assign t[38] = t[56] ? t[61] : t[200];
  assign t[39] = ~(t[62]);
  assign t[3] = t[7] ? t[8] : t[192];
  assign t[40] = t[201] ^ t[63];
  assign t[41] = t[56] ? t[64] : t[202];
  assign t[42] = t[65] ^ t[66];
  assign t[43] = t[67] ^ t[68];
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[71] ^ t[72]);
  assign t[46] = t[73] ^ t[74];
  assign t[47] = t[75] ^ t[76];
  assign t[48] = ~(t[10] ^ t[77]);
  assign t[49] = ~(t[78] & t[79]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[80] ^ t[203];
  assign t[51] = ~(t[195]);
  assign t[52] = t[81] & t[80];
  assign t[53] = ~(t[82]);
  assign t[54] = ~(t[194]);
  assign t[55] = ~(t[83] & t[204]);
  assign t[56] = ~(t[84]);
  assign t[57] = t[199] ^ t[85];
  assign t[58] = t[86] & t[87];
  assign t[59] = ~(t[88] ^ t[36]);
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[73] ^ t[40];
  assign t[61] = t[200] ^ t[89];
  assign t[62] = t[198] ^ t[90];
  assign t[63] = t[56] ? t[91] : t[205];
  assign t[64] = t[202] ^ t[92];
  assign t[65] = t[93] ^ t[94];
  assign t[66] = t[95] & t[96];
  assign t[67] = t[97] ^ t[41];
  assign t[68] = t[65] ^ t[98];
  assign t[69] = t[99] ^ t[100];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[101] & t[102];
  assign t[71] = t[103] ^ t[23];
  assign t[72] = t[104] ^ t[105];
  assign t[73] = t[62] ^ t[19];
  assign t[74] = t[36] ^ t[106];
  assign t[75] = t[107] ^ t[108];
  assign t[76] = t[109] ^ t[94];
  assign t[77] = t[110] ^ t[111];
  assign t[78] = ~(t[81] | t[80]);
  assign t[79] = ~(t[112] | t[51]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[206]);
  assign t[81] = ~(t[203]);
  assign t[82] = ~(t[15]);
  assign t[83] = ~(t[201]);
  assign t[84] = ~(t[7]);
  assign t[85] = t[30] ? x[50] : x[49];
  assign t[86] = ~(t[113]);
  assign t[87] = ~(t[38]);
  assign t[88] = t[38] ^ t[62];
  assign t[89] = t[30] ? x[52] : x[51];
  assign t[8] = t[192] ^ t[16];
  assign t[90] = t[56] ? t[114] : t[207];
  assign t[91] = t[205] ^ t[115];
  assign t[92] = t[82] ? x[57] : x[56];
  assign t[93] = t[116] & t[117];
  assign t[94] = t[118] & t[119];
  assign t[95] = ~(t[120] ^ t[65]);
  assign t[96] = t[67] ^ t[119];
  assign t[97] = t[56] ? t[121] : t[208];
  assign t[98] = t[122] & t[123];
  assign t[99] = t[124];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind105(x, y);
 input [116:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[124] ? t[125] : t[190];
  assign t[101] = t[124] ? t[126] : t[191];
  assign t[102] = ~(t[69] ^ t[127]);
  assign t[103] = t[128] ^ t[129];
  assign t[104] = t[60] ? t[130] : t[192];
  assign t[105] = ~(t[74] ^ t[131]);
  assign t[106] = t[132] ^ t[133];
  assign t[107] = t[134] ? x[75] : x[74];
  assign t[108] = ~(t[133]);
  assign t[109] = ~(t[135]);
  assign t[10] = t[19] ^ t[20];
  assign t[110] = ~(t[71]);
  assign t[111] = t[187] ^ t[136];
  assign t[112] = t[135] ^ t[71];
  assign t[113] = ~(t[172]);
  assign t[114] = t[30] ? x[77] : x[76];
  assign t[115] = t[30] ? x[79] : x[78];
  assign t[116] = t[188] ^ t[137];
  assign t[117] = t[30] ? x[81] : x[80];
  assign t[118] = ~(t[138]);
  assign t[119] = t[60] ? t[139] : t[193];
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[189] ^ t[140];
  assign t[121] = t[141] ^ t[20];
  assign t[122] = t[142] & t[143];
  assign t[123] = t[144] & t[145];
  assign t[124] = ~(t[87]);
  assign t[125] = t[190] ^ t[146];
  assign t[126] = t[191] ^ t[147];
  assign t[127] = t[148] ^ t[149];
  assign t[128] = t[101] ^ t[150];
  assign t[129] = t[124] ? t[151] : t[194];
  assign t[12] = ~(t[23] ^ t[24]);
  assign t[130] = t[192] ^ t[152];
  assign t[131] = t[45] ^ t[135];
  assign t[132] = t[135] ^ t[25];
  assign t[133] = t[111] ^ t[71];
  assign t[134] = ~(t[138]);
  assign t[135] = t[60] ? t[153] : t[195];
  assign t[136] = t[60] ? t[154] : t[196];
  assign t[137] = t[134] ? x[95] : x[94];
  assign t[138] = ~(t[30]);
  assign t[139] = t[193] ^ t[155];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[118] ? x[97] : x[96];
  assign t[141] = t[156] & t[157];
  assign t[142] = ~(t[141] ^ t[158]);
  assign t[143] = t[19] ^ t[159];
  assign t[144] = ~(t[160] ^ t[41]);
  assign t[145] = t[21] ^ t[93];
  assign t[146] = t[161] ? x[99] : x[98];
  assign t[147] = t[161] ? x[101] : x[100];
  assign t[148] = t[162] & t[163];
  assign t[149] = t[164] & t[129];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[124] ? t[165] : t[197];
  assign t[151] = t[194] ^ t[166];
  assign t[152] = t[134] ? x[106] : x[105];
  assign t[153] = t[195] ^ t[167];
  assign t[154] = t[196] ^ t[168];
  assign t[155] = t[118] ? x[108] : x[107];
  assign t[156] = ~(t[159]);
  assign t[157] = ~(t[35]);
  assign t[158] = t[97] ^ t[35];
  assign t[159] = t[38] ^ t[58];
  assign t[15] = t[172] | t[29];
  assign t[160] = t[119] ^ t[39];
  assign t[161] = ~(t[138]);
  assign t[162] = ~(t[169]);
  assign t[163] = ~(t[100]);
  assign t[164] = ~(t[101]);
  assign t[165] = t[197] ^ t[170];
  assign t[166] = t[161] ? x[110] : x[109];
  assign t[167] = t[134] ? x[112] : x[111];
  assign t[168] = t[134] ? x[114] : x[113];
  assign t[169] = t[129] ^ t[101];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[161] ? x[116] : x[115];
  assign t[171] = t[198] ^ x[4];
  assign t[172] = t[199] ^ x[7];
  assign t[173] = t[200] ^ x[12];
  assign t[174] = t[201] ^ x[15];
  assign t[175] = t[202] ^ x[18];
  assign t[176] = t[203] ^ x[21];
  assign t[177] = t[204] ^ x[24];
  assign t[178] = t[205] ^ x[27];
  assign t[179] = t[206] ^ x[30];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[207] ^ x[33];
  assign t[181] = t[208] ^ x[36];
  assign t[182] = t[209] ^ x[39];
  assign t[183] = t[210] ^ x[42];
  assign t[184] = t[211] ^ x[45];
  assign t[185] = t[212] ^ x[48];
  assign t[186] = t[213] ^ x[51];
  assign t[187] = t[214] ^ x[54];
  assign t[188] = t[215] ^ x[57];
  assign t[189] = t[216] ^ x[64];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[217] ^ x[67];
  assign t[191] = t[218] ^ x[70];
  assign t[192] = t[219] ^ x[73];
  assign t[193] = t[220] ^ x[84];
  assign t[194] = t[221] ^ x[87];
  assign t[195] = t[222] ^ x[90];
  assign t[196] = t[223] ^ x[93];
  assign t[197] = t[224] ^ x[104];
  assign t[198] = (x[2] & x[3]);
  assign t[199] = (x[5] & x[6]);
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[10] & x[11]);
  assign t[201] = (x[13] & x[14]);
  assign t[202] = (x[16] & x[17]);
  assign t[203] = (x[19] & x[20]);
  assign t[204] = (x[22] & x[23]);
  assign t[205] = (x[25] & x[26]);
  assign t[206] = (x[28] & x[29]);
  assign t[207] = (x[31] & x[32]);
  assign t[208] = (x[34] & x[35]);
  assign t[209] = (x[37] & x[38]);
  assign t[20] = t[37] & t[38];
  assign t[210] = (x[40] & x[41]);
  assign t[211] = (x[43] & x[44]);
  assign t[212] = (x[46] & x[47]);
  assign t[213] = (x[49] & x[50]);
  assign t[214] = (x[52] & x[53]);
  assign t[215] = (x[55] & x[56]);
  assign t[216] = (x[62] & x[63]);
  assign t[217] = (x[65] & x[66]);
  assign t[218] = (x[68] & x[69]);
  assign t[219] = (x[71] & x[72]);
  assign t[21] = t[39] ^ t[40];
  assign t[220] = (x[82] & x[83]);
  assign t[221] = (x[85] & x[86]);
  assign t[222] = (x[88] & x[89]);
  assign t[223] = (x[91] & x[92]);
  assign t[224] = (x[102] & x[103]);
  assign t[22] = t[41] ^ t[42];
  assign t[23] = ~(t[43] ^ t[44]);
  assign t[24] = t[45] ^ t[46];
  assign t[25] = t[173] ^ t[47];
  assign t[26] = t[48] ^ t[49];
  assign t[27] = ~(t[29] & t[50]);
  assign t[28] = ~(t[174] ^ t[51]);
  assign t[29] = ~(t[52] & t[53]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[15]);
  assign t[31] = ~(t[175]);
  assign t[32] = ~(t[176]);
  assign t[33] = ~(t[177]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = t[56];
  assign t[36] = t[57];
  assign t[37] = ~(t[58]);
  assign t[38] = t[59];
  assign t[39] = t[60] ? t[61] : t[178];
  assign t[3] = t[7] ? t[8] : t[171];
  assign t[40] = t[60] ? t[62] : t[179];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[67] ^ t[68];
  assign t[44] = t[69] ^ t[70];
  assign t[45] = t[71] ^ t[25];
  assign t[46] = t[48] ^ t[72];
  assign t[47] = t[60] ? t[73] : t[180];
  assign t[48] = t[74] ^ t[75];
  assign t[49] = t[76] & t[77];
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[78] & t[79]);
  assign t[51] = t[80] ^ t[181];
  assign t[52] = ~(t[174]);
  assign t[53] = t[81] & t[80];
  assign t[54] = ~(t[173]);
  assign t[55] = ~(t[82] & t[182]);
  assign t[56] = t[60] ? t[83] : t[183];
  assign t[57] = t[60] ? t[84] : t[184];
  assign t[58] = ~t[85];
  assign t[59] = t[60] ? t[86] : t[185];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = ~(t[87]);
  assign t[61] = t[178] ^ t[88];
  assign t[62] = t[179] ^ t[89];
  assign t[63] = t[90] & t[91];
  assign t[64] = t[92] & t[93];
  assign t[65] = ~(t[63] ^ t[94]);
  assign t[66] = t[95] ^ t[96];
  assign t[67] = t[97] ^ t[98];
  assign t[68] = t[40] ^ t[99];
  assign t[69] = t[100] ^ t[101];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[102] & t[103];
  assign t[71] = t[177] ^ t[104];
  assign t[72] = t[105] & t[106];
  assign t[73] = t[180] ^ t[107];
  assign t[74] = t[108] & t[109];
  assign t[75] = t[110] & t[111];
  assign t[76] = ~(t[112] ^ t[48]);
  assign t[77] = t[45] ^ t[111];
  assign t[78] = ~(t[81] | t[80]);
  assign t[79] = ~(t[113] | t[52]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[186]);
  assign t[81] = ~(t[181]);
  assign t[82] = ~(t[187]);
  assign t[83] = t[183] ^ t[114];
  assign t[84] = t[184] ^ t[115];
  assign t[85] = t[60] ? t[116] : t[188];
  assign t[86] = t[185] ^ t[117];
  assign t[87] = ~(t[7]);
  assign t[88] = t[118] ? x[59] : x[58];
  assign t[89] = t[30] ? x[61] : x[60];
  assign t[8] = t[171] ^ t[16];
  assign t[90] = ~(t[96]);
  assign t[91] = ~(t[119]);
  assign t[92] = ~(t[39]);
  assign t[93] = t[60] ? t[120] : t[189];
  assign t[94] = t[21] ^ t[119];
  assign t[95] = t[119] ^ t[40];
  assign t[96] = t[93] ^ t[39];
  assign t[97] = t[58] ^ t[36];
  assign t[98] = t[121] ^ t[122];
  assign t[99] = t[41] ^ t[123];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind106(x, y);
 input [116:0] x;
 output y;

 wire [225:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[30] ? x[64] : x[63];
  assign t[101] = t[30] ? x[66] : x[65];
  assign t[102] = t[134] & t[135];
  assign t[103] = t[136] & t[70];
  assign t[104] = t[7] ? t[137] : t[191];
  assign t[105] = t[184] ^ t[138];
  assign t[106] = t[185] ^ t[139];
  assign t[107] = t[186] ^ t[140];
  assign t[108] = ~(t[114]);
  assign t[109] = ~(t[92]);
  assign t[10] = ~(t[19] ^ t[20]);
  assign t[110] = ~(t[43]);
  assign t[111] = t[141];
  assign t[112] = t[23] ^ t[92];
  assign t[113] = t[92] ^ t[44];
  assign t[114] = t[111] ^ t[43];
  assign t[115] = ~(t[55]);
  assign t[116] = ~(t[142]);
  assign t[117] = ~(t[128]);
  assign t[118] = ~(t[129]);
  assign t[119] = t[47] ? t[143] : t[192];
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[129] ^ t[25];
  assign t[121] = ~(t[173]);
  assign t[122] = ~(t[77]);
  assign t[123] = t[189] ^ t[144];
  assign t[124] = t[176] ^ t[145];
  assign t[125] = t[122] ? t[146] : t[193];
  assign t[126] = t[47] ? t[147] : t[194];
  assign t[127] = t[148] & t[149];
  assign t[128] = t[47] ? t[150] : t[195];
  assign t[129] = t[47] ? t[151] : t[196];
  assign t[12] = t[23] ^ t[24];
  assign t[130] = t[190] ^ t[152];
  assign t[131] = t[153] & t[154];
  assign t[132] = ~(t[155] ^ t[98]);
  assign t[133] = t[156] ^ t[91];
  assign t[134] = ~(t[157]);
  assign t[135] = ~(t[39]);
  assign t[136] = ~(t[40]);
  assign t[137] = t[191] ^ t[158];
  assign t[138] = t[87] ? x[86] : x[85];
  assign t[139] = t[115] ? x[88] : x[87];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[115] ? x[90] : x[89];
  assign t[141] = t[7] ? t[159] : t[197];
  assign t[142] = t[119] ^ t[129];
  assign t[143] = t[192] ^ t[160];
  assign t[144] = t[161] ? x[95] : x[94];
  assign t[145] = t[122] ? t[162] : t[198];
  assign t[146] = t[193] ^ t[163];
  assign t[147] = t[194] ^ t[164];
  assign t[148] = ~(t[102] ^ t[165]);
  assign t[149] = t[166] ^ t[157];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[195] ^ t[167];
  assign t[151] = t[196] ^ t[168];
  assign t[152] = t[161] ? x[100] : x[99];
  assign t[153] = ~(t[169]);
  assign t[154] = ~(t[89]);
  assign t[155] = t[89] ^ t[124];
  assign t[156] = t[124] ^ t[64];
  assign t[157] = t[70] ^ t[40];
  assign t[158] = t[87] ? x[102] : x[101];
  assign t[159] = t[197] ^ t[170];
  assign t[15] = t[173] | t[29];
  assign t[160] = t[115] ? x[104] : x[103];
  assign t[161] = ~(t[55]);
  assign t[162] = t[198] ^ t[171];
  assign t[163] = t[161] ? x[106] : x[105];
  assign t[164] = t[115] ? x[108] : x[107];
  assign t[165] = t[69] ^ t[39];
  assign t[166] = t[39] ^ t[104];
  assign t[167] = t[115] ? x[110] : x[109];
  assign t[168] = t[115] ? x[112] : x[111];
  assign t[169] = t[91] ^ t[124];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[115] ? x[114] : x[113];
  assign t[171] = t[161] ? x[116] : x[115];
  assign t[172] = t[199] ^ x[4];
  assign t[173] = t[200] ^ x[7];
  assign t[174] = t[201] ^ x[12];
  assign t[175] = t[202] ^ x[15];
  assign t[176] = t[203] ^ x[18];
  assign t[177] = t[204] ^ x[21];
  assign t[178] = t[205] ^ x[24];
  assign t[179] = t[206] ^ x[27];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[207] ^ x[30];
  assign t[181] = t[208] ^ x[33];
  assign t[182] = t[209] ^ x[36];
  assign t[183] = t[210] ^ x[39];
  assign t[184] = t[211] ^ x[42];
  assign t[185] = t[212] ^ x[45];
  assign t[186] = t[213] ^ x[48];
  assign t[187] = t[214] ^ x[53];
  assign t[188] = t[215] ^ x[56];
  assign t[189] = t[216] ^ x[59];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[217] ^ x[62];
  assign t[191] = t[218] ^ x[69];
  assign t[192] = t[219] ^ x[72];
  assign t[193] = t[220] ^ x[75];
  assign t[194] = t[221] ^ x[78];
  assign t[195] = t[222] ^ x[81];
  assign t[196] = t[223] ^ x[84];
  assign t[197] = t[224] ^ x[93];
  assign t[198] = t[225] ^ x[98];
  assign t[199] = (x[2] & x[3]);
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[5] & x[6]);
  assign t[201] = (x[10] & x[11]);
  assign t[202] = (x[13] & x[14]);
  assign t[203] = (x[16] & x[17]);
  assign t[204] = (x[19] & x[20]);
  assign t[205] = (x[22] & x[23]);
  assign t[206] = (x[25] & x[26]);
  assign t[207] = (x[28] & x[29]);
  assign t[208] = (x[31] & x[32]);
  assign t[209] = (x[34] & x[35]);
  assign t[20] = ~(t[37] ^ t[38]);
  assign t[210] = (x[37] & x[38]);
  assign t[211] = (x[40] & x[41]);
  assign t[212] = (x[43] & x[44]);
  assign t[213] = (x[46] & x[47]);
  assign t[214] = (x[51] & x[52]);
  assign t[215] = (x[54] & x[55]);
  assign t[216] = (x[57] & x[58]);
  assign t[217] = (x[60] & x[61]);
  assign t[218] = (x[67] & x[68]);
  assign t[219] = (x[70] & x[71]);
  assign t[21] = t[39] ^ t[40];
  assign t[220] = (x[73] & x[74]);
  assign t[221] = (x[76] & x[77]);
  assign t[222] = (x[79] & x[80]);
  assign t[223] = (x[82] & x[83]);
  assign t[224] = (x[91] & x[92]);
  assign t[225] = (x[96] & x[97]);
  assign t[22] = t[41] & t[42];
  assign t[23] = t[43] ^ t[44];
  assign t[24] = t[45] ^ t[46];
  assign t[25] = t[47] ? t[48] : t[174];
  assign t[26] = t[49] ^ t[50];
  assign t[27] = ~(t[29] & t[51]);
  assign t[28] = ~(t[175] ^ t[52]);
  assign t[29] = ~(t[53] & t[54]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[55]);
  assign t[31] = ~(t[176]);
  assign t[32] = ~(t[177]);
  assign t[33] = ~(t[178]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = t[58] ^ t[59];
  assign t[36] = t[60] ^ t[61];
  assign t[37] = t[62] ^ t[63];
  assign t[38] = t[64] ^ t[65];
  assign t[39] = t[7] ? t[66] : t[179];
  assign t[3] = t[7] ? t[8] : t[172];
  assign t[40] = t[7] ? t[67] : t[180];
  assign t[41] = ~(t[21] ^ t[68]);
  assign t[42] = t[69] ^ t[70];
  assign t[43] = ~t[71];
  assign t[44] = ~t[72];
  assign t[45] = t[73] ^ t[74];
  assign t[46] = t[75] & t[76];
  assign t[47] = ~(t[77]);
  assign t[48] = t[174] ^ t[78];
  assign t[49] = t[79] ^ t[80];
  assign t[4] = ~(t[9]);
  assign t[50] = t[81] & t[82];
  assign t[51] = ~(t[83] & t[84]);
  assign t[52] = t[85] ^ t[181];
  assign t[53] = ~(t[175]);
  assign t[54] = t[86] & t[85];
  assign t[55] = ~(t[87]);
  assign t[56] = ~(t[182]);
  assign t[57] = ~(t[88] & t[183]);
  assign t[58] = t[89] ^ t[64];
  assign t[59] = t[90] & t[91];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[92] ^ t[43];
  assign t[61] = t[93] & t[94];
  assign t[62] = t[69] ^ t[95];
  assign t[63] = t[96] ^ t[50];
  assign t[64] = t[183] ^ t[97];
  assign t[65] = t[98] ^ t[99];
  assign t[66] = t[179] ^ t[100];
  assign t[67] = t[180] ^ t[101];
  assign t[68] = t[102] ^ t[103];
  assign t[69] = t[40] ^ t[104];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[7] ? t[105] : t[184];
  assign t[71] = t[47] ? t[106] : t[185];
  assign t[72] = t[47] ? t[107] : t[186];
  assign t[73] = t[108] & t[109];
  assign t[74] = t[110] & t[111];
  assign t[75] = ~(t[73] ^ t[112]);
  assign t[76] = t[113] ^ t[114];
  assign t[77] = ~(t[7]);
  assign t[78] = t[115] ? x[50] : x[49];
  assign t[79] = t[116] & t[117];
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = t[118] & t[119];
  assign t[81] = ~(t[96] ^ t[49]);
  assign t[82] = t[120] ^ t[119];
  assign t[83] = ~(t[86] | t[85]);
  assign t[84] = ~(t[121] | t[53]);
  assign t[85] = ~(t[187]);
  assign t[86] = ~(t[181]);
  assign t[87] = ~(t[15]);
  assign t[88] = ~(t[188]);
  assign t[89] = t[122] ? t[123] : t[189];
  assign t[8] = t[172] ^ t[16];
  assign t[90] = ~(t[124]);
  assign t[91] = t[177] ^ t[125];
  assign t[92] = t[126];
  assign t[93] = ~(t[60] ^ t[45]);
  assign t[94] = t[23] ^ t[111];
  assign t[95] = t[68] ^ t[127];
  assign t[96] = t[128] ^ t[129];
  assign t[97] = t[122] ? t[130] : t[190];
  assign t[98] = t[131] ^ t[59];
  assign t[99] = t[132] & t[133];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind107(x, y);
 input [116:0] x;
 output y;

 wire [234:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[30] ? x[72] : x[71];
  assign t[101] = t[195] ^ t[129];
  assign t[102] = t[130] & t[131];
  assign t[103] = ~(t[102] ^ t[132]);
  assign t[104] = t[60] ^ t[133];
  assign t[105] = t[134] & t[135];
  assign t[106] = ~(t[115] ^ t[71]);
  assign t[107] = t[136] ^ t[42];
  assign t[108] = t[196] ^ t[137];
  assign t[109] = t[197] ^ t[138];
  assign t[10] = ~(t[19] ^ t[20]);
  assign t[110] = t[139] & t[140];
  assign t[111] = t[7] ? t[141] : t[202];
  assign t[112] = ~(t[182]);
  assign t[113] = t[94] ? t[142] : t[203];
  assign t[114] = ~(t[47]);
  assign t[115] = t[39] ^ t[66];
  assign t[116] = t[192] ^ t[143];
  assign t[117] = t[119] ^ t[144];
  assign t[118] = t[184] ^ t[145];
  assign t[119] = t[146] ^ t[147];
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[148] & t[149];
  assign t[121] = t[200] ^ t[150];
  assign t[122] = t[201] ^ t[151];
  assign t[123] = ~(t[7]);
  assign t[124] = t[152] ? x[80] : x[79];
  assign t[125] = ~(t[153] ^ t[69]);
  assign t[126] = t[43] ^ t[93];
  assign t[127] = ~(t[154]);
  assign t[128] = t[127] ? x[82] : x[81];
  assign t[129] = t[152] ? x[84] : x[83];
  assign t[12] = t[23] ^ t[24];
  assign t[130] = ~(t[133]);
  assign t[131] = ~(t[91]);
  assign t[132] = t[43] ^ t[91];
  assign t[133] = t[93] ^ t[68];
  assign t[134] = ~(t[155]);
  assign t[135] = ~(t[39]);
  assign t[136] = t[66] ^ t[40];
  assign t[137] = t[152] ? x[86] : x[85];
  assign t[138] = t[152] ? x[88] : x[87];
  assign t[139] = ~(t[156]);
  assign t[13] = t[25] ^ t[26];
  assign t[140] = ~(t[46]);
  assign t[141] = t[202] ^ t[157];
  assign t[142] = t[203] ^ t[158];
  assign t[143] = t[159] ? t[160] : t[204];
  assign t[144] = t[161] & t[162];
  assign t[145] = t[159] ? t[163] : t[205];
  assign t[146] = t[164] & t[165];
  assign t[147] = t[166] & t[167];
  assign t[148] = ~(t[146] ^ t[168]);
  assign t[149] = t[169] ^ t[170];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[152] ? x[96] : x[95];
  assign t[151] = t[152] ? x[98] : x[97];
  assign t[152] = ~(t[154]);
  assign t[153] = t[91] ^ t[68];
  assign t[154] = ~(t[30]);
  assign t[155] = t[42] ^ t[66];
  assign t[156] = t[77] ^ t[47];
  assign t[157] = t[152] ? x[100] : x[99];
  assign t[158] = t[152] ? x[102] : x[101];
  assign t[159] = ~(t[123]);
  assign t[15] = t[182] | t[29];
  assign t[160] = t[204] ^ t[171];
  assign t[161] = ~(t[172] ^ t[119]);
  assign t[162] = t[89] ^ t[167];
  assign t[163] = t[205] ^ t[173];
  assign t[164] = ~(t[170]);
  assign t[165] = ~(t[174]);
  assign t[166] = ~(t[118]);
  assign t[167] = t[185] ^ t[175];
  assign t[168] = t[89] ^ t[174];
  assign t[169] = t[174] ^ t[116];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[167] ^ t[118];
  assign t[171] = t[176] ? x[104] : x[103];
  assign t[172] = t[174] ^ t[118];
  assign t[173] = t[176] ? x[106] : x[105];
  assign t[174] = t[159] ? t[177] : t[206];
  assign t[175] = t[159] ? t[178] : t[207];
  assign t[176] = ~(t[154]);
  assign t[177] = t[206] ^ t[179];
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[176] ? x[114] : x[113];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[176] ? x[116] : x[115];
  assign t[181] = t[208] ^ x[4];
  assign t[182] = t[209] ^ x[7];
  assign t[183] = t[210] ^ x[12];
  assign t[184] = t[211] ^ x[15];
  assign t[185] = t[212] ^ x[18];
  assign t[186] = t[213] ^ x[21];
  assign t[187] = t[214] ^ x[24];
  assign t[188] = t[215] ^ x[27];
  assign t[189] = t[216] ^ x[30];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[217] ^ x[33];
  assign t[191] = t[218] ^ x[36];
  assign t[192] = t[219] ^ x[39];
  assign t[193] = t[220] ^ x[42];
  assign t[194] = t[221] ^ x[45];
  assign t[195] = t[222] ^ x[48];
  assign t[196] = t[223] ^ x[51];
  assign t[197] = t[224] ^ x[54];
  assign t[198] = t[225] ^ x[57];
  assign t[199] = t[226] ^ x[60];
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[63];
  assign t[201] = t[228] ^ x[66];
  assign t[202] = t[229] ^ x[75];
  assign t[203] = t[230] ^ x[78];
  assign t[204] = t[231] ^ x[91];
  assign t[205] = t[232] ^ x[94];
  assign t[206] = t[233] ^ x[109];
  assign t[207] = t[234] ^ x[112];
  assign t[208] = (x[2] & x[3]);
  assign t[209] = (x[5] & x[6]);
  assign t[20] = ~(t[37] ^ t[38]);
  assign t[210] = (x[10] & x[11]);
  assign t[211] = (x[13] & x[14]);
  assign t[212] = (x[16] & x[17]);
  assign t[213] = (x[19] & x[20]);
  assign t[214] = (x[22] & x[23]);
  assign t[215] = (x[25] & x[26]);
  assign t[216] = (x[28] & x[29]);
  assign t[217] = (x[31] & x[32]);
  assign t[218] = (x[34] & x[35]);
  assign t[219] = (x[37] & x[38]);
  assign t[21] = t[39] ^ t[40];
  assign t[220] = (x[40] & x[41]);
  assign t[221] = (x[43] & x[44]);
  assign t[222] = (x[46] & x[47]);
  assign t[223] = (x[49] & x[50]);
  assign t[224] = (x[52] & x[53]);
  assign t[225] = (x[55] & x[56]);
  assign t[226] = (x[58] & x[59]);
  assign t[227] = (x[61] & x[62]);
  assign t[228] = (x[64] & x[65]);
  assign t[229] = (x[73] & x[74]);
  assign t[22] = t[41] & t[42];
  assign t[230] = (x[76] & x[77]);
  assign t[231] = (x[89] & x[90]);
  assign t[232] = (x[92] & x[93]);
  assign t[233] = (x[107] & x[108]);
  assign t[234] = (x[110] & x[111]);
  assign t[23] = t[43] ^ t[44];
  assign t[24] = t[40] ^ t[45];
  assign t[25] = t[46] ^ t[47];
  assign t[26] = t[48] & t[49];
  assign t[27] = ~(t[29] & t[50]);
  assign t[28] = ~(t[183] ^ t[51]);
  assign t[29] = ~(t[52] & t[53]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[15]);
  assign t[31] = ~(t[184]);
  assign t[32] = ~(t[185]);
  assign t[33] = ~(t[186]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = t[56] ^ t[57];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[62] ^ t[63];
  assign t[39] = t[7] ? t[64] : t[187];
  assign t[3] = t[7] ? t[8] : t[181];
  assign t[40] = t[7] ? t[65] : t[188];
  assign t[41] = ~(t[66]);
  assign t[42] = t[7] ? t[67] : t[189];
  assign t[43] = t[68] ^ t[62];
  assign t[44] = t[69] ^ t[70];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = t[73];
  assign t[47] = ~t[74];
  assign t[48] = ~(t[25] ^ t[75]);
  assign t[49] = t[76] ^ t[77];
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[78] & t[79]);
  assign t[51] = t[80] ^ t[190];
  assign t[52] = ~(t[183]);
  assign t[53] = t[81] & t[80];
  assign t[54] = ~(t[191]);
  assign t[55] = ~(t[82] & t[192]);
  assign t[56] = t[83] ^ t[84];
  assign t[57] = t[85] ^ t[86];
  assign t[58] = ~(t[87] ^ t[88]);
  assign t[59] = t[89] ^ t[90];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[91] ^ t[62];
  assign t[61] = t[92] & t[93];
  assign t[62] = t[94] ? t[95] : t[193];
  assign t[63] = t[69] ^ t[96];
  assign t[64] = t[187] ^ t[97];
  assign t[65] = t[188] ^ t[98];
  assign t[66] = t[7] ? t[99] : t[194];
  assign t[67] = t[189] ^ t[100];
  assign t[68] = t[94] ? t[101] : t[195];
  assign t[69] = t[102] ^ t[61];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[103] & t[104];
  assign t[71] = t[105] ^ t[22];
  assign t[72] = t[106] & t[107];
  assign t[73] = t[94] ? t[108] : t[196];
  assign t[74] = t[94] ? t[109] : t[197];
  assign t[75] = t[110] ^ t[86];
  assign t[76] = t[47] ^ t[83];
  assign t[77] = t[111];
  assign t[78] = ~(t[81] | t[80]);
  assign t[79] = ~(t[112] | t[52]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[198]);
  assign t[81] = ~(t[190]);
  assign t[82] = ~(t[199]);
  assign t[83] = ~t[113];
  assign t[84] = t[75] ^ t[26];
  assign t[85] = t[46] ^ t[83];
  assign t[86] = t[114] & t[77];
  assign t[87] = t[115] ^ t[72];
  assign t[88] = t[116] ^ t[117];
  assign t[89] = t[118] ^ t[116];
  assign t[8] = t[181] ^ t[16];
  assign t[90] = t[119] ^ t[120];
  assign t[91] = t[94] ? t[121] : t[200];
  assign t[92] = ~(t[68]);
  assign t[93] = t[94] ? t[122] : t[201];
  assign t[94] = ~(t[123]);
  assign t[95] = t[193] ^ t[124];
  assign t[96] = t[125] & t[126];
  assign t[97] = t[127] ? x[68] : x[67];
  assign t[98] = t[30] ? x[70] : x[69];
  assign t[99] = t[194] ^ t[128];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind108(x, y);
 input [116:0] x;
 output y;

 wire [245:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[56] ? t[127] : t[210];
  assign t[101] = ~(t[69] ^ t[128]);
  assign t[102] = t[129] ^ t[130];
  assign t[103] = t[129] ^ t[131];
  assign t[104] = t[132] ^ t[133];
  assign t[105] = t[134] & t[135];
  assign t[106] = t[136] & t[137];
  assign t[107] = t[133] ^ t[138];
  assign t[108] = t[139] ^ t[140];
  assign t[109] = t[141] ^ t[41];
  assign t[10] = t[19] ^ t[20];
  assign t[110] = t[56] ? t[142] : t[211];
  assign t[111] = t[128] ^ t[70];
  assign t[112] = ~(t[193]);
  assign t[113] = ~(t[53]);
  assign t[114] = t[40] ^ t[62];
  assign t[115] = t[113] ? x[69] : x[68];
  assign t[116] = t[207] ^ t[143];
  assign t[117] = t[113] ? x[71] : x[70];
  assign t[118] = ~(t[144]);
  assign t[119] = ~(t[141]);
  assign t[11] = t[21] ^ t[22];
  assign t[120] = ~(t[97]);
  assign t[121] = t[7] ? t[145] : t[212];
  assign t[122] = t[141] ^ t[97];
  assign t[123] = t[208] ^ t[146];
  assign t[124] = ~(t[93] ^ t[147]);
  assign t[125] = t[109] ^ t[144];
  assign t[126] = t[209] ^ t[148];
  assign t[127] = t[210] ^ t[149];
  assign t[128] = t[150] ^ t[151];
  assign t[129] = t[100] ^ t[110];
  assign t[12] = ~(t[23] ^ t[24]);
  assign t[130] = t[56] ? t[152] : t[213];
  assign t[131] = t[128] ^ t[153];
  assign t[132] = t[154] ? t[155] : t[214];
  assign t[133] = t[195] ^ t[156];
  assign t[134] = ~(t[104] ^ t[139]);
  assign t[135] = t[107] ^ t[157];
  assign t[136] = ~(t[58] ^ t[158]);
  assign t[137] = t[21] ^ t[114];
  assign t[138] = t[202] ^ t[159];
  assign t[139] = t[160] ^ t[161];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[162] & t[163];
  assign t[141] = t[7] ? t[164] : t[215];
  assign t[142] = t[211] ^ t[165];
  assign t[143] = t[113] ? x[85] : x[84];
  assign t[144] = t[121] ^ t[97];
  assign t[145] = t[212] ^ t[166];
  assign t[146] = t[30] ? x[87] : x[86];
  assign t[147] = t[67] ^ t[141];
  assign t[148] = t[113] ? x[89] : x[88];
  assign t[149] = t[113] ? x[91] : x[90];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[167] & t[168];
  assign t[151] = t[169] & t[130];
  assign t[152] = t[213] ^ t[170];
  assign t[153] = t[171] & t[172];
  assign t[154] = ~(t[84]);
  assign t[155] = t[214] ^ t[173];
  assign t[156] = t[154] ? t[174] : t[216];
  assign t[157] = t[196] ^ t[175];
  assign t[158] = t[73] ^ t[38];
  assign t[159] = t[154] ? t[176] : t[217];
  assign t[15] = t[193] | t[29];
  assign t[160] = t[177] & t[178];
  assign t[161] = t[179] & t[157];
  assign t[162] = ~(t[160] ^ t[180]);
  assign t[163] = t[181] ^ t[182];
  assign t[164] = t[215] ^ t[183];
  assign t[165] = t[113] ? x[99] : x[98];
  assign t[166] = t[82] ? x[101] : x[100];
  assign t[167] = ~(t[184]);
  assign t[168] = ~(t[99]);
  assign t[169] = ~(t[100]);
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[113] ? x[103] : x[102];
  assign t[171] = ~(t[150] ^ t[185]);
  assign t[172] = t[186] ^ t[184];
  assign t[173] = t[187] ? x[105] : x[104];
  assign t[174] = t[216] ^ t[188];
  assign t[175] = t[154] ? t[189] : t[218];
  assign t[176] = t[217] ^ t[190];
  assign t[177] = ~(t[182]);
  assign t[178] = ~(t[132]);
  assign t[179] = ~(t[133]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[107] ^ t[132];
  assign t[181] = t[132] ^ t[138];
  assign t[182] = t[157] ^ t[133];
  assign t[183] = t[30] ? x[110] : x[109];
  assign t[184] = t[130] ^ t[100];
  assign t[185] = t[129] ^ t[99];
  assign t[186] = t[99] ^ t[110];
  assign t[187] = ~(t[53]);
  assign t[188] = t[187] ? x[112] : x[111];
  assign t[189] = t[218] ^ t[191];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[187] ? x[114] : x[113];
  assign t[191] = t[187] ? x[116] : x[115];
  assign t[192] = t[219] ^ x[4];
  assign t[193] = t[220] ^ x[7];
  assign t[194] = t[221] ^ x[12];
  assign t[195] = t[222] ^ x[15];
  assign t[196] = t[223] ^ x[18];
  assign t[197] = t[224] ^ x[21];
  assign t[198] = t[225] ^ x[24];
  assign t[199] = t[226] ^ x[27];
  assign t[19] = ~t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[30];
  assign t[201] = t[228] ^ x[33];
  assign t[202] = t[229] ^ x[36];
  assign t[203] = t[230] ^ x[39];
  assign t[204] = t[231] ^ x[42];
  assign t[205] = t[232] ^ x[45];
  assign t[206] = t[233] ^ x[48];
  assign t[207] = t[234] ^ x[53];
  assign t[208] = t[235] ^ x[58];
  assign t[209] = t[236] ^ x[61];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[64];
  assign t[211] = t[238] ^ x[67];
  assign t[212] = t[239] ^ x[74];
  assign t[213] = t[240] ^ x[77];
  assign t[214] = t[241] ^ x[80];
  assign t[215] = t[242] ^ x[83];
  assign t[216] = t[243] ^ x[94];
  assign t[217] = t[244] ^ x[97];
  assign t[218] = t[245] ^ x[108];
  assign t[219] = (x[2] & x[3]);
  assign t[21] = t[38] ^ t[19];
  assign t[220] = (x[5] & x[6]);
  assign t[221] = (x[10] & x[11]);
  assign t[222] = (x[13] & x[14]);
  assign t[223] = (x[16] & x[17]);
  assign t[224] = (x[19] & x[20]);
  assign t[225] = (x[22] & x[23]);
  assign t[226] = (x[25] & x[26]);
  assign t[227] = (x[28] & x[29]);
  assign t[228] = (x[31] & x[32]);
  assign t[229] = (x[34] & x[35]);
  assign t[22] = t[39] & t[40];
  assign t[230] = (x[37] & x[38]);
  assign t[231] = (x[40] & x[41]);
  assign t[232] = (x[43] & x[44]);
  assign t[233] = (x[46] & x[47]);
  assign t[234] = (x[51] & x[52]);
  assign t[235] = (x[56] & x[57]);
  assign t[236] = (x[59] & x[60]);
  assign t[237] = (x[62] & x[63]);
  assign t[238] = (x[65] & x[66]);
  assign t[239] = (x[72] & x[73]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (x[75] & x[76]);
  assign t[241] = (x[78] & x[79]);
  assign t[242] = (x[81] & x[82]);
  assign t[243] = (x[92] & x[93]);
  assign t[244] = (x[95] & x[96]);
  assign t[245] = (x[106] & x[107]);
  assign t[24] = t[43] ^ t[44];
  assign t[25] = ~(t[45] ^ t[46]);
  assign t[26] = ~(t[47] ^ t[48]);
  assign t[27] = ~(t[29] & t[49]);
  assign t[28] = ~(t[194] ^ t[50]);
  assign t[29] = ~(t[51] & t[52]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = ~(t[53]);
  assign t[31] = ~(t[195]);
  assign t[32] = ~(t[196]);
  assign t[33] = ~(t[197]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = t[56] ? t[57] : t[198];
  assign t[36] = t[58] ^ t[22];
  assign t[37] = t[59] & t[60];
  assign t[38] = t[61];
  assign t[39] = ~(t[62]);
  assign t[3] = t[7] ? t[8] : t[192];
  assign t[40] = t[63];
  assign t[41] = t[7] ? t[64] : t[199];
  assign t[42] = t[65] ^ t[66];
  assign t[43] = t[67] ^ t[68];
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[71] ^ t[72]);
  assign t[46] = t[73] ^ t[74];
  assign t[47] = t[75] ^ t[76];
  assign t[48] = ~(t[10] ^ t[77]);
  assign t[49] = ~(t[78] & t[79]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[80] ^ t[200];
  assign t[51] = ~(t[194]);
  assign t[52] = t[81] & t[80];
  assign t[53] = ~(t[82]);
  assign t[54] = ~(t[201]);
  assign t[55] = ~(t[83] & t[202]);
  assign t[56] = ~(t[84]);
  assign t[57] = t[198] ^ t[85];
  assign t[58] = t[86] & t[87];
  assign t[59] = ~(t[88] ^ t[36]);
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[73] ^ t[40];
  assign t[61] = t[56] ? t[89] : t[203];
  assign t[62] = ~t[90];
  assign t[63] = t[7] ? t[91] : t[204];
  assign t[64] = t[199] ^ t[92];
  assign t[65] = t[93] ^ t[94];
  assign t[66] = t[95] & t[96];
  assign t[67] = t[97] ^ t[41];
  assign t[68] = t[65] ^ t[98];
  assign t[69] = t[99] ^ t[100];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[101] & t[102];
  assign t[71] = t[103] ^ t[23];
  assign t[72] = t[104] ^ t[105];
  assign t[73] = t[62] ^ t[19];
  assign t[74] = t[36] ^ t[106];
  assign t[75] = t[107] ^ t[108];
  assign t[76] = t[109] ^ t[94];
  assign t[77] = t[110] ^ t[111];
  assign t[78] = ~(t[81] | t[80]);
  assign t[79] = ~(t[112] | t[51]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[205]);
  assign t[81] = ~(t[200]);
  assign t[82] = ~(t[15]);
  assign t[83] = ~(t[206]);
  assign t[84] = ~(t[7]);
  assign t[85] = t[113] ? x[50] : x[49];
  assign t[86] = ~(t[114]);
  assign t[87] = ~(t[38]);
  assign t[88] = t[38] ^ t[62];
  assign t[89] = t[203] ^ t[115];
  assign t[8] = t[192] ^ t[16];
  assign t[90] = t[56] ? t[116] : t[207];
  assign t[91] = t[204] ^ t[117];
  assign t[92] = t[82] ? x[55] : x[54];
  assign t[93] = t[118] & t[119];
  assign t[94] = t[120] & t[121];
  assign t[95] = ~(t[122] ^ t[65]);
  assign t[96] = t[67] ^ t[121];
  assign t[97] = t[7] ? t[123] : t[208];
  assign t[98] = t[124] & t[125];
  assign t[99] = t[56] ? t[126] : t[209];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind109(x, y);
 input [116:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[70] ^ t[126]);
  assign t[101] = t[127] ^ t[128];
  assign t[102] = t[112] ? x[72] : x[71];
  assign t[103] = ~(t[128]);
  assign t[104] = ~(t[129]);
  assign t[105] = ~(t[67]);
  assign t[106] = t[130];
  assign t[107] = t[129] ^ t[67];
  assign t[108] = ~(t[131] & t[132]);
  assign t[109] = t[133] ^ t[190];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = ~(t[185]);
  assign t[111] = t[134] & t[133];
  assign t[112] = ~(t[49]);
  assign t[113] = t[112] ? x[77] : x[76];
  assign t[114] = ~(t[49]);
  assign t[115] = t[26] ? t[135] : t[191];
  assign t[116] = t[187] ^ t[136];
  assign t[117] = t[137] ^ t[19];
  assign t[118] = t[138] & t[139];
  assign t[119] = t[140] & t[141];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[188] ^ t[142];
  assign t[121] = t[7] ? t[143] : t[192];
  assign t[122] = t[144] ^ t[145];
  assign t[123] = t[96] ^ t[146];
  assign t[124] = t[173] ^ t[147];
  assign t[125] = t[189] ^ t[148];
  assign t[126] = t[42] ^ t[129];
  assign t[127] = t[129] ^ t[24];
  assign t[128] = t[106] ^ t[67];
  assign t[129] = t[149];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[26] ? t[150] : t[193];
  assign t[131] = ~(t[134] | t[133]);
  assign t[132] = ~(t[151] | t[110]);
  assign t[133] = ~(t[194]);
  assign t[134] = ~(t[190]);
  assign t[135] = t[191] ^ t[152];
  assign t[136] = t[77] ? x[91] : x[90];
  assign t[137] = t[153] & t[154];
  assign t[138] = ~(t[137] ^ t[155]);
  assign t[139] = t[18] ^ t[156];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[157] ^ t[38]);
  assign t[141] = t[20] ^ t[88];
  assign t[142] = t[27] ? x[93] : x[92];
  assign t[143] = t[192] ^ t[158];
  assign t[144] = t[159] & t[160];
  assign t[145] = t[161] & t[124];
  assign t[146] = t[183] ^ t[162];
  assign t[147] = t[7] ? t[163] : t[195];
  assign t[148] = t[112] ? x[98] : x[97];
  assign t[149] = t[52] ? t[164] : t[196];
  assign t[14] = ~(t[26]);
  assign t[150] = t[193] ^ t[165];
  assign t[151] = ~(t[181]);
  assign t[152] = t[114] ? x[103] : x[102];
  assign t[153] = ~(t[156]);
  assign t[154] = ~(t[32]);
  assign t[155] = t[92] ^ t[32];
  assign t[156] = t[35] ^ t[55];
  assign t[157] = t[115] ^ t[36];
  assign t[158] = t[27] ? x[105] : x[104];
  assign t[159] = ~(t[166]);
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = ~(t[95]);
  assign t[161] = ~(t[96]);
  assign t[162] = t[7] ? t[167] : t[197];
  assign t[163] = t[195] ^ t[168];
  assign t[164] = t[196] ^ t[169];
  assign t[165] = t[112] ? x[110] : x[109];
  assign t[166] = t[124] ^ t[96];
  assign t[167] = t[197] ^ t[170];
  assign t[168] = t[27] ? x[112] : x[111];
  assign t[169] = t[112] ? x[114] : x[113];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[27] ? x[116] : x[115];
  assign t[171] = t[198] ^ x[4];
  assign t[172] = t[199] ^ x[9];
  assign t[173] = t[200] ^ x[12];
  assign t[174] = t[201] ^ x[15];
  assign t[175] = t[202] ^ x[18];
  assign t[176] = t[203] ^ x[21];
  assign t[177] = t[204] ^ x[24];
  assign t[178] = t[205] ^ x[27];
  assign t[179] = t[206] ^ x[30];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[207] ^ x[33];
  assign t[181] = t[208] ^ x[36];
  assign t[182] = t[209] ^ x[39];
  assign t[183] = t[210] ^ x[42];
  assign t[184] = t[211] ^ x[45];
  assign t[185] = t[212] ^ x[48];
  assign t[186] = t[213] ^ x[51];
  assign t[187] = t[214] ^ x[64];
  assign t[188] = t[215] ^ x[67];
  assign t[189] = t[216] ^ x[70];
  assign t[18] = t[32] ^ t[33];
  assign t[190] = t[217] ^ x[75];
  assign t[191] = t[218] ^ x[80];
  assign t[192] = t[219] ^ x[83];
  assign t[193] = t[220] ^ x[86];
  assign t[194] = t[221] ^ x[89];
  assign t[195] = t[222] ^ x[96];
  assign t[196] = t[223] ^ x[101];
  assign t[197] = t[224] ^ x[108];
  assign t[198] = (x[2] & x[3]);
  assign t[199] = (x[7] & x[8]);
  assign t[19] = t[34] & t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[10] & x[11]);
  assign t[201] = (x[13] & x[14]);
  assign t[202] = (x[16] & x[17]);
  assign t[203] = (x[19] & x[20]);
  assign t[204] = (x[22] & x[23]);
  assign t[205] = (x[25] & x[26]);
  assign t[206] = (x[28] & x[29]);
  assign t[207] = (x[31] & x[32]);
  assign t[208] = (x[34] & x[35]);
  assign t[209] = (x[37] & x[38]);
  assign t[20] = t[36] ^ t[37];
  assign t[210] = (x[40] & x[41]);
  assign t[211] = (x[43] & x[44]);
  assign t[212] = (x[46] & x[47]);
  assign t[213] = (x[49] & x[50]);
  assign t[214] = (x[62] & x[63]);
  assign t[215] = (x[65] & x[66]);
  assign t[216] = (x[68] & x[69]);
  assign t[217] = (x[73] & x[74]);
  assign t[218] = (x[78] & x[79]);
  assign t[219] = (x[81] & x[82]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = (x[84] & x[85]);
  assign t[221] = (x[87] & x[88]);
  assign t[222] = (x[94] & x[95]);
  assign t[223] = (x[99] & x[100]);
  assign t[224] = (x[106] & x[107]);
  assign t[22] = ~(t[40] ^ t[41]);
  assign t[23] = t[42] ^ t[43];
  assign t[24] = ~t[44];
  assign t[25] = t[45] ^ t[46];
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49]);
  assign t[28] = ~(t[172]);
  assign t[29] = ~(t[173]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[174]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = t[52] ? t[53] : t[175];
  assign t[33] = t[52] ? t[54] : t[176];
  assign t[34] = ~(t[55]);
  assign t[35] = t[52] ? t[56] : t[177];
  assign t[36] = t[26] ? t[57] : t[178];
  assign t[37] = t[26] ? t[58] : t[179];
  assign t[38] = t[59] ^ t[60];
  assign t[39] = t[61] & t[62];
  assign t[3] = t[7] ? t[8] : t[171];
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] ^ t[24];
  assign t[43] = t[45] ^ t[68];
  assign t[44] = t[52] ? t[69] : t[180];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] & t[73];
  assign t[47] = ~(t[74] & t[75]);
  assign t[48] = t[181] | t[76];
  assign t[49] = ~(t[77]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[182]);
  assign t[51] = ~(t[78] & t[183]);
  assign t[52] = ~(t[14]);
  assign t[53] = t[175] ^ t[79];
  assign t[54] = t[176] ^ t[80];
  assign t[55] = t[52] ? t[81] : t[184];
  assign t[56] = t[177] ^ t[82];
  assign t[57] = t[178] ^ t[83];
  assign t[58] = t[179] ^ t[84];
  assign t[59] = t[85] & t[86];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[87] & t[88];
  assign t[61] = ~(t[59] ^ t[89]);
  assign t[62] = t[90] ^ t[91];
  assign t[63] = t[92] ^ t[93];
  assign t[64] = t[37] ^ t[94];
  assign t[65] = t[95] ^ t[96];
  assign t[66] = t[97] & t[98];
  assign t[67] = ~t[99];
  assign t[68] = t[100] & t[101];
  assign t[69] = t[180] ^ t[102];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[103] & t[104];
  assign t[71] = t[105] & t[106];
  assign t[72] = ~(t[107] ^ t[45]);
  assign t[73] = t[42] ^ t[106];
  assign t[74] = ~(t[76] & t[108]);
  assign t[75] = ~(t[185] ^ t[109]);
  assign t[76] = ~(t[110] & t[111]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[186]);
  assign t[79] = t[112] ? x[53] : x[52];
  assign t[7] = ~(t[14]);
  assign t[80] = t[112] ? x[55] : x[54];
  assign t[81] = t[184] ^ t[113];
  assign t[82] = t[112] ? x[57] : x[56];
  assign t[83] = t[114] ? x[59] : x[58];
  assign t[84] = t[77] ? x[61] : x[60];
  assign t[85] = ~(t[91]);
  assign t[86] = ~(t[115]);
  assign t[87] = ~(t[36]);
  assign t[88] = t[26] ? t[116] : t[187];
  assign t[89] = t[20] ^ t[115];
  assign t[8] = t[171] ^ t[15];
  assign t[90] = t[115] ^ t[37];
  assign t[91] = t[88] ^ t[36];
  assign t[92] = t[55] ^ t[33];
  assign t[93] = t[117] ^ t[118];
  assign t[94] = t[38] ^ t[119];
  assign t[95] = t[7] ? t[120] : t[188];
  assign t[96] = t[172] ^ t[121];
  assign t[97] = ~(t[65] ^ t[122]);
  assign t[98] = t[123] ^ t[124];
  assign t[99] = t[52] ? t[125] : t[189];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind110(x, y);
 input [116:0] x;
 output y;

 wire [225:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[133] & t[134];
  assign t[101] = t[135] & t[69];
  assign t[102] = t[183] ^ t[136];
  assign t[103] = t[7] ? t[137] : t[190];
  assign t[104] = t[131] ? x[66] : x[65];
  assign t[105] = t[131] ? x[68] : x[67];
  assign t[106] = ~(t[112]);
  assign t[107] = ~(t[90]);
  assign t[108] = ~(t[43]);
  assign t[109] = t[47] ? t[138] : t[191];
  assign t[10] = ~(t[19] ^ t[20]);
  assign t[110] = t[23] ^ t[90];
  assign t[111] = t[90] ^ t[44];
  assign t[112] = t[109] ^ t[43];
  assign t[113] = ~(t[139]);
  assign t[114] = ~(t[140]);
  assign t[115] = ~(t[125]);
  assign t[116] = ~(t[126]);
  assign t[117] = t[47] ? t[141] : t[192];
  assign t[118] = t[126] ^ t[25];
  assign t[119] = ~(t[173]);
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[7] ? t[142] : t[193];
  assign t[121] = t[143];
  assign t[122] = t[7] ? t[144] : t[194];
  assign t[123] = t[188] ^ t[145];
  assign t[124] = t[146] & t[147];
  assign t[125] = t[47] ? t[148] : t[195];
  assign t[126] = t[47] ? t[149] : t[196];
  assign t[127] = t[189] ^ t[150];
  assign t[128] = t[151] & t[152];
  assign t[129] = ~(t[153] ^ t[96]);
  assign t[12] = t[23] ^ t[24];
  assign t[130] = t[154] ^ t[89];
  assign t[131] = ~(t[139]);
  assign t[132] = t[131] ? x[88] : x[87];
  assign t[133] = ~(t[155]);
  assign t[134] = ~(t[39]);
  assign t[135] = ~(t[40]);
  assign t[136] = t[156] ? t[157] : t[197];
  assign t[137] = t[190] ^ t[158];
  assign t[138] = t[191] ^ t[159];
  assign t[139] = ~(t[30]);
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[117] ^ t[126];
  assign t[141] = t[192] ^ t[160];
  assign t[142] = t[193] ^ t[161];
  assign t[143] = t[7] ? t[162] : t[198];
  assign t[144] = t[194] ^ t[163];
  assign t[145] = t[131] ? x[96] : x[95];
  assign t[146] = ~(t[100] ^ t[164]);
  assign t[147] = t[165] ^ t[155];
  assign t[148] = t[195] ^ t[166];
  assign t[149] = t[196] ^ t[167];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[30] ? x[98] : x[97];
  assign t[151] = ~(t[168]);
  assign t[152] = ~(t[87]);
  assign t[153] = t[87] ^ t[121];
  assign t[154] = t[121] ^ t[63];
  assign t[155] = t[69] ^ t[40];
  assign t[156] = ~(t[76]);
  assign t[157] = t[197] ^ t[169];
  assign t[158] = t[30] ? x[100] : x[99];
  assign t[159] = t[131] ? x[102] : x[101];
  assign t[15] = t[173] | t[29];
  assign t[160] = t[113] ? x[104] : x[103];
  assign t[161] = t[30] ? x[106] : x[105];
  assign t[162] = t[198] ^ t[170];
  assign t[163] = t[171] ? x[108] : x[107];
  assign t[164] = t[68] ^ t[39];
  assign t[165] = t[39] ^ t[102];
  assign t[166] = t[113] ? x[110] : x[109];
  assign t[167] = t[113] ? x[112] : x[111];
  assign t[168] = t[89] ^ t[121];
  assign t[169] = t[171] ? x[114] : x[113];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[171] ? x[116] : x[115];
  assign t[171] = ~(t[139]);
  assign t[172] = t[199] ^ x[4];
  assign t[173] = t[200] ^ x[7];
  assign t[174] = t[201] ^ x[12];
  assign t[175] = t[202] ^ x[15];
  assign t[176] = t[203] ^ x[18];
  assign t[177] = t[204] ^ x[21];
  assign t[178] = t[205] ^ x[24];
  assign t[179] = t[206] ^ x[27];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[207] ^ x[30];
  assign t[181] = t[208] ^ x[33];
  assign t[182] = t[209] ^ x[36];
  assign t[183] = t[210] ^ x[39];
  assign t[184] = t[211] ^ x[42];
  assign t[185] = t[212] ^ x[45];
  assign t[186] = t[213] ^ x[48];
  assign t[187] = t[214] ^ x[53];
  assign t[188] = t[215] ^ x[56];
  assign t[189] = t[216] ^ x[59];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[217] ^ x[64];
  assign t[191] = t[218] ^ x[71];
  assign t[192] = t[219] ^ x[74];
  assign t[193] = t[220] ^ x[77];
  assign t[194] = t[221] ^ x[80];
  assign t[195] = t[222] ^ x[83];
  assign t[196] = t[223] ^ x[86];
  assign t[197] = t[224] ^ x[91];
  assign t[198] = t[225] ^ x[94];
  assign t[199] = (x[2] & x[3]);
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[5] & x[6]);
  assign t[201] = (x[10] & x[11]);
  assign t[202] = (x[13] & x[14]);
  assign t[203] = (x[16] & x[17]);
  assign t[204] = (x[19] & x[20]);
  assign t[205] = (x[22] & x[23]);
  assign t[206] = (x[25] & x[26]);
  assign t[207] = (x[28] & x[29]);
  assign t[208] = (x[31] & x[32]);
  assign t[209] = (x[34] & x[35]);
  assign t[20] = ~(t[37] ^ t[38]);
  assign t[210] = (x[37] & x[38]);
  assign t[211] = (x[40] & x[41]);
  assign t[212] = (x[43] & x[44]);
  assign t[213] = (x[46] & x[47]);
  assign t[214] = (x[51] & x[52]);
  assign t[215] = (x[54] & x[55]);
  assign t[216] = (x[57] & x[58]);
  assign t[217] = (x[62] & x[63]);
  assign t[218] = (x[69] & x[70]);
  assign t[219] = (x[72] & x[73]);
  assign t[21] = t[39] ^ t[40];
  assign t[220] = (x[75] & x[76]);
  assign t[221] = (x[78] & x[79]);
  assign t[222] = (x[81] & x[82]);
  assign t[223] = (x[84] & x[85]);
  assign t[224] = (x[89] & x[90]);
  assign t[225] = (x[92] & x[93]);
  assign t[22] = t[41] & t[42];
  assign t[23] = t[43] ^ t[44];
  assign t[24] = t[45] ^ t[46];
  assign t[25] = t[47] ? t[48] : t[174];
  assign t[26] = t[49] ^ t[50];
  assign t[27] = ~(t[29] & t[51]);
  assign t[28] = ~(t[175] ^ t[52]);
  assign t[29] = ~(t[53] & t[54]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[15]);
  assign t[31] = ~(t[176]);
  assign t[32] = ~(t[177]);
  assign t[33] = ~(t[178]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = t[57] ^ t[58];
  assign t[36] = t[59] ^ t[60];
  assign t[37] = t[61] ^ t[62];
  assign t[38] = t[63] ^ t[64];
  assign t[39] = t[7] ? t[65] : t[179];
  assign t[3] = t[7] ? t[8] : t[172];
  assign t[40] = t[178] ^ t[66];
  assign t[41] = ~(t[21] ^ t[67]);
  assign t[42] = t[68] ^ t[69];
  assign t[43] = t[47] ? t[70] : t[180];
  assign t[44] = t[47] ? t[71] : t[181];
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] & t[75];
  assign t[47] = ~(t[76]);
  assign t[48] = t[174] ^ t[77];
  assign t[49] = t[78] ^ t[79];
  assign t[4] = ~(t[9]);
  assign t[50] = t[80] & t[81];
  assign t[51] = ~(t[82] & t[83]);
  assign t[52] = t[84] ^ t[182];
  assign t[53] = ~(t[175]);
  assign t[54] = t[85] & t[84];
  assign t[55] = ~(t[183]);
  assign t[56] = ~(t[86] & t[184]);
  assign t[57] = t[87] ^ t[63];
  assign t[58] = t[88] & t[89];
  assign t[59] = t[90] ^ t[43];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[91] & t[92];
  assign t[61] = t[68] ^ t[93];
  assign t[62] = t[94] ^ t[50];
  assign t[63] = t[95];
  assign t[64] = t[96] ^ t[97];
  assign t[65] = t[179] ^ t[98];
  assign t[66] = t[7] ? t[99] : t[185];
  assign t[67] = t[100] ^ t[101];
  assign t[68] = t[40] ^ t[102];
  assign t[69] = t[186] ^ t[103];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[180] ^ t[104];
  assign t[71] = t[181] ^ t[105];
  assign t[72] = t[106] & t[107];
  assign t[73] = t[108] & t[109];
  assign t[74] = ~(t[72] ^ t[110]);
  assign t[75] = t[111] ^ t[112];
  assign t[76] = ~(t[7]);
  assign t[77] = t[113] ? x[50] : x[49];
  assign t[78] = t[114] & t[115];
  assign t[79] = t[116] & t[117];
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[94] ^ t[49]);
  assign t[81] = t[118] ^ t[117];
  assign t[82] = ~(t[85] | t[84]);
  assign t[83] = ~(t[119] | t[53]);
  assign t[84] = ~(t[187]);
  assign t[85] = ~(t[182]);
  assign t[86] = ~(t[186]);
  assign t[87] = ~t[120];
  assign t[88] = ~(t[121]);
  assign t[89] = t[122];
  assign t[8] = t[172] ^ t[16];
  assign t[90] = t[47] ? t[123] : t[188];
  assign t[91] = ~(t[59] ^ t[45]);
  assign t[92] = t[23] ^ t[109];
  assign t[93] = t[67] ^ t[124];
  assign t[94] = t[125] ^ t[126];
  assign t[95] = t[7] ? t[127] : t[189];
  assign t[96] = t[128] ^ t[58];
  assign t[97] = t[129] & t[130];
  assign t[98] = t[131] ? x[61] : x[60];
  assign t[99] = t[185] ^ t[132];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind111(x, y);
 input [116:0] x;
 output y;

 wire [234:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[111]);
  assign t[101] = t[195] ^ t[130];
  assign t[102] = t[7] ? t[131] : t[203];
  assign t[103] = t[196] ^ t[132];
  assign t[104] = t[197] ^ t[133];
  assign t[105] = t[134] & t[135];
  assign t[106] = ~(t[105] ^ t[136]);
  assign t[107] = t[61] ^ t[137];
  assign t[108] = t[138] & t[139];
  assign t[109] = ~(t[119] ^ t[72]);
  assign t[10] = ~(t[19] ^ t[20]);
  assign t[110] = t[140] ^ t[42];
  assign t[111] = ~(t[7]);
  assign t[112] = t[30] ? x[76] : x[75];
  assign t[113] = t[30] ? x[78] : x[77];
  assign t[114] = t[141] & t[142];
  assign t[115] = t[198] ^ t[143];
  assign t[116] = ~(t[182]);
  assign t[117] = t[200] ^ t[144];
  assign t[118] = ~(t[47]);
  assign t[119] = t[39] ^ t[67];
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[145];
  assign t[121] = t[123] ^ t[146];
  assign t[122] = t[147];
  assign t[123] = t[148] ^ t[149];
  assign t[124] = t[150] & t[151];
  assign t[125] = t[201] ^ t[152];
  assign t[126] = t[202] ^ t[153];
  assign t[127] = t[154] ? x[80] : x[79];
  assign t[128] = ~(t[155] ^ t[70]);
  assign t[129] = t[43] ^ t[96];
  assign t[12] = t[23] ^ t[24];
  assign t[130] = t[156] ? x[82] : x[81];
  assign t[131] = t[203] ^ t[157];
  assign t[132] = t[84] ? x[84] : x[83];
  assign t[133] = t[154] ? x[86] : x[85];
  assign t[134] = ~(t[137]);
  assign t[135] = ~(t[94]);
  assign t[136] = t[43] ^ t[94];
  assign t[137] = t[96] ^ t[69];
  assign t[138] = ~(t[158]);
  assign t[139] = ~(t[39]);
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[67] ^ t[40];
  assign t[141] = ~(t[159]);
  assign t[142] = ~(t[46]);
  assign t[143] = t[30] ? x[88] : x[87];
  assign t[144] = t[30] ? x[90] : x[89];
  assign t[145] = t[7] ? t[160] : t[204];
  assign t[146] = t[161] & t[162];
  assign t[147] = t[7] ? t[163] : t[205];
  assign t[148] = t[164] & t[165];
  assign t[149] = t[166] & t[167];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = ~(t[148] ^ t[168]);
  assign t[151] = t[169] ^ t[170];
  assign t[152] = t[154] ? x[98] : x[97];
  assign t[153] = t[154] ? x[100] : x[99];
  assign t[154] = ~(t[54]);
  assign t[155] = t[94] ^ t[69];
  assign t[156] = ~(t[54]);
  assign t[157] = t[30] ? x[102] : x[101];
  assign t[158] = t[42] ^ t[67];
  assign t[159] = t[79] ^ t[47];
  assign t[15] = t[182] | t[29];
  assign t[160] = t[204] ^ t[171];
  assign t[161] = ~(t[172] ^ t[123]);
  assign t[162] = t[92] ^ t[167];
  assign t[163] = t[205] ^ t[173];
  assign t[164] = ~(t[170]);
  assign t[165] = ~(t[174]);
  assign t[166] = ~(t[122]);
  assign t[167] = t[175];
  assign t[168] = t[92] ^ t[174];
  assign t[169] = t[174] ^ t[120];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[167] ^ t[122];
  assign t[171] = t[84] ? x[104] : x[103];
  assign t[172] = t[174] ^ t[122];
  assign t[173] = t[156] ? x[106] : x[105];
  assign t[174] = ~t[176];
  assign t[175] = t[7] ? t[177] : t[206];
  assign t[176] = t[7] ? t[178] : t[207];
  assign t[177] = t[206] ^ t[179];
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[156] ? x[114] : x[113];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[84] ? x[116] : x[115];
  assign t[181] = t[208] ^ x[4];
  assign t[182] = t[209] ^ x[7];
  assign t[183] = t[210] ^ x[12];
  assign t[184] = t[211] ^ x[15];
  assign t[185] = t[212] ^ x[18];
  assign t[186] = t[213] ^ x[21];
  assign t[187] = t[214] ^ x[24];
  assign t[188] = t[215] ^ x[27];
  assign t[189] = t[216] ^ x[30];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[217] ^ x[33];
  assign t[191] = t[218] ^ x[36];
  assign t[192] = t[219] ^ x[39];
  assign t[193] = t[220] ^ x[42];
  assign t[194] = t[221] ^ x[45];
  assign t[195] = t[222] ^ x[48];
  assign t[196] = t[223] ^ x[51];
  assign t[197] = t[224] ^ x[54];
  assign t[198] = t[225] ^ x[57];
  assign t[199] = t[226] ^ x[60];
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[63];
  assign t[201] = t[228] ^ x[66];
  assign t[202] = t[229] ^ x[69];
  assign t[203] = t[230] ^ x[74];
  assign t[204] = t[231] ^ x[93];
  assign t[205] = t[232] ^ x[96];
  assign t[206] = t[233] ^ x[109];
  assign t[207] = t[234] ^ x[112];
  assign t[208] = (x[2] & x[3]);
  assign t[209] = (x[5] & x[6]);
  assign t[20] = ~(t[37] ^ t[38]);
  assign t[210] = (x[10] & x[11]);
  assign t[211] = (x[13] & x[14]);
  assign t[212] = (x[16] & x[17]);
  assign t[213] = (x[19] & x[20]);
  assign t[214] = (x[22] & x[23]);
  assign t[215] = (x[25] & x[26]);
  assign t[216] = (x[28] & x[29]);
  assign t[217] = (x[31] & x[32]);
  assign t[218] = (x[34] & x[35]);
  assign t[219] = (x[37] & x[38]);
  assign t[21] = t[39] ^ t[40];
  assign t[220] = (x[40] & x[41]);
  assign t[221] = (x[43] & x[44]);
  assign t[222] = (x[46] & x[47]);
  assign t[223] = (x[49] & x[50]);
  assign t[224] = (x[52] & x[53]);
  assign t[225] = (x[55] & x[56]);
  assign t[226] = (x[58] & x[59]);
  assign t[227] = (x[61] & x[62]);
  assign t[228] = (x[64] & x[65]);
  assign t[229] = (x[67] & x[68]);
  assign t[22] = t[41] & t[42];
  assign t[230] = (x[72] & x[73]);
  assign t[231] = (x[91] & x[92]);
  assign t[232] = (x[94] & x[95]);
  assign t[233] = (x[107] & x[108]);
  assign t[234] = (x[110] & x[111]);
  assign t[23] = t[43] ^ t[44];
  assign t[24] = t[40] ^ t[45];
  assign t[25] = t[46] ^ t[47];
  assign t[26] = t[48] & t[49];
  assign t[27] = ~(t[29] & t[50]);
  assign t[28] = ~(t[183] ^ t[51]);
  assign t[29] = ~(t[52] & t[53]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[54]);
  assign t[31] = ~(t[184]);
  assign t[32] = ~(t[185]);
  assign t[33] = ~(t[186]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = t[57] ^ t[58];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[37] = t[61] ^ t[62];
  assign t[38] = t[63] ^ t[64];
  assign t[39] = t[7] ? t[65] : t[187];
  assign t[3] = t[7] ? t[8] : t[181];
  assign t[40] = t[188] ^ t[66];
  assign t[41] = ~(t[67]);
  assign t[42] = t[189] ^ t[68];
  assign t[43] = t[69] ^ t[63];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] ? t[75] : t[190];
  assign t[47] = t[74] ? t[76] : t[191];
  assign t[48] = ~(t[25] ^ t[77]);
  assign t[49] = t[78] ^ t[79];
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[80] & t[81]);
  assign t[51] = t[82] ^ t[192];
  assign t[52] = ~(t[183]);
  assign t[53] = t[83] & t[82];
  assign t[54] = ~(t[84]);
  assign t[55] = ~(t[188]);
  assign t[56] = ~(t[85] & t[193]);
  assign t[57] = t[86] ^ t[87];
  assign t[58] = t[88] ^ t[89];
  assign t[59] = ~(t[90] ^ t[91]);
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[94] ^ t[63];
  assign t[62] = t[95] & t[96];
  assign t[63] = t[74] ? t[97] : t[194];
  assign t[64] = t[70] ^ t[98];
  assign t[65] = t[187] ^ t[99];
  assign t[66] = t[100] ? t[101] : t[195];
  assign t[67] = t[186] ^ t[102];
  assign t[68] = t[7] ? t[103] : t[196];
  assign t[69] = t[74] ? t[104] : t[197];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[105] ^ t[62];
  assign t[71] = t[106] & t[107];
  assign t[72] = t[108] ^ t[22];
  assign t[73] = t[109] & t[110];
  assign t[74] = ~(t[111]);
  assign t[75] = t[190] ^ t[112];
  assign t[76] = t[191] ^ t[113];
  assign t[77] = t[114] ^ t[89];
  assign t[78] = t[47] ^ t[86];
  assign t[79] = t[74] ? t[115] : t[198];
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[83] | t[82]);
  assign t[81] = ~(t[116] | t[52]);
  assign t[82] = ~(t[199]);
  assign t[83] = ~(t[192]);
  assign t[84] = ~(t[15]);
  assign t[85] = ~(t[189]);
  assign t[86] = t[74] ? t[117] : t[200];
  assign t[87] = t[77] ^ t[26];
  assign t[88] = t[46] ^ t[86];
  assign t[89] = t[118] & t[79];
  assign t[8] = t[181] ^ t[16];
  assign t[90] = t[119] ^ t[73];
  assign t[91] = t[120] ^ t[121];
  assign t[92] = t[122] ^ t[120];
  assign t[93] = t[123] ^ t[124];
  assign t[94] = t[74] ? t[125] : t[201];
  assign t[95] = ~(t[69]);
  assign t[96] = t[74] ? t[126] : t[202];
  assign t[97] = t[194] ^ t[127];
  assign t[98] = t[128] & t[129];
  assign t[99] = t[30] ? x[71] : x[70];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind112(x, y);
 input [116:0] x;
 output y;

 wire [245:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[35] ? t[125] : t[208];
  assign t[101] = t[35] ? t[126] : t[209];
  assign t[102] = ~(t[70] ^ t[127]);
  assign t[103] = t[128] ^ t[129];
  assign t[104] = t[128] ^ t[130];
  assign t[105] = t[131] ^ t[132];
  assign t[106] = t[133] & t[134];
  assign t[107] = t[135] & t[136];
  assign t[108] = t[132] ^ t[137];
  assign t[109] = t[138] ^ t[139];
  assign t[10] = t[19] ^ t[20];
  assign t[110] = t[140] ^ t[42];
  assign t[111] = t[35] ? t[141] : t[210];
  assign t[112] = t[127] ^ t[71];
  assign t[113] = ~(t[193]);
  assign t[114] = t[41] ^ t[63];
  assign t[115] = t[85] ? x[68] : x[67];
  assign t[116] = t[142] ? x[70] : x[69];
  assign t[117] = ~(t[143]);
  assign t[118] = ~(t[140]);
  assign t[119] = ~(t[98]);
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[207] ^ t[144];
  assign t[121] = t[140] ^ t[98];
  assign t[122] = t[7] ? t[145] : t[211];
  assign t[123] = ~(t[94] ^ t[146]);
  assign t[124] = t[110] ^ t[143];
  assign t[125] = t[208] ^ t[147];
  assign t[126] = t[209] ^ t[148];
  assign t[127] = t[149] ^ t[150];
  assign t[128] = t[101] ^ t[111];
  assign t[129] = t[35] ? t[151] : t[212];
  assign t[12] = ~(t[23] ^ t[24]);
  assign t[130] = t[127] ^ t[152];
  assign t[131] = ~t[153];
  assign t[132] = t[154];
  assign t[133] = ~(t[105] ^ t[138]);
  assign t[134] = t[108] ^ t[155];
  assign t[135] = ~(t[59] ^ t[156]);
  assign t[136] = t[21] ^ t[114];
  assign t[137] = t[157];
  assign t[138] = t[158] ^ t[159];
  assign t[139] = t[160] & t[161];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[7] ? t[162] : t[213];
  assign t[141] = t[210] ^ t[163];
  assign t[142] = ~(t[54]);
  assign t[143] = t[120] ^ t[98];
  assign t[144] = t[7] ? t[164] : t[214];
  assign t[145] = t[211] ^ t[165];
  assign t[146] = t[68] ^ t[140];
  assign t[147] = t[30] ? x[84] : x[83];
  assign t[148] = t[30] ? x[86] : x[85];
  assign t[149] = t[166] & t[167];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[168] & t[129];
  assign t[151] = t[212] ^ t[169];
  assign t[152] = t[170] & t[171];
  assign t[153] = t[7] ? t[172] : t[215];
  assign t[154] = t[7] ? t[173] : t[216];
  assign t[155] = t[174];
  assign t[156] = t[74] ^ t[39];
  assign t[157] = t[7] ? t[175] : t[217];
  assign t[158] = t[176] & t[177];
  assign t[159] = t[178] & t[155];
  assign t[15] = t[193] | t[29];
  assign t[160] = ~(t[158] ^ t[179]);
  assign t[161] = t[180] ^ t[181];
  assign t[162] = t[213] ^ t[182];
  assign t[163] = t[30] ? x[97] : x[96];
  assign t[164] = t[214] ^ t[183];
  assign t[165] = t[85] ? x[99] : x[98];
  assign t[166] = ~(t[184]);
  assign t[167] = ~(t[100]);
  assign t[168] = ~(t[101]);
  assign t[169] = t[30] ? x[101] : x[100];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = ~(t[149] ^ t[185]);
  assign t[171] = t[186] ^ t[184];
  assign t[172] = t[215] ^ t[187];
  assign t[173] = t[216] ^ t[188];
  assign t[174] = t[7] ? t[189] : t[218];
  assign t[175] = t[217] ^ t[190];
  assign t[176] = ~(t[181]);
  assign t[177] = ~(t[131]);
  assign t[178] = ~(t[132]);
  assign t[179] = t[108] ^ t[131];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[131] ^ t[137];
  assign t[181] = t[155] ^ t[132];
  assign t[182] = t[85] ? x[106] : x[105];
  assign t[183] = t[83] ? x[108] : x[107];
  assign t[184] = t[129] ^ t[101];
  assign t[185] = t[128] ^ t[100];
  assign t[186] = t[100] ^ t[111];
  assign t[187] = t[83] ? x[110] : x[109];
  assign t[188] = t[142] ? x[112] : x[111];
  assign t[189] = t[218] ^ t[191];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[83] ? x[114] : x[113];
  assign t[191] = t[142] ? x[116] : x[115];
  assign t[192] = t[219] ^ x[4];
  assign t[193] = t[220] ^ x[7];
  assign t[194] = t[221] ^ x[12];
  assign t[195] = t[222] ^ x[15];
  assign t[196] = t[223] ^ x[18];
  assign t[197] = t[224] ^ x[21];
  assign t[198] = t[225] ^ x[24];
  assign t[199] = t[226] ^ x[27];
  assign t[19] = t[35] ? t[36] : t[194];
  assign t[1] = ~(t[4]);
  assign t[200] = t[227] ^ x[30];
  assign t[201] = t[228] ^ x[33];
  assign t[202] = t[229] ^ x[36];
  assign t[203] = t[230] ^ x[39];
  assign t[204] = t[231] ^ x[44];
  assign t[205] = t[232] ^ x[47];
  assign t[206] = t[233] ^ x[50];
  assign t[207] = t[234] ^ x[53];
  assign t[208] = t[235] ^ x[60];
  assign t[209] = t[236] ^ x[63];
  assign t[20] = t[37] ^ t[38];
  assign t[210] = t[237] ^ x[66];
  assign t[211] = t[238] ^ x[73];
  assign t[212] = t[239] ^ x[76];
  assign t[213] = t[240] ^ x[79];
  assign t[214] = t[241] ^ x[82];
  assign t[215] = t[242] ^ x[89];
  assign t[216] = t[243] ^ x[92];
  assign t[217] = t[244] ^ x[95];
  assign t[218] = t[245] ^ x[104];
  assign t[219] = (x[2] & x[3]);
  assign t[21] = t[39] ^ t[19];
  assign t[220] = (x[5] & x[6]);
  assign t[221] = (x[10] & x[11]);
  assign t[222] = (x[13] & x[14]);
  assign t[223] = (x[16] & x[17]);
  assign t[224] = (x[19] & x[20]);
  assign t[225] = (x[22] & x[23]);
  assign t[226] = (x[25] & x[26]);
  assign t[227] = (x[28] & x[29]);
  assign t[228] = (x[31] & x[32]);
  assign t[229] = (x[34] & x[35]);
  assign t[22] = t[40] & t[41];
  assign t[230] = (x[37] & x[38]);
  assign t[231] = (x[42] & x[43]);
  assign t[232] = (x[45] & x[46]);
  assign t[233] = (x[48] & x[49]);
  assign t[234] = (x[51] & x[52]);
  assign t[235] = (x[58] & x[59]);
  assign t[236] = (x[61] & x[62]);
  assign t[237] = (x[64] & x[65]);
  assign t[238] = (x[71] & x[72]);
  assign t[239] = (x[74] & x[75]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (x[77] & x[78]);
  assign t[241] = (x[80] & x[81]);
  assign t[242] = (x[87] & x[88]);
  assign t[243] = (x[90] & x[91]);
  assign t[244] = (x[93] & x[94]);
  assign t[245] = (x[102] & x[103]);
  assign t[24] = t[44] ^ t[45];
  assign t[25] = ~(t[46] ^ t[47]);
  assign t[26] = ~(t[48] ^ t[49]);
  assign t[27] = ~(t[29] & t[50]);
  assign t[28] = ~(t[195] ^ t[51]);
  assign t[29] = ~(t[52] & t[53]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = ~(t[54]);
  assign t[31] = ~(t[196]);
  assign t[32] = ~(t[197]);
  assign t[33] = ~(t[198]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = ~(t[57]);
  assign t[36] = t[194] ^ t[58];
  assign t[37] = t[59] ^ t[22];
  assign t[38] = t[60] & t[61];
  assign t[39] = t[35] ? t[62] : t[199];
  assign t[3] = t[7] ? t[8] : t[192];
  assign t[40] = ~(t[63]);
  assign t[41] = t[35] ? t[64] : t[200];
  assign t[42] = t[201] ^ t[65];
  assign t[43] = t[66] ^ t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] ^ t[73]);
  assign t[47] = t[74] ^ t[75];
  assign t[48] = t[76] ^ t[77];
  assign t[49] = ~(t[10] ^ t[78]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[79] & t[80]);
  assign t[51] = t[81] ^ t[202];
  assign t[52] = ~(t[195]);
  assign t[53] = t[82] & t[81];
  assign t[54] = ~(t[83]);
  assign t[55] = ~(t[201]);
  assign t[56] = ~(t[84] & t[203]);
  assign t[57] = ~(t[7]);
  assign t[58] = t[85] ? x[41] : x[40];
  assign t[59] = t[86] & t[87];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = ~(t[88] ^ t[37]);
  assign t[61] = t[74] ^ t[41];
  assign t[62] = t[199] ^ t[89];
  assign t[63] = t[35] ? t[90] : t[204];
  assign t[64] = t[200] ^ t[91];
  assign t[65] = t[92] ? t[93] : t[205];
  assign t[66] = t[94] ^ t[95];
  assign t[67] = t[96] & t[97];
  assign t[68] = t[98] ^ t[42];
  assign t[69] = t[66] ^ t[99];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[100] ^ t[101];
  assign t[71] = t[102] & t[103];
  assign t[72] = t[104] ^ t[23];
  assign t[73] = t[105] ^ t[106];
  assign t[74] = t[63] ^ t[19];
  assign t[75] = t[37] ^ t[107];
  assign t[76] = t[108] ^ t[109];
  assign t[77] = t[110] ^ t[95];
  assign t[78] = t[111] ^ t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[113] | t[52]);
  assign t[81] = ~(t[206]);
  assign t[82] = ~(t[202]);
  assign t[83] = ~(t[15]);
  assign t[84] = ~(t[207]);
  assign t[85] = ~(t[54]);
  assign t[86] = ~(t[114]);
  assign t[87] = ~(t[39]);
  assign t[88] = t[39] ^ t[63];
  assign t[89] = t[85] ? x[55] : x[54];
  assign t[8] = t[192] ^ t[16];
  assign t[90] = t[204] ^ t[115];
  assign t[91] = t[85] ? x[57] : x[56];
  assign t[92] = ~(t[57]);
  assign t[93] = t[205] ^ t[116];
  assign t[94] = t[117] & t[118];
  assign t[95] = t[119] & t[120];
  assign t[96] = ~(t[121] ^ t[66]);
  assign t[97] = t[68] ^ t[120];
  assign t[98] = t[198] ^ t[122];
  assign t[99] = t[123] & t[124];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind113(x, y);
 input [116:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[41] ^ t[123];
  assign t[101] = ~t[124];
  assign t[102] = t[125];
  assign t[103] = ~(t[69] ^ t[126]);
  assign t[104] = t[127] ^ t[128];
  assign t[105] = t[187] ^ t[129];
  assign t[106] = ~(t[75] ^ t[130]);
  assign t[107] = t[131] ^ t[132];
  assign t[108] = ~(t[133]);
  assign t[109] = ~(t[132]);
  assign t[10] = t[19] ^ t[20];
  assign t[110] = ~(t[134]);
  assign t[111] = ~(t[71]);
  assign t[112] = t[47] ? t[135] : t[190];
  assign t[113] = t[134] ^ t[71];
  assign t[114] = ~(t[172]);
  assign t[115] = ~(t[133]);
  assign t[116] = t[115] ? x[73] : x[72];
  assign t[117] = t[108] ? x[75] : x[74];
  assign t[118] = t[136] ? x[77] : x[76];
  assign t[119] = t[7] ? t[137] : t[191];
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[7] ? t[138] : t[192];
  assign t[121] = t[139] ^ t[20];
  assign t[122] = t[140] & t[141];
  assign t[123] = t[142] & t[143];
  assign t[124] = t[7] ? t[144] : t[193];
  assign t[125] = t[7] ? t[145] : t[194];
  assign t[126] = t[146] ^ t[147];
  assign t[127] = t[102] ^ t[148];
  assign t[128] = t[149];
  assign t[129] = t[108] ? x[91] : x[90];
  assign t[12] = ~(t[23] ^ t[24]);
  assign t[130] = t[45] ^ t[134];
  assign t[131] = t[134] ^ t[25];
  assign t[132] = t[112] ^ t[71];
  assign t[133] = ~(t[30]);
  assign t[134] = t[47] ? t[150] : t[195];
  assign t[135] = t[190] ^ t[151];
  assign t[136] = ~(t[133]);
  assign t[137] = t[191] ^ t[152];
  assign t[138] = t[192] ^ t[153];
  assign t[139] = t[154] & t[155];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = ~(t[139] ^ t[156]);
  assign t[141] = t[19] ^ t[157];
  assign t[142] = ~(t[158] ^ t[41]);
  assign t[143] = t[21] ^ t[94];
  assign t[144] = t[193] ^ t[159];
  assign t[145] = t[194] ^ t[160];
  assign t[146] = t[161] & t[162];
  assign t[147] = t[163] & t[128];
  assign t[148] = t[164];
  assign t[149] = t[7] ? t[165] : t[196];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[195] ^ t[166];
  assign t[151] = t[108] ? x[99] : x[98];
  assign t[152] = t[108] ? x[101] : x[100];
  assign t[153] = t[30] ? x[103] : x[102];
  assign t[154] = ~(t[157]);
  assign t[155] = ~(t[35]);
  assign t[156] = t[98] ^ t[35];
  assign t[157] = t[38] ^ t[59];
  assign t[158] = t[119] ^ t[39];
  assign t[159] = t[30] ? x[105] : x[104];
  assign t[15] = t[172] | t[29];
  assign t[160] = t[136] ? x[107] : x[106];
  assign t[161] = ~(t[167]);
  assign t[162] = ~(t[101]);
  assign t[163] = ~(t[102]);
  assign t[164] = t[7] ? t[168] : t[197];
  assign t[165] = t[196] ^ t[169];
  assign t[166] = t[108] ? x[112] : x[111];
  assign t[167] = t[128] ^ t[102];
  assign t[168] = t[197] ^ t[170];
  assign t[169] = t[136] ? x[114] : x[113];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[30] ? x[116] : x[115];
  assign t[171] = t[198] ^ x[4];
  assign t[172] = t[199] ^ x[7];
  assign t[173] = t[200] ^ x[12];
  assign t[174] = t[201] ^ x[15];
  assign t[175] = t[202] ^ x[18];
  assign t[176] = t[203] ^ x[21];
  assign t[177] = t[204] ^ x[24];
  assign t[178] = t[205] ^ x[27];
  assign t[179] = t[206] ^ x[30];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[207] ^ x[33];
  assign t[181] = t[208] ^ x[36];
  assign t[182] = t[209] ^ x[39];
  assign t[183] = t[210] ^ x[42];
  assign t[184] = t[211] ^ x[45];
  assign t[185] = t[212] ^ x[48];
  assign t[186] = t[213] ^ x[51];
  assign t[187] = t[214] ^ x[54];
  assign t[188] = t[215] ^ x[59];
  assign t[189] = t[216] ^ x[62];
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = t[217] ^ x[71];
  assign t[191] = t[218] ^ x[80];
  assign t[192] = t[219] ^ x[83];
  assign t[193] = t[220] ^ x[86];
  assign t[194] = t[221] ^ x[89];
  assign t[195] = t[222] ^ x[94];
  assign t[196] = t[223] ^ x[97];
  assign t[197] = t[224] ^ x[110];
  assign t[198] = (x[2] & x[3]);
  assign t[199] = (x[5] & x[6]);
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[10] & x[11]);
  assign t[201] = (x[13] & x[14]);
  assign t[202] = (x[16] & x[17]);
  assign t[203] = (x[19] & x[20]);
  assign t[204] = (x[22] & x[23]);
  assign t[205] = (x[25] & x[26]);
  assign t[206] = (x[28] & x[29]);
  assign t[207] = (x[31] & x[32]);
  assign t[208] = (x[34] & x[35]);
  assign t[209] = (x[37] & x[38]);
  assign t[20] = t[37] & t[38];
  assign t[210] = (x[40] & x[41]);
  assign t[211] = (x[43] & x[44]);
  assign t[212] = (x[46] & x[47]);
  assign t[213] = (x[49] & x[50]);
  assign t[214] = (x[52] & x[53]);
  assign t[215] = (x[57] & x[58]);
  assign t[216] = (x[60] & x[61]);
  assign t[217] = (x[69] & x[70]);
  assign t[218] = (x[78] & x[79]);
  assign t[219] = (x[81] & x[82]);
  assign t[21] = t[39] ^ t[40];
  assign t[220] = (x[84] & x[85]);
  assign t[221] = (x[87] & x[88]);
  assign t[222] = (x[92] & x[93]);
  assign t[223] = (x[95] & x[96]);
  assign t[224] = (x[108] & x[109]);
  assign t[22] = t[41] ^ t[42];
  assign t[23] = ~(t[43] ^ t[44]);
  assign t[24] = t[45] ^ t[46];
  assign t[25] = t[47] ? t[48] : t[173];
  assign t[26] = t[49] ^ t[50];
  assign t[27] = ~(t[29] & t[51]);
  assign t[28] = ~(t[174] ^ t[52]);
  assign t[29] = ~(t[53] & t[54]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[15]);
  assign t[31] = ~(t[175]);
  assign t[32] = ~(t[176]);
  assign t[33] = ~(t[177]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = t[47] ? t[57] : t[178];
  assign t[36] = t[47] ? t[58] : t[179];
  assign t[37] = ~(t[59]);
  assign t[38] = t[47] ? t[60] : t[180];
  assign t[39] = t[177] ^ t[61];
  assign t[3] = t[7] ? t[8] : t[171];
  assign t[40] = t[181] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[67] ^ t[68];
  assign t[44] = t[69] ^ t[70];
  assign t[45] = t[71] ^ t[25];
  assign t[46] = t[49] ^ t[72];
  assign t[47] = ~(t[73]);
  assign t[48] = t[173] ^ t[74];
  assign t[49] = t[75] ^ t[76];
  assign t[4] = ~(t[9]);
  assign t[50] = t[77] & t[78];
  assign t[51] = ~(t[79] & t[80]);
  assign t[52] = t[81] ^ t[182];
  assign t[53] = ~(t[174]);
  assign t[54] = t[82] & t[81];
  assign t[55] = ~(t[181]);
  assign t[56] = ~(t[83] & t[183]);
  assign t[57] = t[178] ^ t[84];
  assign t[58] = t[179] ^ t[85];
  assign t[59] = t[47] ? t[86] : t[184];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[180] ^ t[87];
  assign t[61] = t[7] ? t[88] : t[185];
  assign t[62] = t[89] ? t[90] : t[186];
  assign t[63] = t[91] & t[92];
  assign t[64] = t[93] & t[94];
  assign t[65] = ~(t[63] ^ t[95]);
  assign t[66] = t[96] ^ t[97];
  assign t[67] = t[98] ^ t[99];
  assign t[68] = t[40] ^ t[100];
  assign t[69] = t[101] ^ t[102];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[103] & t[104];
  assign t[71] = t[47] ? t[105] : t[187];
  assign t[72] = t[106] & t[107];
  assign t[73] = ~(t[7]);
  assign t[74] = t[108] ? x[56] : x[55];
  assign t[75] = t[109] & t[110];
  assign t[76] = t[111] & t[112];
  assign t[77] = ~(t[113] ^ t[49]);
  assign t[78] = t[45] ^ t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[114] | t[53]);
  assign t[81] = ~(t[188]);
  assign t[82] = ~(t[182]);
  assign t[83] = ~(t[189]);
  assign t[84] = t[115] ? x[64] : x[63];
  assign t[85] = t[115] ? x[66] : x[65];
  assign t[86] = t[184] ^ t[116];
  assign t[87] = t[115] ? x[68] : x[67];
  assign t[88] = t[185] ^ t[117];
  assign t[89] = ~(t[73]);
  assign t[8] = t[171] ^ t[16];
  assign t[90] = t[186] ^ t[118];
  assign t[91] = ~(t[97]);
  assign t[92] = ~(t[119]);
  assign t[93] = ~(t[39]);
  assign t[94] = t[189] ^ t[120];
  assign t[95] = t[21] ^ t[119];
  assign t[96] = t[119] ^ t[40];
  assign t[97] = t[94] ^ t[39];
  assign t[98] = t[59] ^ t[36];
  assign t[99] = t[121] ^ t[122];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind114(x, y);
 input [111:0] x;
 output y;

 wire [202:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[167] ^ t[127];
  assign t[101] = ~(t[107]);
  assign t[102] = ~(t[128]);
  assign t[103] = ~(t[51]);
  assign t[104] = t[155] ^ t[129];
  assign t[105] = t[32] ^ t[128];
  assign t[106] = t[128] ^ t[52];
  assign t[107] = t[104] ^ t[51];
  assign t[108] = t[74] ? x[71] : x[70];
  assign t[109] = ~(t[130]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = ~(t[131]);
  assign t[111] = ~(t[132]);
  assign t[112] = t[133];
  assign t[113] = t[131] ^ t[132];
  assign t[114] = t[132] ^ t[34];
  assign t[115] = ~(t[134]);
  assign t[116] = ~(t[3]);
  assign t[117] = ~(t[36]);
  assign t[118] = t[168] ^ t[135];
  assign t[119] = t[27] ? x[73] : x[72];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[169] ^ t[136];
  assign t[121] = t[92] ? x[75] : x[74];
  assign t[122] = ~(t[125] | t[124]);
  assign t[123] = ~(t[137] | t[97]);
  assign t[124] = ~(t[171]);
  assign t[125] = ~(t[170]);
  assign t[126] = t[138] ? x[80] : x[79];
  assign t[127] = t[74] ? x[82] : x[81];
  assign t[128] = t[39] ? t[139] : t[172];
  assign t[129] = t[39] ? t[140] : t[173];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[112] ^ t[132];
  assign t[131] = ~t[141];
  assign t[132] = t[142];
  assign t[133] = t[26] ? t[143] : t[174];
  assign t[134] = t[61] ^ t[36];
  assign t[135] = t[27] ? x[93] : x[92];
  assign t[136] = t[92] ? x[95] : x[94];
  assign t[137] = ~(t[158]);
  assign t[138] = ~(t[48]);
  assign t[139] = t[172] ^ t[144];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[173] ^ t[145];
  assign t[141] = t[26] ? t[146] : t[175];
  assign t[142] = t[26] ? t[147] : t[176];
  assign t[143] = t[174] ^ t[148];
  assign t[144] = t[74] ? x[103] : x[102];
  assign t[145] = t[138] ? x[105] : x[104];
  assign t[146] = t[175] ^ t[149];
  assign t[147] = t[176] ^ t[150];
  assign t[148] = t[92] ? x[107] : x[106];
  assign t[149] = t[74] ? x[109] : x[108];
  assign t[14] = ~(t[26]);
  assign t[150] = t[138] ? x[111] : x[110];
  assign t[151] = t[177] ^ x[4];
  assign t[152] = t[178] ^ x[9];
  assign t[153] = t[179] ^ x[12];
  assign t[154] = t[180] ^ x[15];
  assign t[155] = t[181] ^ x[18];
  assign t[156] = t[182] ^ x[21];
  assign t[157] = t[183] ^ x[24];
  assign t[158] = t[184] ^ x[27];
  assign t[159] = t[185] ^ x[30];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[186] ^ x[33];
  assign t[161] = t[187] ^ x[36];
  assign t[162] = t[188] ^ x[39];
  assign t[163] = t[189] ^ x[46];
  assign t[164] = t[190] ^ x[49];
  assign t[165] = t[191] ^ x[52];
  assign t[166] = t[192] ^ x[55];
  assign t[167] = t[193] ^ x[58];
  assign t[168] = t[194] ^ x[63];
  assign t[169] = t[195] ^ x[66];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[196] ^ x[69];
  assign t[171] = t[197] ^ x[78];
  assign t[172] = t[198] ^ x[85];
  assign t[173] = t[199] ^ x[88];
  assign t[174] = t[200] ^ x[91];
  assign t[175] = t[201] ^ x[98];
  assign t[176] = t[202] ^ x[101];
  assign t[177] = (x[2] & x[3]);
  assign t[178] = (x[7] & x[8]);
  assign t[179] = (x[10] & x[11]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = (x[13] & x[14]);
  assign t[181] = (x[16] & x[17]);
  assign t[182] = (x[19] & x[20]);
  assign t[183] = (x[22] & x[23]);
  assign t[184] = (x[25] & x[26]);
  assign t[185] = (x[28] & x[29]);
  assign t[186] = (x[31] & x[32]);
  assign t[187] = (x[34] & x[35]);
  assign t[188] = (x[37] & x[38]);
  assign t[189] = (x[44] & x[45]);
  assign t[18] = t[32] ^ t[33];
  assign t[190] = (x[47] & x[48]);
  assign t[191] = (x[50] & x[51]);
  assign t[192] = (x[53] & x[54]);
  assign t[193] = (x[56] & x[57]);
  assign t[194] = (x[61] & x[62]);
  assign t[195] = (x[64] & x[65]);
  assign t[196] = (x[67] & x[68]);
  assign t[197] = (x[76] & x[77]);
  assign t[198] = (x[83] & x[84]);
  assign t[199] = (x[86] & x[87]);
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[89] & x[90]);
  assign t[201] = (x[96] & x[97]);
  assign t[202] = (x[99] & x[100]);
  assign t[20] = t[3] ^ t[36];
  assign t[21] = t[37] & t[38];
  assign t[22] = t[39] ? t[40] : t[152];
  assign t[23] = t[39] ? t[41] : t[153];
  assign t[24] = t[42] ^ t[43];
  assign t[25] = t[44] & t[45];
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[154]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[156]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[51] ^ t[52];
  assign t[33] = t[53] ^ t[54];
  assign t[34] = ~t[55];
  assign t[35] = t[56] ^ t[57];
  assign t[36] = t[7] ? t[58] : t[157];
  assign t[37] = ~(t[20] ^ t[59]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = ~(t[14]);
  assign t[3] = t[7] ? t[8] : t[151];
  assign t[40] = t[152] ^ t[62];
  assign t[41] = t[153] ^ t[63];
  assign t[42] = t[64] & t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = ~(t[42] ^ t[68]);
  assign t[45] = t[69] ^ t[70];
  assign t[46] = ~(t[71] & t[72]);
  assign t[47] = t[158] | t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = ~(t[159]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[75] & t[160]);
  assign t[51] = t[154] ^ t[76];
  assign t[52] = t[160] ^ t[77];
  assign t[53] = t[78] ^ t[79];
  assign t[54] = t[80] & t[81];
  assign t[55] = t[26] ? t[82] : t[161];
  assign t[56] = t[83] ^ t[84];
  assign t[57] = t[85] & t[86];
  assign t[58] = t[157] ^ t[87];
  assign t[59] = t[88] ^ t[89];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[36] ^ t[90];
  assign t[61] = t[7] ? t[91] : t[162];
  assign t[62] = t[92] ? x[41] : x[40];
  assign t[63] = t[92] ? x[43] : x[42];
  assign t[64] = ~(t[70]);
  assign t[65] = ~(t[93]);
  assign t[66] = ~(t[22]);
  assign t[67] = t[39] ? t[94] : t[163];
  assign t[68] = t[12] ^ t[93];
  assign t[69] = t[93] ^ t[23];
  assign t[6] = t[12] ^ t[13];
  assign t[70] = t[67] ^ t[22];
  assign t[71] = ~(t[73] & t[95]);
  assign t[72] = ~(t[164] ^ t[96]);
  assign t[73] = ~(t[97] & t[98]);
  assign t[74] = ~(t[47]);
  assign t[75] = ~(t[165]);
  assign t[76] = t[26] ? t[99] : t[166];
  assign t[77] = t[39] ? t[100] : t[167];
  assign t[78] = t[101] & t[102];
  assign t[79] = t[103] & t[104];
  assign t[7] = ~(t[14]);
  assign t[80] = ~(t[78] ^ t[105]);
  assign t[81] = t[106] ^ t[107];
  assign t[82] = t[161] ^ t[108];
  assign t[83] = t[109] & t[110];
  assign t[84] = t[111] & t[112];
  assign t[85] = ~(t[113] ^ t[56]);
  assign t[86] = t[114] ^ t[112];
  assign t[87] = t[27] ? x[60] : x[59];
  assign t[88] = t[115] & t[116];
  assign t[89] = t[117] & t[61];
  assign t[8] = t[151] ^ t[15];
  assign t[90] = t[7] ? t[118] : t[168];
  assign t[91] = t[162] ^ t[119];
  assign t[92] = ~(t[48]);
  assign t[93] = t[39] ? t[120] : t[169];
  assign t[94] = t[163] ^ t[121];
  assign t[95] = ~(t[122] & t[123]);
  assign t[96] = t[124] ^ t[170];
  assign t[97] = ~(t[164]);
  assign t[98] = t[125] & t[124];
  assign t[99] = t[166] ^ t[126];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind115(x, y);
 input [111:0] x;
 output y;

 wire [203:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[166]);
  assign t[101] = t[128] & t[127];
  assign t[102] = t[27] ? x[76] : x[75];
  assign t[103] = ~(t[47]);
  assign t[104] = ~(t[129]);
  assign t[105] = ~(t[34]);
  assign t[106] = ~(t[35]);
  assign t[107] = t[168] ^ t[130];
  assign t[108] = t[103] ? x[78] : x[77];
  assign t[109] = t[169] ^ t[131];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[170] ^ t[132];
  assign t[111] = ~(t[117]);
  assign t[112] = ~(t[133]);
  assign t[113] = ~(t[58]);
  assign t[114] = t[134];
  assign t[115] = t[38] ^ t[133];
  assign t[116] = t[133] ^ t[59];
  assign t[117] = t[114] ^ t[58];
  assign t[118] = t[73] ? x[80] : x[79];
  assign t[119] = t[171] ^ t[135];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[136] & t[137];
  assign t[121] = t[138] & t[93];
  assign t[122] = t[162] ^ t[139];
  assign t[123] = t[52] ? t[140] : t[173];
  assign t[124] = t[3] ^ t[51];
  assign t[125] = ~(t[128] | t[127]);
  assign t[126] = ~(t[141] | t[100]);
  assign t[127] = ~(t[174]);
  assign t[128] = ~(t[172]);
  assign t[129] = t[57] ^ t[35];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[103] ? x[88] : x[87];
  assign t[131] = t[142] ? x[90] : x[89];
  assign t[132] = t[73] ? x[92] : x[91];
  assign t[133] = ~t[143];
  assign t[134] = t[26] ? t[144] : t[175];
  assign t[135] = t[142] ? x[97] : x[96];
  assign t[136] = ~(t[145]);
  assign t[137] = ~(t[62]);
  assign t[138] = ~(t[63]);
  assign t[139] = t[52] ? t[146] : t[176];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[173] ^ t[147];
  assign t[141] = ~(t[160]);
  assign t[142] = ~(t[47]);
  assign t[143] = t[26] ? t[148] : t[177];
  assign t[144] = t[175] ^ t[149];
  assign t[145] = t[93] ^ t[63];
  assign t[146] = t[176] ^ t[150];
  assign t[147] = t[142] ? x[105] : x[104];
  assign t[148] = t[177] ^ t[151];
  assign t[149] = t[103] ? x[107] : x[106];
  assign t[14] = ~(t[26]);
  assign t[150] = t[73] ? x[109] : x[108];
  assign t[151] = t[73] ? x[111] : x[110];
  assign t[152] = t[178] ^ x[4];
  assign t[153] = t[179] ^ x[9];
  assign t[154] = t[180] ^ x[12];
  assign t[155] = t[181] ^ x[15];
  assign t[156] = t[182] ^ x[18];
  assign t[157] = t[183] ^ x[21];
  assign t[158] = t[184] ^ x[24];
  assign t[159] = t[185] ^ x[27];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[186] ^ x[30];
  assign t[161] = t[187] ^ x[33];
  assign t[162] = t[188] ^ x[36];
  assign t[163] = t[189] ^ x[39];
  assign t[164] = t[190] ^ x[42];
  assign t[165] = t[191] ^ x[45];
  assign t[166] = t[192] ^ x[50];
  assign t[167] = t[193] ^ x[53];
  assign t[168] = t[194] ^ x[62];
  assign t[169] = t[195] ^ x[65];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[196] ^ x[68];
  assign t[171] = t[197] ^ x[71];
  assign t[172] = t[198] ^ x[74];
  assign t[173] = t[199] ^ x[83];
  assign t[174] = t[200] ^ x[86];
  assign t[175] = t[201] ^ x[95];
  assign t[176] = t[202] ^ x[100];
  assign t[177] = t[203] ^ x[103];
  assign t[178] = (x[2] & x[3]);
  assign t[179] = (x[7] & x[8]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = (x[10] & x[11]);
  assign t[181] = (x[13] & x[14]);
  assign t[182] = (x[16] & x[17]);
  assign t[183] = (x[19] & x[20]);
  assign t[184] = (x[22] & x[23]);
  assign t[185] = (x[25] & x[26]);
  assign t[186] = (x[28] & x[29]);
  assign t[187] = (x[31] & x[32]);
  assign t[188] = (x[34] & x[35]);
  assign t[189] = (x[37] & x[38]);
  assign t[18] = t[32] ^ t[24];
  assign t[190] = (x[40] & x[41]);
  assign t[191] = (x[43] & x[44]);
  assign t[192] = (x[48] & x[49]);
  assign t[193] = (x[51] & x[52]);
  assign t[194] = (x[60] & x[61]);
  assign t[195] = (x[63] & x[64]);
  assign t[196] = (x[66] & x[67]);
  assign t[197] = (x[69] & x[70]);
  assign t[198] = (x[72] & x[73]);
  assign t[199] = (x[81] & x[82]);
  assign t[19] = t[33] & t[3];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[84] & x[85]);
  assign t[201] = (x[93] & x[94]);
  assign t[202] = (x[98] & x[99]);
  assign t[203] = (x[101] & x[102]);
  assign t[20] = t[34] ^ t[35];
  assign t[21] = t[36] & t[37];
  assign t[22] = t[38] ^ t[39];
  assign t[23] = t[40] ^ t[41];
  assign t[24] = t[7] ? t[42] : t[153];
  assign t[25] = t[43] ^ t[44];
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[154]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[156]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = t[7] ? t[50] : t[157];
  assign t[33] = ~(t[51]);
  assign t[34] = t[52] ? t[53] : t[158];
  assign t[35] = t[52] ? t[54] : t[159];
  assign t[36] = ~(t[20] ^ t[55]);
  assign t[37] = t[56] ^ t[57];
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[60] ^ t[61];
  assign t[3] = t[7] ? t[8] : t[152];
  assign t[40] = t[62] ^ t[63];
  assign t[41] = t[64] & t[65];
  assign t[42] = t[153] ^ t[66];
  assign t[43] = t[67] ^ t[19];
  assign t[44] = t[68] & t[69];
  assign t[45] = ~(t[70] & t[71]);
  assign t[46] = t[160] | t[72];
  assign t[47] = ~(t[73]);
  assign t[48] = ~(t[161]);
  assign t[49] = ~(t[74] & t[162]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[157] ^ t[75];
  assign t[51] = t[7] ? t[76] : t[163];
  assign t[52] = ~(t[14]);
  assign t[53] = t[158] ^ t[77];
  assign t[54] = t[159] ^ t[78];
  assign t[55] = t[79] ^ t[80];
  assign t[56] = t[35] ^ t[81];
  assign t[57] = t[52] ? t[82] : t[164];
  assign t[58] = t[83];
  assign t[59] = ~t[84];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[85] ^ t[86];
  assign t[61] = t[87] & t[88];
  assign t[62] = t[52] ? t[89] : t[165];
  assign t[63] = t[154] ^ t[90];
  assign t[64] = ~(t[40] ^ t[91]);
  assign t[65] = t[92] ^ t[93];
  assign t[66] = t[27] ? x[47] : x[46];
  assign t[67] = t[94] & t[95];
  assign t[68] = ~(t[96] ^ t[43]);
  assign t[69] = t[97] ^ t[3];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[72] & t[98]);
  assign t[71] = ~(t[166] ^ t[99]);
  assign t[72] = ~(t[100] & t[101]);
  assign t[73] = ~(t[46]);
  assign t[74] = ~(t[167]);
  assign t[75] = t[27] ? x[55] : x[54];
  assign t[76] = t[163] ^ t[102];
  assign t[77] = t[103] ? x[57] : x[56];
  assign t[78] = t[103] ? x[59] : x[58];
  assign t[79] = t[104] & t[105];
  assign t[7] = ~(t[14]);
  assign t[80] = t[106] & t[57];
  assign t[81] = t[52] ? t[107] : t[168];
  assign t[82] = t[164] ^ t[108];
  assign t[83] = t[26] ? t[109] : t[169];
  assign t[84] = t[26] ? t[110] : t[170];
  assign t[85] = t[111] & t[112];
  assign t[86] = t[113] & t[114];
  assign t[87] = ~(t[85] ^ t[115]);
  assign t[88] = t[116] ^ t[117];
  assign t[89] = t[165] ^ t[118];
  assign t[8] = t[152] ^ t[15];
  assign t[90] = t[26] ? t[119] : t[171];
  assign t[91] = t[120] ^ t[121];
  assign t[92] = t[63] ^ t[122];
  assign t[93] = t[155] ^ t[123];
  assign t[94] = ~(t[124]);
  assign t[95] = ~(t[32]);
  assign t[96] = t[32] ^ t[51];
  assign t[97] = t[51] ^ t[24];
  assign t[98] = ~(t[125] & t[126]);
  assign t[99] = t[127] ^ t[172];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind116(x, y);
 input [111:0] x;
 output y;

 wire [214:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[65] ^ t[24];
  assign t[101] = ~(t[131] & t[132]);
  assign t[102] = t[133] ^ t[181];
  assign t[103] = ~(t[177]);
  assign t[104] = t[134] & t[133];
  assign t[105] = ~(t[48]);
  assign t[106] = ~(t[135]);
  assign t[107] = ~(t[55]);
  assign t[108] = t[55] ^ t[81];
  assign t[109] = t[81] ^ t[32];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[105] ? x[68] : x[67];
  assign t[111] = t[179] ^ t[136];
  assign t[112] = t[105] ? x[70] : x[69];
  assign t[113] = t[26] ? t[137] : t[182];
  assign t[114] = t[26] ? t[138] : t[183];
  assign t[115] = t[139] ^ t[140];
  assign t[116] = t[84] ^ t[141];
  assign t[117] = t[142];
  assign t[118] = t[27] ? x[78] : x[77];
  assign t[119] = ~(t[143] ^ t[62]);
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[38] ^ t[124];
  assign t[121] = ~(t[127]);
  assign t[122] = ~(t[144]);
  assign t[123] = ~(t[3]);
  assign t[124] = t[7] ? t[145] : t[184];
  assign t[125] = t[38] ^ t[144];
  assign t[126] = t[144] ^ t[60];
  assign t[127] = t[124] ^ t[3];
  assign t[128] = t[180] ^ t[146];
  assign t[129] = t[147] ? x[83] : x[82];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[42] ^ t[65];
  assign t[131] = ~(t[134] | t[133]);
  assign t[132] = ~(t[148] | t[103]);
  assign t[133] = ~(t[185]);
  assign t[134] = ~(t[181]);
  assign t[135] = t[57] ^ t[81];
  assign t[136] = t[105] ? x[88] : x[87];
  assign t[137] = t[182] ^ t[149];
  assign t[138] = t[183] ^ t[150];
  assign t[139] = t[151] & t[152];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[153] & t[117];
  assign t[141] = ~t[154];
  assign t[142] = t[26] ? t[155] : t[186];
  assign t[143] = t[144] ^ t[3];
  assign t[144] = t[7] ? t[156] : t[187];
  assign t[145] = t[184] ^ t[157];
  assign t[146] = t[147] ? x[96] : x[95];
  assign t[147] = ~(t[48]);
  assign t[148] = ~(t[171]);
  assign t[149] = t[74] ? x[98] : x[97];
  assign t[14] = ~(t[26]);
  assign t[150] = t[147] ? x[100] : x[99];
  assign t[151] = ~(t[158]);
  assign t[152] = ~(t[83]);
  assign t[153] = ~(t[84]);
  assign t[154] = t[26] ? t[159] : t[188];
  assign t[155] = t[186] ^ t[160];
  assign t[156] = t[187] ^ t[161];
  assign t[157] = t[27] ? x[105] : x[104];
  assign t[158] = t[117] ^ t[84];
  assign t[159] = t[188] ^ t[162];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[105] ? x[107] : x[106];
  assign t[161] = t[27] ? x[109] : x[108];
  assign t[162] = t[74] ? x[111] : x[110];
  assign t[163] = t[189] ^ x[4];
  assign t[164] = t[190] ^ x[9];
  assign t[165] = t[191] ^ x[12];
  assign t[166] = t[192] ^ x[15];
  assign t[167] = t[193] ^ x[18];
  assign t[168] = t[194] ^ x[21];
  assign t[169] = t[195] ^ x[24];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[196] ^ x[27];
  assign t[171] = t[197] ^ x[30];
  assign t[172] = t[198] ^ x[33];
  assign t[173] = t[199] ^ x[36];
  assign t[174] = t[200] ^ x[39];
  assign t[175] = t[201] ^ x[42];
  assign t[176] = t[202] ^ x[45];
  assign t[177] = t[203] ^ x[48];
  assign t[178] = t[204] ^ x[51];
  assign t[179] = t[205] ^ x[56];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[206] ^ x[61];
  assign t[181] = t[207] ^ x[66];
  assign t[182] = t[208] ^ x[73];
  assign t[183] = t[209] ^ x[76];
  assign t[184] = t[210] ^ x[81];
  assign t[185] = t[211] ^ x[86];
  assign t[186] = t[212] ^ x[91];
  assign t[187] = t[213] ^ x[94];
  assign t[188] = t[214] ^ x[103];
  assign t[189] = (x[2] & x[3]);
  assign t[18] = t[32] ^ t[33];
  assign t[190] = (x[7] & x[8]);
  assign t[191] = (x[10] & x[11]);
  assign t[192] = (x[13] & x[14]);
  assign t[193] = (x[16] & x[17]);
  assign t[194] = (x[19] & x[20]);
  assign t[195] = (x[22] & x[23]);
  assign t[196] = (x[25] & x[26]);
  assign t[197] = (x[28] & x[29]);
  assign t[198] = (x[31] & x[32]);
  assign t[199] = (x[34] & x[35]);
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[37] & x[38]);
  assign t[201] = (x[40] & x[41]);
  assign t[202] = (x[43] & x[44]);
  assign t[203] = (x[46] & x[47]);
  assign t[204] = (x[49] & x[50]);
  assign t[205] = (x[54] & x[55]);
  assign t[206] = (x[59] & x[60]);
  assign t[207] = (x[64] & x[65]);
  assign t[208] = (x[71] & x[72]);
  assign t[209] = (x[74] & x[75]);
  assign t[20] = ~(t[36] ^ t[37]);
  assign t[210] = (x[79] & x[80]);
  assign t[211] = (x[84] & x[85]);
  assign t[212] = (x[89] & x[90]);
  assign t[213] = (x[92] & x[93]);
  assign t[214] = (x[101] & x[102]);
  assign t[21] = t[38] ^ t[39];
  assign t[22] = t[40] ^ t[24];
  assign t[23] = t[41] & t[42];
  assign t[24] = t[164] ^ t[43];
  assign t[25] = t[44] ^ t[45];
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[165]);
  assign t[29] = ~(t[166]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[167]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[51] ? t[52] : t[168];
  assign t[33] = t[53] ^ t[54];
  assign t[34] = t[55] ^ t[32];
  assign t[35] = t[56] & t[57];
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[3] ^ t[60];
  assign t[39] = t[62] ^ t[63];
  assign t[3] = t[7] ? t[8] : t[163];
  assign t[40] = t[51] ? t[64] : t[169];
  assign t[41] = ~(t[65]);
  assign t[42] = t[166] ^ t[66];
  assign t[43] = t[51] ? t[67] : t[170];
  assign t[44] = t[68] ^ t[23];
  assign t[45] = t[69] & t[70];
  assign t[46] = ~(t[71] & t[72]);
  assign t[47] = t[171] | t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = ~(t[172]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[75] & t[164]);
  assign t[51] = ~(t[14]);
  assign t[52] = t[168] ^ t[76];
  assign t[53] = t[77] ^ t[35];
  assign t[54] = t[78] & t[79];
  assign t[55] = t[51] ? t[80] : t[173];
  assign t[56] = ~(t[81]);
  assign t[57] = t[51] ? t[82] : t[174];
  assign t[58] = t[83] ^ t[84];
  assign t[59] = t[85] & t[86];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[7] ? t[87] : t[175];
  assign t[61] = t[62] ^ t[88];
  assign t[62] = t[89] ^ t[90];
  assign t[63] = t[91] & t[92];
  assign t[64] = t[169] ^ t[93];
  assign t[65] = t[165] ^ t[94];
  assign t[66] = t[51] ? t[95] : t[176];
  assign t[67] = t[170] ^ t[96];
  assign t[68] = t[97] & t[98];
  assign t[69] = ~(t[99] ^ t[44]);
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[100] ^ t[42];
  assign t[71] = ~(t[73] & t[101]);
  assign t[72] = ~(t[177] ^ t[102]);
  assign t[73] = ~(t[103] & t[104]);
  assign t[74] = ~(t[47]);
  assign t[75] = ~(t[178]);
  assign t[76] = t[105] ? x[53] : x[52];
  assign t[77] = t[106] & t[107];
  assign t[78] = ~(t[108] ^ t[53]);
  assign t[79] = t[109] ^ t[57];
  assign t[7] = ~(t[14]);
  assign t[80] = t[173] ^ t[110];
  assign t[81] = t[51] ? t[111] : t[179];
  assign t[82] = t[174] ^ t[112];
  assign t[83] = ~t[113];
  assign t[84] = t[114];
  assign t[85] = ~(t[58] ^ t[115]);
  assign t[86] = t[116] ^ t[117];
  assign t[87] = t[175] ^ t[118];
  assign t[88] = t[119] & t[120];
  assign t[89] = t[121] & t[122];
  assign t[8] = t[163] ^ t[15];
  assign t[90] = t[123] & t[124];
  assign t[91] = ~(t[89] ^ t[125]);
  assign t[92] = t[126] ^ t[127];
  assign t[93] = t[74] ? x[58] : x[57];
  assign t[94] = t[26] ? t[128] : t[180];
  assign t[95] = t[176] ^ t[129];
  assign t[96] = t[74] ? x[63] : x[62];
  assign t[97] = ~(t[130]);
  assign t[98] = ~(t[40]);
  assign t[99] = t[40] ^ t[65];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind117(x, y);
 input [111:0] x;
 output y;

 wire [192:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[117] ^ t[24];
  assign t[101] = ~(t[119] & t[120]);
  assign t[102] = t[121] ^ t[159];
  assign t[103] = ~(t[154]);
  assign t[104] = t[122] & t[121];
  assign t[105] = t[7] ? t[123] : t[160];
  assign t[106] = t[156] ^ t[124];
  assign t[107] = t[73] ? x[71] : x[70];
  assign t[108] = t[73] ? x[73] : x[72];
  assign t[109] = t[157] ^ t[125];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[87] ? x[75] : x[74];
  assign t[111] = t[91] ^ t[113];
  assign t[112] = t[39] ? t[126] : t[161];
  assign t[113] = t[39] ? t[127] : t[162];
  assign t[114] = t[158] ^ t[128];
  assign t[115] = t[98] ^ t[117];
  assign t[116] = t[39] ? t[129] : t[163];
  assign t[117] = t[144] ^ t[130];
  assign t[118] = t[39] ? t[131] : t[164];
  assign t[119] = ~(t[122] | t[121]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = ~(t[132] | t[103]);
  assign t[121] = ~(t[165]);
  assign t[122] = ~(t[159]);
  assign t[123] = t[160] ^ t[133];
  assign t[124] = t[27] ? x[92] : x[91];
  assign t[125] = t[134] ? x[94] : x[93];
  assign t[126] = t[161] ^ t[135];
  assign t[127] = t[162] ^ t[136];
  assign t[128] = t[87] ? x[96] : x[95];
  assign t[129] = t[163] ^ t[137];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[26] ? t[138] : t[166];
  assign t[131] = t[164] ^ t[139];
  assign t[132] = ~(t[149]);
  assign t[133] = t[27] ? x[101] : x[100];
  assign t[134] = ~(t[48]);
  assign t[135] = t[87] ? x[103] : x[102];
  assign t[136] = t[87] ? x[105] : x[104];
  assign t[137] = t[73] ? x[107] : x[106];
  assign t[138] = t[166] ^ t[140];
  assign t[139] = t[134] ? x[109] : x[108];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[134] ? x[111] : x[110];
  assign t[141] = t[167] ^ x[4];
  assign t[142] = t[168] ^ x[9];
  assign t[143] = t[169] ^ x[12];
  assign t[144] = t[170] ^ x[15];
  assign t[145] = t[171] ^ x[18];
  assign t[146] = t[172] ^ x[21];
  assign t[147] = t[173] ^ x[24];
  assign t[148] = t[174] ^ x[27];
  assign t[149] = t[175] ^ x[30];
  assign t[14] = ~(t[26]);
  assign t[150] = t[176] ^ x[33];
  assign t[151] = t[177] ^ x[36];
  assign t[152] = t[178] ^ x[39];
  assign t[153] = t[179] ^ x[42];
  assign t[154] = t[180] ^ x[47];
  assign t[155] = t[181] ^ x[50];
  assign t[156] = t[182] ^ x[55];
  assign t[157] = t[183] ^ x[58];
  assign t[158] = t[184] ^ x[61];
  assign t[159] = t[185] ^ x[66];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[186] ^ x[69];
  assign t[161] = t[187] ^ x[78];
  assign t[162] = t[188] ^ x[81];
  assign t[163] = t[189] ^ x[84];
  assign t[164] = t[190] ^ x[87];
  assign t[165] = t[191] ^ x[90];
  assign t[166] = t[192] ^ x[99];
  assign t[167] = (x[2] & x[3]);
  assign t[168] = (x[7] & x[8]);
  assign t[169] = (x[10] & x[11]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = (x[13] & x[14]);
  assign t[171] = (x[16] & x[17]);
  assign t[172] = (x[19] & x[20]);
  assign t[173] = (x[22] & x[23]);
  assign t[174] = (x[25] & x[26]);
  assign t[175] = (x[28] & x[29]);
  assign t[176] = (x[31] & x[32]);
  assign t[177] = (x[34] & x[35]);
  assign t[178] = (x[37] & x[38]);
  assign t[179] = (x[40] & x[41]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = (x[45] & x[46]);
  assign t[181] = (x[48] & x[49]);
  assign t[182] = (x[53] & x[54]);
  assign t[183] = (x[56] & x[57]);
  assign t[184] = (x[59] & x[60]);
  assign t[185] = (x[64] & x[65]);
  assign t[186] = (x[67] & x[68]);
  assign t[187] = (x[76] & x[77]);
  assign t[188] = (x[79] & x[80]);
  assign t[189] = (x[82] & x[83]);
  assign t[18] = t[32] ^ t[3];
  assign t[190] = (x[85] & x[86]);
  assign t[191] = (x[88] & x[89]);
  assign t[192] = (x[97] & x[98]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = ~(t[4]);
  assign t[20] = t[35] ^ t[36];
  assign t[21] = t[37] & t[38];
  assign t[22] = t[39] ? t[40] : t[142];
  assign t[23] = t[41] ^ t[42];
  assign t[24] = t[143] ^ t[43];
  assign t[25] = t[44] ^ t[45];
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[144]);
  assign t[29] = ~(t[145]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[146]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[7] ? t[51] : t[147];
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[54] & t[55];
  assign t[35] = ~t[56];
  assign t[36] = ~t[57];
  assign t[37] = ~(t[58]);
  assign t[38] = t[59];
  assign t[39] = ~(t[14]);
  assign t[3] = t[7] ? t[8] : t[141];
  assign t[40] = t[142] ^ t[60];
  assign t[41] = t[61] ^ t[62];
  assign t[42] = t[63] & t[64];
  assign t[43] = t[39] ? t[65] : t[148];
  assign t[44] = t[66] ^ t[67];
  assign t[45] = t[68] & t[69];
  assign t[46] = ~(t[70] & t[71]);
  assign t[47] = t[149] | t[72];
  assign t[48] = ~(t[73]);
  assign t[49] = ~(t[150]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[74] & t[143]);
  assign t[51] = t[147] ^ t[75];
  assign t[52] = t[76] & t[77];
  assign t[53] = t[78] & t[79];
  assign t[54] = ~(t[52] ^ t[80]);
  assign t[55] = t[81] ^ t[82];
  assign t[56] = t[26] ? t[83] : t[151];
  assign t[57] = t[26] ? t[84] : t[152];
  assign t[58] = t[85];
  assign t[59] = t[26] ? t[86] : t[153];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[87] ? x[44] : x[43];
  assign t[61] = t[88] & t[89];
  assign t[62] = t[90] & t[91];
  assign t[63] = ~(t[92] ^ t[41]);
  assign t[64] = t[93] ^ t[91];
  assign t[65] = t[148] ^ t[94];
  assign t[66] = t[95] & t[96];
  assign t[67] = t[97] & t[98];
  assign t[68] = ~(t[99] ^ t[44]);
  assign t[69] = t[100] ^ t[98];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[72] & t[101]);
  assign t[71] = ~(t[154] ^ t[102]);
  assign t[72] = ~(t[103] & t[104]);
  assign t[73] = ~(t[47]);
  assign t[74] = ~(t[155]);
  assign t[75] = t[27] ? x[52] : x[51];
  assign t[76] = ~(t[82]);
  assign t[77] = ~(t[105]);
  assign t[78] = ~(t[32]);
  assign t[79] = t[7] ? t[106] : t[156];
  assign t[7] = ~(t[14]);
  assign t[80] = t[18] ^ t[105];
  assign t[81] = t[105] ^ t[3];
  assign t[82] = t[79] ^ t[32];
  assign t[83] = t[151] ^ t[107];
  assign t[84] = t[152] ^ t[108];
  assign t[85] = t[26] ? t[109] : t[157];
  assign t[86] = t[153] ^ t[110];
  assign t[87] = ~(t[48]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[112]);
  assign t[8] = t[141] ^ t[15];
  assign t[90] = ~(t[113]);
  assign t[91] = t[39] ? t[114] : t[158];
  assign t[92] = t[112] ^ t[113];
  assign t[93] = t[113] ^ t[22];
  assign t[94] = t[73] ? x[63] : x[62];
  assign t[95] = ~(t[115]);
  assign t[96] = ~(t[116]);
  assign t[97] = ~(t[117]);
  assign t[98] = t[145] ^ t[118];
  assign t[99] = t[116] ^ t[117];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind118(x, y);
 input [111:0] x;
 output y;

 wire [202:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[165] ^ t[127];
  assign t[101] = t[166] ^ t[128];
  assign t[102] = ~(t[108]);
  assign t[103] = ~(t[129]);
  assign t[104] = ~(t[50]);
  assign t[105] = t[130];
  assign t[106] = t[32] ^ t[129];
  assign t[107] = t[129] ^ t[51];
  assign t[108] = t[105] ^ t[50];
  assign t[109] = ~(t[131]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = ~(t[132]);
  assign t[111] = ~(t[133]);
  assign t[112] = t[54] ? t[134] : t[171];
  assign t[113] = t[132] ^ t[133];
  assign t[114] = t[133] ^ t[34];
  assign t[115] = ~(t[135]);
  assign t[116] = ~(t[3]);
  assign t[117] = ~(t[36]);
  assign t[118] = t[167] ^ t[136];
  assign t[119] = t[27] ? x[76] : x[75];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = ~(t[47]);
  assign t[121] = t[168] ^ t[137];
  assign t[122] = t[169] ^ t[138];
  assign t[123] = ~(t[126] | t[125]);
  assign t[124] = ~(t[139] | t[98]);
  assign t[125] = ~(t[172]);
  assign t[126] = ~(t[170]);
  assign t[127] = t[120] ? x[81] : x[80];
  assign t[128] = t[74] ? x[83] : x[82];
  assign t[129] = t[140];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[54] ? t[141] : t[173];
  assign t[131] = t[112] ^ t[133];
  assign t[132] = t[54] ? t[142] : t[174];
  assign t[133] = t[54] ? t[143] : t[175];
  assign t[134] = t[171] ^ t[144];
  assign t[135] = t[61] ^ t[36];
  assign t[136] = t[27] ? x[94] : x[93];
  assign t[137] = t[120] ? x[96] : x[95];
  assign t[138] = t[120] ? x[98] : x[97];
  assign t[139] = ~(t[160]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[54] ? t[145] : t[176];
  assign t[141] = t[173] ^ t[146];
  assign t[142] = t[174] ^ t[147];
  assign t[143] = t[175] ^ t[148];
  assign t[144] = t[149] ? x[103] : x[102];
  assign t[145] = t[176] ^ t[150];
  assign t[146] = t[74] ? x[105] : x[104];
  assign t[147] = t[149] ? x[107] : x[106];
  assign t[148] = t[149] ? x[109] : x[108];
  assign t[149] = ~(t[47]);
  assign t[14] = ~(t[26]);
  assign t[150] = t[74] ? x[111] : x[110];
  assign t[151] = t[177] ^ x[4];
  assign t[152] = t[178] ^ x[9];
  assign t[153] = t[179] ^ x[12];
  assign t[154] = t[180] ^ x[15];
  assign t[155] = t[181] ^ x[18];
  assign t[156] = t[182] ^ x[21];
  assign t[157] = t[183] ^ x[24];
  assign t[158] = t[184] ^ x[27];
  assign t[159] = t[185] ^ x[30];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[186] ^ x[33];
  assign t[161] = t[187] ^ x[36];
  assign t[162] = t[188] ^ x[39];
  assign t[163] = t[189] ^ x[42];
  assign t[164] = t[190] ^ x[45];
  assign t[165] = t[191] ^ x[48];
  assign t[166] = t[192] ^ x[51];
  assign t[167] = t[193] ^ x[58];
  assign t[168] = t[194] ^ x[65];
  assign t[169] = t[195] ^ x[68];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[196] ^ x[71];
  assign t[171] = t[197] ^ x[74];
  assign t[172] = t[198] ^ x[79];
  assign t[173] = t[199] ^ x[86];
  assign t[174] = t[200] ^ x[89];
  assign t[175] = t[201] ^ x[92];
  assign t[176] = t[202] ^ x[101];
  assign t[177] = (x[2] & x[3]);
  assign t[178] = (x[7] & x[8]);
  assign t[179] = (x[10] & x[11]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = (x[13] & x[14]);
  assign t[181] = (x[16] & x[17]);
  assign t[182] = (x[19] & x[20]);
  assign t[183] = (x[22] & x[23]);
  assign t[184] = (x[25] & x[26]);
  assign t[185] = (x[28] & x[29]);
  assign t[186] = (x[31] & x[32]);
  assign t[187] = (x[34] & x[35]);
  assign t[188] = (x[37] & x[38]);
  assign t[189] = (x[40] & x[41]);
  assign t[18] = t[32] ^ t[33];
  assign t[190] = (x[43] & x[44]);
  assign t[191] = (x[46] & x[47]);
  assign t[192] = (x[49] & x[50]);
  assign t[193] = (x[56] & x[57]);
  assign t[194] = (x[63] & x[64]);
  assign t[195] = (x[66] & x[67]);
  assign t[196] = (x[69] & x[70]);
  assign t[197] = (x[72] & x[73]);
  assign t[198] = (x[77] & x[78]);
  assign t[199] = (x[84] & x[85]);
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[87] & x[88]);
  assign t[201] = (x[90] & x[91]);
  assign t[202] = (x[99] & x[100]);
  assign t[20] = t[3] ^ t[36];
  assign t[21] = t[37] & t[38];
  assign t[22] = t[152] ^ t[39];
  assign t[23] = t[153] ^ t[40];
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[43] & t[44];
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[154]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[152]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = t[50] ^ t[51];
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[54] ? t[55] : t[156];
  assign t[35] = t[56] ^ t[57];
  assign t[36] = t[7] ? t[58] : t[157];
  assign t[37] = ~(t[20] ^ t[59]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[54] ? t[62] : t[158];
  assign t[3] = t[7] ? t[8] : t[151];
  assign t[40] = t[54] ? t[63] : t[159];
  assign t[41] = t[64] & t[65];
  assign t[42] = t[66] & t[67];
  assign t[43] = ~(t[41] ^ t[68]);
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[71] & t[72]);
  assign t[46] = t[160] | t[73];
  assign t[47] = ~(t[74]);
  assign t[48] = ~(t[153]);
  assign t[49] = ~(t[75] & t[161]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~t[76];
  assign t[51] = t[77];
  assign t[52] = t[78] ^ t[79];
  assign t[53] = t[80] & t[81];
  assign t[54] = ~(t[14]);
  assign t[55] = t[156] ^ t[82];
  assign t[56] = t[83] ^ t[84];
  assign t[57] = t[85] & t[86];
  assign t[58] = t[157] ^ t[87];
  assign t[59] = t[88] ^ t[89];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[36] ^ t[90];
  assign t[61] = t[7] ? t[91] : t[162];
  assign t[62] = t[158] ^ t[92];
  assign t[63] = t[159] ^ t[93];
  assign t[64] = ~(t[70]);
  assign t[65] = ~(t[94]);
  assign t[66] = ~(t[22]);
  assign t[67] = t[163] ^ t[95];
  assign t[68] = t[12] ^ t[94];
  assign t[69] = t[94] ^ t[23];
  assign t[6] = t[12] ^ t[13];
  assign t[70] = t[67] ^ t[22];
  assign t[71] = ~(t[73] & t[96]);
  assign t[72] = ~(t[164] ^ t[97]);
  assign t[73] = ~(t[98] & t[99]);
  assign t[74] = ~(t[46]);
  assign t[75] = ~(t[163]);
  assign t[76] = t[54] ? t[100] : t[165];
  assign t[77] = t[54] ? t[101] : t[166];
  assign t[78] = t[102] & t[103];
  assign t[79] = t[104] & t[105];
  assign t[7] = ~(t[14]);
  assign t[80] = ~(t[78] ^ t[106]);
  assign t[81] = t[107] ^ t[108];
  assign t[82] = t[74] ? x[53] : x[52];
  assign t[83] = t[109] & t[110];
  assign t[84] = t[111] & t[112];
  assign t[85] = ~(t[113] ^ t[56]);
  assign t[86] = t[114] ^ t[112];
  assign t[87] = t[27] ? x[55] : x[54];
  assign t[88] = t[115] & t[116];
  assign t[89] = t[117] & t[61];
  assign t[8] = t[151] ^ t[15];
  assign t[90] = t[7] ? t[118] : t[167];
  assign t[91] = t[162] ^ t[119];
  assign t[92] = t[120] ? x[60] : x[59];
  assign t[93] = t[120] ? x[62] : x[61];
  assign t[94] = t[54] ? t[121] : t[168];
  assign t[95] = t[54] ? t[122] : t[169];
  assign t[96] = ~(t[123] & t[124]);
  assign t[97] = t[125] ^ t[170];
  assign t[98] = ~(t[164]);
  assign t[99] = t[126] & t[125];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind119(x, y);
 input [111:0] x;
 output y;

 wire [203:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[167]);
  assign t[101] = t[129] & t[128];
  assign t[102] = t[27] ? x[71] : x[70];
  assign t[103] = ~(t[47]);
  assign t[104] = t[103] ? x[73] : x[72];
  assign t[105] = ~(t[130]);
  assign t[106] = ~(t[34]);
  assign t[107] = ~(t[35]);
  assign t[108] = t[52] ? t[131] : t[172];
  assign t[109] = t[168] ^ t[132];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[133] ? x[78] : x[77];
  assign t[111] = t[73] ? x[80] : x[79];
  assign t[112] = ~(t[118]);
  assign t[113] = ~(t[134]);
  assign t[114] = ~(t[58]);
  assign t[115] = t[52] ? t[135] : t[173];
  assign t[116] = t[38] ^ t[134];
  assign t[117] = t[134] ^ t[59];
  assign t[118] = t[115] ^ t[58];
  assign t[119] = t[169] ^ t[136];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[170] ^ t[137];
  assign t[121] = t[138] & t[139];
  assign t[122] = t[140] & t[93];
  assign t[123] = t[141];
  assign t[124] = t[52] ? t[142] : t[174];
  assign t[125] = t[3] ^ t[51];
  assign t[126] = ~(t[129] | t[128]);
  assign t[127] = ~(t[143] | t[100]);
  assign t[128] = ~(t[175]);
  assign t[129] = ~(t[171]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[57] ^ t[35];
  assign t[131] = t[172] ^ t[144];
  assign t[132] = t[103] ? x[91] : x[90];
  assign t[133] = ~(t[47]);
  assign t[134] = t[52] ? t[145] : t[176];
  assign t[135] = t[173] ^ t[146];
  assign t[136] = t[73] ? x[96] : x[95];
  assign t[137] = t[103] ? x[98] : x[97];
  assign t[138] = ~(t[147]);
  assign t[139] = ~(t[62]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[63]);
  assign t[141] = t[52] ? t[148] : t[177];
  assign t[142] = t[174] ^ t[149];
  assign t[143] = ~(t[159]);
  assign t[144] = t[103] ? x[103] : x[102];
  assign t[145] = t[176] ^ t[150];
  assign t[146] = t[133] ? x[105] : x[104];
  assign t[147] = t[93] ^ t[63];
  assign t[148] = t[177] ^ t[151];
  assign t[149] = t[73] ? x[107] : x[106];
  assign t[14] = ~(t[26]);
  assign t[150] = t[133] ? x[109] : x[108];
  assign t[151] = t[73] ? x[111] : x[110];
  assign t[152] = t[178] ^ x[4];
  assign t[153] = t[179] ^ x[9];
  assign t[154] = t[180] ^ x[12];
  assign t[155] = t[181] ^ x[15];
  assign t[156] = t[182] ^ x[18];
  assign t[157] = t[183] ^ x[21];
  assign t[158] = t[184] ^ x[24];
  assign t[159] = t[185] ^ x[27];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[186] ^ x[30];
  assign t[161] = t[187] ^ x[33];
  assign t[162] = t[188] ^ x[36];
  assign t[163] = t[189] ^ x[39];
  assign t[164] = t[190] ^ x[42];
  assign t[165] = t[191] ^ x[45];
  assign t[166] = t[192] ^ x[48];
  assign t[167] = t[193] ^ x[53];
  assign t[168] = t[194] ^ x[60];
  assign t[169] = t[195] ^ x[63];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[196] ^ x[66];
  assign t[171] = t[197] ^ x[69];
  assign t[172] = t[198] ^ x[76];
  assign t[173] = t[199] ^ x[83];
  assign t[174] = t[200] ^ x[86];
  assign t[175] = t[201] ^ x[89];
  assign t[176] = t[202] ^ x[94];
  assign t[177] = t[203] ^ x[101];
  assign t[178] = (x[2] & x[3]);
  assign t[179] = (x[7] & x[8]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = (x[10] & x[11]);
  assign t[181] = (x[13] & x[14]);
  assign t[182] = (x[16] & x[17]);
  assign t[183] = (x[19] & x[20]);
  assign t[184] = (x[22] & x[23]);
  assign t[185] = (x[25] & x[26]);
  assign t[186] = (x[28] & x[29]);
  assign t[187] = (x[31] & x[32]);
  assign t[188] = (x[34] & x[35]);
  assign t[189] = (x[37] & x[38]);
  assign t[18] = t[32] ^ t[24];
  assign t[190] = (x[40] & x[41]);
  assign t[191] = (x[43] & x[44]);
  assign t[192] = (x[46] & x[47]);
  assign t[193] = (x[51] & x[52]);
  assign t[194] = (x[58] & x[59]);
  assign t[195] = (x[61] & x[62]);
  assign t[196] = (x[64] & x[65]);
  assign t[197] = (x[67] & x[68]);
  assign t[198] = (x[74] & x[75]);
  assign t[199] = (x[81] & x[82]);
  assign t[19] = t[33] & t[3];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[84] & x[85]);
  assign t[201] = (x[87] & x[88]);
  assign t[202] = (x[92] & x[93]);
  assign t[203] = (x[99] & x[100]);
  assign t[20] = t[34] ^ t[35];
  assign t[21] = t[36] & t[37];
  assign t[22] = t[38] ^ t[39];
  assign t[23] = t[40] ^ t[41];
  assign t[24] = t[7] ? t[42] : t[153];
  assign t[25] = t[43] ^ t[44];
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[154]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[156]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = t[7] ? t[50] : t[157];
  assign t[33] = ~(t[51]);
  assign t[34] = t[52] ? t[53] : t[158];
  assign t[35] = t[156] ^ t[54];
  assign t[36] = ~(t[20] ^ t[55]);
  assign t[37] = t[56] ^ t[57];
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[60] ^ t[61];
  assign t[3] = t[7] ? t[8] : t[152];
  assign t[40] = t[62] ^ t[63];
  assign t[41] = t[64] & t[65];
  assign t[42] = t[153] ^ t[66];
  assign t[43] = t[67] ^ t[19];
  assign t[44] = t[68] & t[69];
  assign t[45] = ~(t[70] & t[71]);
  assign t[46] = t[159] | t[72];
  assign t[47] = ~(t[73]);
  assign t[48] = ~(t[160]);
  assign t[49] = ~(t[74] & t[161]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[157] ^ t[75];
  assign t[51] = t[7] ? t[76] : t[162];
  assign t[52] = ~(t[14]);
  assign t[53] = t[158] ^ t[77];
  assign t[54] = t[52] ? t[78] : t[163];
  assign t[55] = t[79] ^ t[80];
  assign t[56] = t[35] ^ t[81];
  assign t[57] = t[164] ^ t[82];
  assign t[58] = t[52] ? t[83] : t[165];
  assign t[59] = t[52] ? t[84] : t[166];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[85] ^ t[86];
  assign t[61] = t[87] & t[88];
  assign t[62] = t[89];
  assign t[63] = ~t[90];
  assign t[64] = ~(t[40] ^ t[91]);
  assign t[65] = t[92] ^ t[93];
  assign t[66] = t[27] ? x[50] : x[49];
  assign t[67] = t[94] & t[95];
  assign t[68] = ~(t[96] ^ t[43]);
  assign t[69] = t[97] ^ t[3];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[72] & t[98]);
  assign t[71] = ~(t[167] ^ t[99]);
  assign t[72] = ~(t[100] & t[101]);
  assign t[73] = ~(t[46]);
  assign t[74] = ~(t[164]);
  assign t[75] = t[27] ? x[55] : x[54];
  assign t[76] = t[162] ^ t[102];
  assign t[77] = t[103] ? x[57] : x[56];
  assign t[78] = t[163] ^ t[104];
  assign t[79] = t[105] & t[106];
  assign t[7] = ~(t[14]);
  assign t[80] = t[107] & t[57];
  assign t[81] = t[160] ^ t[108];
  assign t[82] = t[52] ? t[109] : t[168];
  assign t[83] = t[165] ^ t[110];
  assign t[84] = t[166] ^ t[111];
  assign t[85] = t[112] & t[113];
  assign t[86] = t[114] & t[115];
  assign t[87] = ~(t[85] ^ t[116]);
  assign t[88] = t[117] ^ t[118];
  assign t[89] = t[52] ? t[119] : t[169];
  assign t[8] = t[152] ^ t[15];
  assign t[90] = t[52] ? t[120] : t[170];
  assign t[91] = t[121] ^ t[122];
  assign t[92] = t[63] ^ t[123];
  assign t[93] = t[124];
  assign t[94] = ~(t[125]);
  assign t[95] = ~(t[32]);
  assign t[96] = t[32] ^ t[51];
  assign t[97] = t[51] ^ t[24];
  assign t[98] = ~(t[126] & t[127]);
  assign t[99] = t[128] ^ t[171];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind120(x, y);
 input [111:0] x;
 output y;

 wire [214:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[64] ^ t[24];
  assign t[101] = ~(t[132] & t[133]);
  assign t[102] = t[134] ^ t[182];
  assign t[103] = ~(t[177]);
  assign t[104] = t[135] & t[134];
  assign t[105] = t[136] ? x[67] : x[66];
  assign t[106] = ~(t[137]);
  assign t[107] = ~(t[54]);
  assign t[108] = t[54] ^ t[81];
  assign t[109] = t[81] ^ t[32];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[136] ? x[69] : x[68];
  assign t[111] = t[66] ? t[138] : t[183];
  assign t[112] = t[178] ^ t[139];
  assign t[113] = t[179] ^ t[140];
  assign t[114] = t[180] ^ t[141];
  assign t[115] = t[142] ^ t[143];
  assign t[116] = t[84] ^ t[144];
  assign t[117] = t[66] ? t[145] : t[184];
  assign t[118] = t[27] ? x[77] : x[76];
  assign t[119] = ~(t[146] ^ t[61]);
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[38] ^ t[124];
  assign t[121] = ~(t[127]);
  assign t[122] = ~(t[147]);
  assign t[123] = ~(t[3]);
  assign t[124] = t[7] ? t[148] : t[185];
  assign t[125] = t[38] ^ t[147];
  assign t[126] = t[147] ^ t[59];
  assign t[127] = t[124] ^ t[3];
  assign t[128] = t[74] ? x[82] : x[81];
  assign t[129] = t[181] ^ t[149];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[74] ? x[84] : x[83];
  assign t[131] = t[42] ^ t[64];
  assign t[132] = ~(t[135] | t[134]);
  assign t[133] = ~(t[150] | t[103]);
  assign t[134] = ~(t[186]);
  assign t[135] = ~(t[182]);
  assign t[136] = ~(t[48]);
  assign t[137] = t[56] ^ t[81];
  assign t[138] = t[183] ^ t[151];
  assign t[139] = t[136] ? x[89] : x[88];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[152] ? x[91] : x[90];
  assign t[141] = t[152] ? x[93] : x[92];
  assign t[142] = t[153] & t[154];
  assign t[143] = t[155] & t[117];
  assign t[144] = t[66] ? t[156] : t[187];
  assign t[145] = t[184] ^ t[157];
  assign t[146] = t[147] ^ t[3];
  assign t[147] = t[7] ? t[158] : t[188];
  assign t[148] = t[185] ^ t[159];
  assign t[149] = t[136] ? x[101] : x[100];
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[169]);
  assign t[151] = t[136] ? x[103] : x[102];
  assign t[152] = ~(t[48]);
  assign t[153] = ~(t[160]);
  assign t[154] = ~(t[83]);
  assign t[155] = ~(t[84]);
  assign t[156] = t[187] ^ t[161];
  assign t[157] = t[152] ? x[105] : x[104];
  assign t[158] = t[188] ^ t[162];
  assign t[159] = t[27] ? x[107] : x[106];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[117] ^ t[84];
  assign t[161] = t[74] ? x[109] : x[108];
  assign t[162] = t[27] ? x[111] : x[110];
  assign t[163] = t[189] ^ x[4];
  assign t[164] = t[190] ^ x[9];
  assign t[165] = t[191] ^ x[12];
  assign t[166] = t[192] ^ x[15];
  assign t[167] = t[193] ^ x[18];
  assign t[168] = t[194] ^ x[21];
  assign t[169] = t[195] ^ x[24];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[196] ^ x[27];
  assign t[171] = t[197] ^ x[30];
  assign t[172] = t[198] ^ x[33];
  assign t[173] = t[199] ^ x[36];
  assign t[174] = t[200] ^ x[39];
  assign t[175] = t[201] ^ x[42];
  assign t[176] = t[202] ^ x[45];
  assign t[177] = t[203] ^ x[48];
  assign t[178] = t[204] ^ x[51];
  assign t[179] = t[205] ^ x[54];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[206] ^ x[57];
  assign t[181] = t[207] ^ x[60];
  assign t[182] = t[208] ^ x[65];
  assign t[183] = t[209] ^ x[72];
  assign t[184] = t[210] ^ x[75];
  assign t[185] = t[211] ^ x[80];
  assign t[186] = t[212] ^ x[87];
  assign t[187] = t[213] ^ x[96];
  assign t[188] = t[214] ^ x[99];
  assign t[189] = (x[2] & x[3]);
  assign t[18] = t[32] ^ t[33];
  assign t[190] = (x[7] & x[8]);
  assign t[191] = (x[10] & x[11]);
  assign t[192] = (x[13] & x[14]);
  assign t[193] = (x[16] & x[17]);
  assign t[194] = (x[19] & x[20]);
  assign t[195] = (x[22] & x[23]);
  assign t[196] = (x[25] & x[26]);
  assign t[197] = (x[28] & x[29]);
  assign t[198] = (x[31] & x[32]);
  assign t[199] = (x[34] & x[35]);
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[37] & x[38]);
  assign t[201] = (x[40] & x[41]);
  assign t[202] = (x[43] & x[44]);
  assign t[203] = (x[46] & x[47]);
  assign t[204] = (x[49] & x[50]);
  assign t[205] = (x[52] & x[53]);
  assign t[206] = (x[55] & x[56]);
  assign t[207] = (x[58] & x[59]);
  assign t[208] = (x[63] & x[64]);
  assign t[209] = (x[70] & x[71]);
  assign t[20] = ~(t[36] ^ t[37]);
  assign t[210] = (x[73] & x[74]);
  assign t[211] = (x[78] & x[79]);
  assign t[212] = (x[85] & x[86]);
  assign t[213] = (x[94] & x[95]);
  assign t[214] = (x[97] & x[98]);
  assign t[21] = t[38] ^ t[39];
  assign t[22] = t[40] ^ t[24];
  assign t[23] = t[41] & t[42];
  assign t[24] = t[43];
  assign t[25] = t[44] ^ t[45];
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[164]);
  assign t[29] = ~(t[165]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[166]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[167] ^ t[51];
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[54] ^ t[32];
  assign t[35] = t[55] & t[56];
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[3] ^ t[59];
  assign t[39] = t[61] ^ t[62];
  assign t[3] = t[7] ? t[8] : t[163];
  assign t[40] = t[63];
  assign t[41] = ~(t[64]);
  assign t[42] = t[65];
  assign t[43] = t[66] ? t[67] : t[168];
  assign t[44] = t[68] ^ t[23];
  assign t[45] = t[69] & t[70];
  assign t[46] = ~(t[71] & t[72]);
  assign t[47] = t[169] | t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = ~(t[167]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[75] & t[170]);
  assign t[51] = t[66] ? t[76] : t[171];
  assign t[52] = t[77] ^ t[35];
  assign t[53] = t[78] & t[79];
  assign t[54] = t[66] ? t[80] : t[172];
  assign t[55] = ~(t[81]);
  assign t[56] = t[173] ^ t[82];
  assign t[57] = t[83] ^ t[84];
  assign t[58] = t[85] & t[86];
  assign t[59] = t[7] ? t[87] : t[174];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[61] ^ t[88];
  assign t[61] = t[89] ^ t[90];
  assign t[62] = t[91] & t[92];
  assign t[63] = t[66] ? t[93] : t[175];
  assign t[64] = ~t[94];
  assign t[65] = t[66] ? t[95] : t[176];
  assign t[66] = ~(t[14]);
  assign t[67] = t[168] ^ t[96];
  assign t[68] = t[97] & t[98];
  assign t[69] = ~(t[99] ^ t[44]);
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[100] ^ t[42];
  assign t[71] = ~(t[73] & t[101]);
  assign t[72] = ~(t[177] ^ t[102]);
  assign t[73] = ~(t[103] & t[104]);
  assign t[74] = ~(t[47]);
  assign t[75] = ~(t[173]);
  assign t[76] = t[171] ^ t[105];
  assign t[77] = t[106] & t[107];
  assign t[78] = ~(t[108] ^ t[52]);
  assign t[79] = t[109] ^ t[56];
  assign t[7] = ~(t[14]);
  assign t[80] = t[172] ^ t[110];
  assign t[81] = t[166] ^ t[111];
  assign t[82] = t[66] ? t[112] : t[178];
  assign t[83] = t[66] ? t[113] : t[179];
  assign t[84] = t[66] ? t[114] : t[180];
  assign t[85] = ~(t[57] ^ t[115]);
  assign t[86] = t[116] ^ t[117];
  assign t[87] = t[174] ^ t[118];
  assign t[88] = t[119] & t[120];
  assign t[89] = t[121] & t[122];
  assign t[8] = t[163] ^ t[15];
  assign t[90] = t[123] & t[124];
  assign t[91] = ~(t[89] ^ t[125]);
  assign t[92] = t[126] ^ t[127];
  assign t[93] = t[175] ^ t[128];
  assign t[94] = t[66] ? t[129] : t[181];
  assign t[95] = t[176] ^ t[130];
  assign t[96] = t[74] ? x[62] : x[61];
  assign t[97] = ~(t[131]);
  assign t[98] = ~(t[40]);
  assign t[99] = t[40] ^ t[64];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind121(x, y);
 input [111:0] x;
 output y;

 wire [192:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[116] ^ t[24];
  assign t[101] = ~(t[118] & t[119]);
  assign t[102] = t[120] ^ t[158];
  assign t[103] = ~(t[155]);
  assign t[104] = t[121] & t[120];
  assign t[105] = t[7] ? t[122] : t[159];
  assign t[106] = t[157] ^ t[123];
  assign t[107] = ~(t[47]);
  assign t[108] = t[107] ? x[74] : x[73];
  assign t[109] = ~(t[47]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[91] ^ t[112];
  assign t[111] = t[55] ? t[124] : t[160];
  assign t[112] = t[145] ^ t[125];
  assign t[113] = t[55] ? t[126] : t[161];
  assign t[114] = t[98] ^ t[116];
  assign t[115] = t[127];
  assign t[116] = ~t[128];
  assign t[117] = t[55] ? t[129] : t[162];
  assign t[118] = ~(t[121] | t[120]);
  assign t[119] = ~(t[130] | t[103]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = ~(t[163]);
  assign t[121] = ~(t[158]);
  assign t[122] = t[159] ^ t[131];
  assign t[123] = t[27] ? x[88] : x[87];
  assign t[124] = t[160] ^ t[132];
  assign t[125] = t[55] ? t[133] : t[164];
  assign t[126] = t[161] ^ t[134];
  assign t[127] = t[55] ? t[135] : t[165];
  assign t[128] = t[55] ? t[136] : t[166];
  assign t[129] = t[162] ^ t[137];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = ~(t[152]);
  assign t[131] = t[27] ? x[99] : x[98];
  assign t[132] = t[109] ? x[101] : x[100];
  assign t[133] = t[164] ^ t[138];
  assign t[134] = t[109] ? x[103] : x[102];
  assign t[135] = t[165] ^ t[139];
  assign t[136] = t[166] ^ t[140];
  assign t[137] = t[73] ? x[105] : x[104];
  assign t[138] = t[109] ? x[107] : x[106];
  assign t[139] = t[73] ? x[109] : x[108];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[109] ? x[111] : x[110];
  assign t[141] = t[167] ^ x[4];
  assign t[142] = t[168] ^ x[9];
  assign t[143] = t[169] ^ x[12];
  assign t[144] = t[170] ^ x[15];
  assign t[145] = t[171] ^ x[18];
  assign t[146] = t[172] ^ x[21];
  assign t[147] = t[173] ^ x[24];
  assign t[148] = t[174] ^ x[27];
  assign t[149] = t[175] ^ x[30];
  assign t[14] = ~(t[26]);
  assign t[150] = t[176] ^ x[33];
  assign t[151] = t[177] ^ x[36];
  assign t[152] = t[178] ^ x[39];
  assign t[153] = t[179] ^ x[42];
  assign t[154] = t[180] ^ x[45];
  assign t[155] = t[181] ^ x[48];
  assign t[156] = t[182] ^ x[51];
  assign t[157] = t[183] ^ x[56];
  assign t[158] = t[184] ^ x[69];
  assign t[159] = t[185] ^ x[72];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[186] ^ x[77];
  assign t[161] = t[187] ^ x[80];
  assign t[162] = t[188] ^ x[83];
  assign t[163] = t[189] ^ x[86];
  assign t[164] = t[190] ^ x[91];
  assign t[165] = t[191] ^ x[94];
  assign t[166] = t[192] ^ x[97];
  assign t[167] = (x[2] & x[3]);
  assign t[168] = (x[7] & x[8]);
  assign t[169] = (x[10] & x[11]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = (x[13] & x[14]);
  assign t[171] = (x[16] & x[17]);
  assign t[172] = (x[19] & x[20]);
  assign t[173] = (x[22] & x[23]);
  assign t[174] = (x[25] & x[26]);
  assign t[175] = (x[28] & x[29]);
  assign t[176] = (x[31] & x[32]);
  assign t[177] = (x[34] & x[35]);
  assign t[178] = (x[37] & x[38]);
  assign t[179] = (x[40] & x[41]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = (x[43] & x[44]);
  assign t[181] = (x[46] & x[47]);
  assign t[182] = (x[49] & x[50]);
  assign t[183] = (x[54] & x[55]);
  assign t[184] = (x[67] & x[68]);
  assign t[185] = (x[70] & x[71]);
  assign t[186] = (x[75] & x[76]);
  assign t[187] = (x[78] & x[79]);
  assign t[188] = (x[81] & x[82]);
  assign t[189] = (x[84] & x[85]);
  assign t[18] = t[32] ^ t[3];
  assign t[190] = (x[89] & x[90]);
  assign t[191] = (x[92] & x[93]);
  assign t[192] = (x[95] & x[96]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = ~(t[4]);
  assign t[20] = t[35] ^ t[36];
  assign t[21] = t[37] & t[38];
  assign t[22] = t[142] ^ t[39];
  assign t[23] = t[40] ^ t[41];
  assign t[24] = t[42];
  assign t[25] = t[43] ^ t[44];
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[143]);
  assign t[29] = ~(t[144]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[145]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = t[7] ? t[50] : t[146];
  assign t[33] = t[51] ^ t[52];
  assign t[34] = t[53] & t[54];
  assign t[35] = t[55] ? t[56] : t[147];
  assign t[36] = t[55] ? t[57] : t[148];
  assign t[37] = ~(t[58]);
  assign t[38] = t[55] ? t[59] : t[149];
  assign t[39] = t[55] ? t[60] : t[150];
  assign t[3] = t[7] ? t[8] : t[141];
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] & t[64];
  assign t[42] = t[55] ? t[65] : t[151];
  assign t[43] = t[66] ^ t[67];
  assign t[44] = t[68] & t[69];
  assign t[45] = ~(t[70] & t[71]);
  assign t[46] = t[152] | t[72];
  assign t[47] = ~(t[73]);
  assign t[48] = ~(t[142]);
  assign t[49] = ~(t[74] & t[153]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[146] ^ t[75];
  assign t[51] = t[76] & t[77];
  assign t[52] = t[78] & t[79];
  assign t[53] = ~(t[51] ^ t[80]);
  assign t[54] = t[81] ^ t[82];
  assign t[55] = ~(t[14]);
  assign t[56] = t[147] ^ t[83];
  assign t[57] = t[148] ^ t[84];
  assign t[58] = t[55] ? t[85] : t[154];
  assign t[59] = t[149] ^ t[86];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[150] ^ t[87];
  assign t[61] = t[88] & t[89];
  assign t[62] = t[90] & t[91];
  assign t[63] = ~(t[92] ^ t[40]);
  assign t[64] = t[93] ^ t[91];
  assign t[65] = t[151] ^ t[94];
  assign t[66] = t[95] & t[96];
  assign t[67] = t[97] & t[98];
  assign t[68] = ~(t[99] ^ t[43]);
  assign t[69] = t[100] ^ t[98];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[72] & t[101]);
  assign t[71] = ~(t[155] ^ t[102]);
  assign t[72] = ~(t[103] & t[104]);
  assign t[73] = ~(t[46]);
  assign t[74] = ~(t[156]);
  assign t[75] = t[27] ? x[53] : x[52];
  assign t[76] = ~(t[82]);
  assign t[77] = ~(t[105]);
  assign t[78] = ~(t[32]);
  assign t[79] = t[7] ? t[106] : t[157];
  assign t[7] = ~(t[14]);
  assign t[80] = t[18] ^ t[105];
  assign t[81] = t[105] ^ t[3];
  assign t[82] = t[79] ^ t[32];
  assign t[83] = t[107] ? x[58] : x[57];
  assign t[84] = t[73] ? x[60] : x[59];
  assign t[85] = t[154] ^ t[108];
  assign t[86] = t[107] ? x[62] : x[61];
  assign t[87] = t[109] ? x[64] : x[63];
  assign t[88] = ~(t[110]);
  assign t[89] = ~(t[111]);
  assign t[8] = t[141] ^ t[15];
  assign t[90] = ~(t[112]);
  assign t[91] = t[156] ^ t[113];
  assign t[92] = t[111] ^ t[112];
  assign t[93] = t[112] ^ t[22];
  assign t[94] = t[73] ? x[66] : x[65];
  assign t[95] = ~(t[114]);
  assign t[96] = ~(t[115]);
  assign t[97] = ~(t[116]);
  assign t[98] = t[117];
  assign t[99] = t[115] ^ t[116];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind122(x, y);
 input [111:0] x;
 output y;

 wire [202:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[121] ? x[65] : x[64];
  assign t[101] = t[121] ? x[67] : x[66];
  assign t[102] = ~(t[108]);
  assign t[103] = ~(t[128]);
  assign t[104] = ~(t[50]);
  assign t[105] = t[61] ? t[129] : t[169];
  assign t[106] = t[32] ^ t[128];
  assign t[107] = t[128] ^ t[51];
  assign t[108] = t[105] ^ t[50];
  assign t[109] = ~(t[130]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = ~(t[131]);
  assign t[111] = ~(t[132]);
  assign t[112] = t[26] ? t[133] : t[170];
  assign t[113] = t[131] ^ t[132];
  assign t[114] = t[132] ^ t[34];
  assign t[115] = t[27] ? x[75] : x[74];
  assign t[116] = ~(t[134]);
  assign t[117] = ~(t[3]);
  assign t[118] = ~(t[36]);
  assign t[119] = t[7] ? t[135] : t[171];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[166] ^ t[136];
  assign t[121] = ~(t[47]);
  assign t[122] = t[61] ? t[137] : t[172];
  assign t[123] = t[167] ^ t[138];
  assign t[124] = ~(t[127] | t[126]);
  assign t[125] = ~(t[139] | t[98]);
  assign t[126] = ~(t[173]);
  assign t[127] = ~(t[168]);
  assign t[128] = t[61] ? t[140] : t[174];
  assign t[129] = t[169] ^ t[141];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[112] ^ t[132];
  assign t[131] = t[26] ? t[142] : t[175];
  assign t[132] = t[26] ? t[143] : t[176];
  assign t[133] = t[170] ^ t[144];
  assign t[134] = t[60] ^ t[36];
  assign t[135] = t[171] ^ t[145];
  assign t[136] = t[27] ? x[95] : x[94];
  assign t[137] = t[172] ^ t[146];
  assign t[138] = t[121] ? x[97] : x[96];
  assign t[139] = ~(t[158]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[174] ^ t[147];
  assign t[141] = t[121] ? x[99] : x[98];
  assign t[142] = t[175] ^ t[148];
  assign t[143] = t[176] ^ t[149];
  assign t[144] = t[74] ? x[101] : x[100];
  assign t[145] = t[27] ? x[103] : x[102];
  assign t[146] = t[121] ? x[105] : x[104];
  assign t[147] = t[121] ? x[107] : x[106];
  assign t[148] = t[150] ? x[109] : x[108];
  assign t[149] = t[150] ? x[111] : x[110];
  assign t[14] = ~(t[26]);
  assign t[150] = ~(t[47]);
  assign t[151] = t[177] ^ x[4];
  assign t[152] = t[178] ^ x[9];
  assign t[153] = t[179] ^ x[12];
  assign t[154] = t[180] ^ x[15];
  assign t[155] = t[181] ^ x[18];
  assign t[156] = t[182] ^ x[21];
  assign t[157] = t[183] ^ x[24];
  assign t[158] = t[184] ^ x[27];
  assign t[159] = t[185] ^ x[30];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[186] ^ x[33];
  assign t[161] = t[187] ^ x[36];
  assign t[162] = t[188] ^ x[39];
  assign t[163] = t[189] ^ x[42];
  assign t[164] = t[190] ^ x[45];
  assign t[165] = t[191] ^ x[48];
  assign t[166] = t[192] ^ x[53];
  assign t[167] = t[193] ^ x[60];
  assign t[168] = t[194] ^ x[63];
  assign t[169] = t[195] ^ x[70];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[196] ^ x[73];
  assign t[171] = t[197] ^ x[78];
  assign t[172] = t[198] ^ x[81];
  assign t[173] = t[199] ^ x[84];
  assign t[174] = t[200] ^ x[87];
  assign t[175] = t[201] ^ x[90];
  assign t[176] = t[202] ^ x[93];
  assign t[177] = (x[2] & x[3]);
  assign t[178] = (x[7] & x[8]);
  assign t[179] = (x[10] & x[11]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = (x[13] & x[14]);
  assign t[181] = (x[16] & x[17]);
  assign t[182] = (x[19] & x[20]);
  assign t[183] = (x[22] & x[23]);
  assign t[184] = (x[25] & x[26]);
  assign t[185] = (x[28] & x[29]);
  assign t[186] = (x[31] & x[32]);
  assign t[187] = (x[34] & x[35]);
  assign t[188] = (x[37] & x[38]);
  assign t[189] = (x[40] & x[41]);
  assign t[18] = t[32] ^ t[33];
  assign t[190] = (x[43] & x[44]);
  assign t[191] = (x[46] & x[47]);
  assign t[192] = (x[51] & x[52]);
  assign t[193] = (x[58] & x[59]);
  assign t[194] = (x[61] & x[62]);
  assign t[195] = (x[68] & x[69]);
  assign t[196] = (x[71] & x[72]);
  assign t[197] = (x[76] & x[77]);
  assign t[198] = (x[79] & x[80]);
  assign t[199] = (x[82] & x[83]);
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[85] & x[86]);
  assign t[201] = (x[88] & x[89]);
  assign t[202] = (x[91] & x[92]);
  assign t[20] = t[3] ^ t[36];
  assign t[21] = t[37] & t[38];
  assign t[22] = ~t[39];
  assign t[23] = ~t[40];
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[43] & t[44];
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47]);
  assign t[28] = ~(t[152]);
  assign t[29] = ~(t[153]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[154]);
  assign t[31] = ~(t[48] | t[49]);
  assign t[32] = t[50] ^ t[51];
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[26] ? t[54] : t[155];
  assign t[35] = t[55] ^ t[56];
  assign t[36] = t[152] ^ t[57];
  assign t[37] = ~(t[20] ^ t[58]);
  assign t[38] = t[59] ^ t[60];
  assign t[39] = t[61] ? t[62] : t[156];
  assign t[3] = t[7] ? t[8] : t[151];
  assign t[40] = t[61] ? t[63] : t[157];
  assign t[41] = t[64] & t[65];
  assign t[42] = t[66] & t[67];
  assign t[43] = ~(t[41] ^ t[68]);
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[71] & t[72]);
  assign t[46] = t[158] | t[73];
  assign t[47] = ~(t[74]);
  assign t[48] = ~(t[159]);
  assign t[49] = ~(t[75] & t[160]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[61] ? t[76] : t[161];
  assign t[51] = t[61] ? t[77] : t[162];
  assign t[52] = t[78] ^ t[79];
  assign t[53] = t[80] & t[81];
  assign t[54] = t[155] ^ t[82];
  assign t[55] = t[83] ^ t[84];
  assign t[56] = t[85] & t[86];
  assign t[57] = t[7] ? t[87] : t[163];
  assign t[58] = t[88] ^ t[89];
  assign t[59] = t[36] ^ t[90];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[153] ^ t[91];
  assign t[61] = ~(t[14]);
  assign t[62] = t[156] ^ t[92];
  assign t[63] = t[157] ^ t[93];
  assign t[64] = ~(t[70]);
  assign t[65] = ~(t[94]);
  assign t[66] = ~(t[22]);
  assign t[67] = t[95];
  assign t[68] = t[12] ^ t[94];
  assign t[69] = t[94] ^ t[23];
  assign t[6] = t[12] ^ t[13];
  assign t[70] = t[67] ^ t[22];
  assign t[71] = ~(t[73] & t[96]);
  assign t[72] = ~(t[164] ^ t[97]);
  assign t[73] = ~(t[98] & t[99]);
  assign t[74] = ~(t[46]);
  assign t[75] = ~(t[165]);
  assign t[76] = t[161] ^ t[100];
  assign t[77] = t[162] ^ t[101];
  assign t[78] = t[102] & t[103];
  assign t[79] = t[104] & t[105];
  assign t[7] = ~(t[14]);
  assign t[80] = ~(t[78] ^ t[106]);
  assign t[81] = t[107] ^ t[108];
  assign t[82] = t[74] ? x[50] : x[49];
  assign t[83] = t[109] & t[110];
  assign t[84] = t[111] & t[112];
  assign t[85] = ~(t[113] ^ t[55]);
  assign t[86] = t[114] ^ t[112];
  assign t[87] = t[163] ^ t[115];
  assign t[88] = t[116] & t[117];
  assign t[89] = t[118] & t[60];
  assign t[8] = t[151] ^ t[15];
  assign t[90] = t[160] ^ t[119];
  assign t[91] = t[7] ? t[120] : t[166];
  assign t[92] = t[121] ? x[55] : x[54];
  assign t[93] = t[121] ? x[57] : x[56];
  assign t[94] = t[122];
  assign t[95] = t[26] ? t[123] : t[167];
  assign t[96] = ~(t[124] & t[125]);
  assign t[97] = t[126] ^ t[168];
  assign t[98] = ~(t[164]);
  assign t[99] = t[127] & t[126];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind123(x, y);
 input [111:0] x;
 output y;

 wire [203:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = ~(t[128] & t[129]);
  assign t[101] = t[130] ^ t[172];
  assign t[102] = ~(t[167]);
  assign t[103] = t[131] & t[130];
  assign t[104] = t[169] ^ t[132];
  assign t[105] = t[133] ? x[72] : x[71];
  assign t[106] = t[133] ? x[74] : x[73];
  assign t[107] = ~(t[134]);
  assign t[108] = ~(t[35]);
  assign t[109] = ~(t[36]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[77] ? t[135] : t[173];
  assign t[111] = t[170] ^ t[136];
  assign t[112] = t[137] ? x[79] : x[78];
  assign t[113] = t[73] ? x[81] : x[80];
  assign t[114] = ~(t[120]);
  assign t[115] = ~(t[138]);
  assign t[116] = ~(t[58]);
  assign t[117] = t[26] ? t[139] : t[174];
  assign t[118] = t[39] ^ t[138];
  assign t[119] = t[138] ^ t[59];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[117] ^ t[58];
  assign t[121] = t[133] ? x[86] : x[85];
  assign t[122] = t[133] ? x[88] : x[87];
  assign t[123] = t[140] & t[141];
  assign t[124] = t[142] & t[94];
  assign t[125] = t[77] ? t[143] : t[175];
  assign t[126] = t[171] ^ t[144];
  assign t[127] = t[34] ^ t[52];
  assign t[128] = ~(t[131] | t[130]);
  assign t[129] = ~(t[145] | t[102]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = ~(t[176]);
  assign t[131] = ~(t[172]);
  assign t[132] = t[27] ? x[96] : x[95];
  assign t[133] = ~(t[48]);
  assign t[134] = t[57] ^ t[36];
  assign t[135] = t[173] ^ t[146];
  assign t[136] = t[133] ? x[98] : x[97];
  assign t[137] = ~(t[48]);
  assign t[138] = t[26] ? t[147] : t[177];
  assign t[139] = t[174] ^ t[148];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[149]);
  assign t[141] = ~(t[62]);
  assign t[142] = ~(t[63]);
  assign t[143] = t[175] ^ t[150];
  assign t[144] = t[133] ? x[103] : x[102];
  assign t[145] = ~(t[159]);
  assign t[146] = t[133] ? x[105] : x[104];
  assign t[147] = t[177] ^ t[151];
  assign t[148] = t[73] ? x[107] : x[106];
  assign t[149] = t[94] ^ t[63];
  assign t[14] = ~(t[26]);
  assign t[150] = t[133] ? x[109] : x[108];
  assign t[151] = t[137] ? x[111] : x[110];
  assign t[152] = t[178] ^ x[4];
  assign t[153] = t[179] ^ x[9];
  assign t[154] = t[180] ^ x[12];
  assign t[155] = t[181] ^ x[15];
  assign t[156] = t[182] ^ x[18];
  assign t[157] = t[183] ^ x[21];
  assign t[158] = t[184] ^ x[24];
  assign t[159] = t[185] ^ x[27];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[186] ^ x[30];
  assign t[161] = t[187] ^ x[33];
  assign t[162] = t[188] ^ x[36];
  assign t[163] = t[189] ^ x[39];
  assign t[164] = t[190] ^ x[42];
  assign t[165] = t[191] ^ x[45];
  assign t[166] = t[192] ^ x[48];
  assign t[167] = t[193] ^ x[51];
  assign t[168] = t[194] ^ x[54];
  assign t[169] = t[195] ^ x[59];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[196] ^ x[62];
  assign t[171] = t[197] ^ x[65];
  assign t[172] = t[198] ^ x[70];
  assign t[173] = t[199] ^ x[77];
  assign t[174] = t[200] ^ x[84];
  assign t[175] = t[201] ^ x[91];
  assign t[176] = t[202] ^ x[94];
  assign t[177] = t[203] ^ x[101];
  assign t[178] = (x[2] & x[3]);
  assign t[179] = (x[7] & x[8]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = (x[10] & x[11]);
  assign t[181] = (x[13] & x[14]);
  assign t[182] = (x[16] & x[17]);
  assign t[183] = (x[19] & x[20]);
  assign t[184] = (x[22] & x[23]);
  assign t[185] = (x[25] & x[26]);
  assign t[186] = (x[28] & x[29]);
  assign t[187] = (x[31] & x[32]);
  assign t[188] = (x[34] & x[35]);
  assign t[189] = (x[37] & x[38]);
  assign t[18] = t[32] ^ t[24];
  assign t[190] = (x[40] & x[41]);
  assign t[191] = (x[43] & x[44]);
  assign t[192] = (x[46] & x[47]);
  assign t[193] = (x[49] & x[50]);
  assign t[194] = (x[52] & x[53]);
  assign t[195] = (x[57] & x[58]);
  assign t[196] = (x[60] & x[61]);
  assign t[197] = (x[63] & x[64]);
  assign t[198] = (x[68] & x[69]);
  assign t[199] = (x[75] & x[76]);
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[82] & x[83]);
  assign t[201] = (x[89] & x[90]);
  assign t[202] = (x[92] & x[93]);
  assign t[203] = (x[99] & x[100]);
  assign t[20] = t[35] ^ t[36];
  assign t[21] = t[37] & t[38];
  assign t[22] = t[39] ^ t[40];
  assign t[23] = t[41] ^ t[42];
  assign t[24] = t[153] ^ t[43];
  assign t[25] = t[44] ^ t[45];
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48]);
  assign t[28] = ~(t[154]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[156]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = t[7] ? t[51] : t[157];
  assign t[33] = ~(t[52]);
  assign t[34] = t[155] ^ t[3];
  assign t[35] = t[53];
  assign t[36] = ~t[54];
  assign t[37] = ~(t[20] ^ t[55]);
  assign t[38] = t[56] ^ t[57];
  assign t[39] = t[58] ^ t[59];
  assign t[3] = t[7] ? t[8] : t[152];
  assign t[40] = t[60] ^ t[61];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] & t[65];
  assign t[43] = t[7] ? t[66] : t[158];
  assign t[44] = t[67] ^ t[19];
  assign t[45] = t[68] & t[69];
  assign t[46] = ~(t[70] & t[71]);
  assign t[47] = t[159] | t[72];
  assign t[48] = ~(t[73]);
  assign t[49] = ~(t[160]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[74] & t[153]);
  assign t[51] = t[157] ^ t[75];
  assign t[52] = t[154] ^ t[76];
  assign t[53] = t[77] ? t[78] : t[161];
  assign t[54] = t[77] ? t[79] : t[162];
  assign t[55] = t[80] ^ t[81];
  assign t[56] = t[36] ^ t[82];
  assign t[57] = t[83];
  assign t[58] = t[26] ? t[84] : t[163];
  assign t[59] = t[26] ? t[85] : t[164];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[86] ^ t[87];
  assign t[61] = t[88] & t[89];
  assign t[62] = t[77] ? t[90] : t[165];
  assign t[63] = t[77] ? t[91] : t[166];
  assign t[64] = ~(t[41] ^ t[92]);
  assign t[65] = t[93] ^ t[94];
  assign t[66] = t[158] ^ t[95];
  assign t[67] = t[96] & t[97];
  assign t[68] = ~(t[98] ^ t[44]);
  assign t[69] = t[99] ^ t[34];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[72] & t[100]);
  assign t[71] = ~(t[167] ^ t[101]);
  assign t[72] = ~(t[102] & t[103]);
  assign t[73] = ~(t[47]);
  assign t[74] = ~(t[168]);
  assign t[75] = t[27] ? x[56] : x[55];
  assign t[76] = t[7] ? t[104] : t[169];
  assign t[77] = ~(t[14]);
  assign t[78] = t[161] ^ t[105];
  assign t[79] = t[162] ^ t[106];
  assign t[7] = ~(t[14]);
  assign t[80] = t[107] & t[108];
  assign t[81] = t[109] & t[57];
  assign t[82] = ~t[110];
  assign t[83] = t[26] ? t[111] : t[170];
  assign t[84] = t[163] ^ t[112];
  assign t[85] = t[164] ^ t[113];
  assign t[86] = t[114] & t[115];
  assign t[87] = t[116] & t[117];
  assign t[88] = ~(t[86] ^ t[118]);
  assign t[89] = t[119] ^ t[120];
  assign t[8] = t[152] ^ t[15];
  assign t[90] = t[165] ^ t[121];
  assign t[91] = t[166] ^ t[122];
  assign t[92] = t[123] ^ t[124];
  assign t[93] = t[63] ^ t[125];
  assign t[94] = t[77] ? t[126] : t[171];
  assign t[95] = t[27] ? x[67] : x[66];
  assign t[96] = ~(t[127]);
  assign t[97] = ~(t[32]);
  assign t[98] = t[32] ^ t[52];
  assign t[99] = t[52] ^ t[24];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind124(x, y);
 input [111:0] x;
 output y;

 wire [214:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[40] ^ t[66];
  assign t[101] = t[66] ^ t[24];
  assign t[102] = ~(t[131] & t[132]);
  assign t[103] = t[133] ^ t[182];
  assign t[104] = ~(t[175]);
  assign t[105] = t[134] & t[133];
  assign t[106] = t[97] ? x[71] : x[70];
  assign t[107] = ~(t[135]);
  assign t[108] = ~(t[55]);
  assign t[109] = t[55] ^ t[82];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[82] ^ t[32];
  assign t[111] = t[177] ^ t[136];
  assign t[112] = t[43] ? t[137] : t[183];
  assign t[113] = t[178] ^ t[138];
  assign t[114] = t[179] ^ t[139];
  assign t[115] = t[180] ^ t[140];
  assign t[116] = t[141] ^ t[142];
  assign t[117] = t[85] ^ t[143];
  assign t[118] = t[26] ? t[144] : t[184];
  assign t[119] = t[181] ^ t[145];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = ~(t[146] ^ t[63]);
  assign t[121] = t[38] ^ t[125];
  assign t[122] = ~(t[128]);
  assign t[123] = ~(t[147]);
  assign t[124] = ~(t[62]);
  assign t[125] = t[166] ^ t[148];
  assign t[126] = t[38] ^ t[147];
  assign t[127] = t[147] ^ t[60];
  assign t[128] = t[125] ^ t[62];
  assign t[129] = t[97] ? x[79] : x[78];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[42] ^ t[66];
  assign t[131] = ~(t[134] | t[133]);
  assign t[132] = ~(t[149] | t[104]);
  assign t[133] = ~(t[185]);
  assign t[134] = ~(t[182]);
  assign t[135] = t[57] ^ t[82];
  assign t[136] = t[97] ? x[84] : x[83];
  assign t[137] = t[183] ^ t[150];
  assign t[138] = t[97] ? x[86] : x[85];
  assign t[139] = t[151] ? x[88] : x[87];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[151] ? x[90] : x[89];
  assign t[141] = t[152] & t[153];
  assign t[142] = t[154] & t[118];
  assign t[143] = t[26] ? t[155] : t[186];
  assign t[144] = t[184] ^ t[156];
  assign t[145] = t[27] ? x[95] : x[94];
  assign t[146] = t[147] ^ t[62];
  assign t[147] = t[7] ? t[157] : t[187];
  assign t[148] = t[7] ? t[158] : t[188];
  assign t[149] = ~(t[170]);
  assign t[14] = ~(t[26]);
  assign t[150] = t[97] ? x[103] : x[102];
  assign t[151] = ~(t[49]);
  assign t[152] = ~(t[159]);
  assign t[153] = ~(t[84]);
  assign t[154] = ~(t[85]);
  assign t[155] = t[186] ^ t[160];
  assign t[156] = t[75] ? x[105] : x[104];
  assign t[157] = t[187] ^ t[161];
  assign t[158] = t[188] ^ t[162];
  assign t[159] = t[118] ^ t[85];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[75] ? x[107] : x[106];
  assign t[161] = t[27] ? x[109] : x[108];
  assign t[162] = t[27] ? x[111] : x[110];
  assign t[163] = t[189] ^ x[4];
  assign t[164] = t[190] ^ x[9];
  assign t[165] = t[191] ^ x[12];
  assign t[166] = t[192] ^ x[15];
  assign t[167] = t[193] ^ x[18];
  assign t[168] = t[194] ^ x[21];
  assign t[169] = t[195] ^ x[24];
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = t[196] ^ x[27];
  assign t[171] = t[197] ^ x[30];
  assign t[172] = t[198] ^ x[33];
  assign t[173] = t[199] ^ x[36];
  assign t[174] = t[200] ^ x[39];
  assign t[175] = t[201] ^ x[44];
  assign t[176] = t[202] ^ x[47];
  assign t[177] = t[203] ^ x[50];
  assign t[178] = t[204] ^ x[53];
  assign t[179] = t[205] ^ x[56];
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = t[206] ^ x[59];
  assign t[181] = t[207] ^ x[62];
  assign t[182] = t[208] ^ x[69];
  assign t[183] = t[209] ^ x[74];
  assign t[184] = t[210] ^ x[77];
  assign t[185] = t[211] ^ x[82];
  assign t[186] = t[212] ^ x[93];
  assign t[187] = t[213] ^ x[98];
  assign t[188] = t[214] ^ x[101];
  assign t[189] = (x[2] & x[3]);
  assign t[18] = t[32] ^ t[33];
  assign t[190] = (x[7] & x[8]);
  assign t[191] = (x[10] & x[11]);
  assign t[192] = (x[13] & x[14]);
  assign t[193] = (x[16] & x[17]);
  assign t[194] = (x[19] & x[20]);
  assign t[195] = (x[22] & x[23]);
  assign t[196] = (x[25] & x[26]);
  assign t[197] = (x[28] & x[29]);
  assign t[198] = (x[31] & x[32]);
  assign t[199] = (x[34] & x[35]);
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[37] & x[38]);
  assign t[201] = (x[42] & x[43]);
  assign t[202] = (x[45] & x[46]);
  assign t[203] = (x[48] & x[49]);
  assign t[204] = (x[51] & x[52]);
  assign t[205] = (x[54] & x[55]);
  assign t[206] = (x[57] & x[58]);
  assign t[207] = (x[60] & x[61]);
  assign t[208] = (x[67] & x[68]);
  assign t[209] = (x[72] & x[73]);
  assign t[20] = ~(t[36] ^ t[37]);
  assign t[210] = (x[75] & x[76]);
  assign t[211] = (x[80] & x[81]);
  assign t[212] = (x[91] & x[92]);
  assign t[213] = (x[96] & x[97]);
  assign t[214] = (x[99] & x[100]);
  assign t[21] = t[38] ^ t[39];
  assign t[22] = t[40] ^ t[24];
  assign t[23] = t[41] & t[42];
  assign t[24] = t[43] ? t[44] : t[164];
  assign t[25] = t[45] ^ t[46];
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49]);
  assign t[28] = ~(t[165]);
  assign t[29] = ~(t[166]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[167]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~t[52];
  assign t[33] = t[53] ^ t[54];
  assign t[34] = t[55] ^ t[32];
  assign t[35] = t[56] & t[57];
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[62] ^ t[60];
  assign t[39] = t[63] ^ t[64];
  assign t[3] = t[7] ? t[8] : t[163];
  assign t[40] = t[43] ? t[65] : t[168];
  assign t[41] = ~(t[66]);
  assign t[42] = t[43] ? t[67] : t[169];
  assign t[43] = ~(t[14]);
  assign t[44] = t[164] ^ t[68];
  assign t[45] = t[69] ^ t[23];
  assign t[46] = t[70] & t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[170] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[171]);
  assign t[51] = ~(t[76] & t[172]);
  assign t[52] = t[43] ? t[77] : t[173];
  assign t[53] = t[78] ^ t[35];
  assign t[54] = t[79] & t[80];
  assign t[55] = t[81];
  assign t[56] = ~(t[82]);
  assign t[57] = t[83];
  assign t[58] = t[84] ^ t[85];
  assign t[59] = t[86] & t[87];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[172] ^ t[88];
  assign t[61] = t[63] ^ t[89];
  assign t[62] = t[165] ^ t[3];
  assign t[63] = t[90] ^ t[91];
  assign t[64] = t[92] & t[93];
  assign t[65] = t[168] ^ t[94];
  assign t[66] = t[43] ? t[95] : t[174];
  assign t[67] = t[169] ^ t[96];
  assign t[68] = t[97] ? x[41] : x[40];
  assign t[69] = t[98] & t[99];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[100] ^ t[45]);
  assign t[71] = t[101] ^ t[42];
  assign t[72] = ~(t[74] & t[102]);
  assign t[73] = ~(t[175] ^ t[103]);
  assign t[74] = ~(t[104] & t[105]);
  assign t[75] = ~(t[48]);
  assign t[76] = ~(t[176]);
  assign t[77] = t[173] ^ t[106];
  assign t[78] = t[107] & t[108];
  assign t[79] = ~(t[109] ^ t[53]);
  assign t[7] = ~(t[14]);
  assign t[80] = t[110] ^ t[57];
  assign t[81] = t[43] ? t[111] : t[177];
  assign t[82] = ~t[112];
  assign t[83] = t[26] ? t[113] : t[178];
  assign t[84] = t[26] ? t[114] : t[179];
  assign t[85] = t[26] ? t[115] : t[180];
  assign t[86] = ~(t[58] ^ t[116]);
  assign t[87] = t[117] ^ t[118];
  assign t[88] = t[7] ? t[119] : t[181];
  assign t[89] = t[120] & t[121];
  assign t[8] = t[163] ^ t[15];
  assign t[90] = t[122] & t[123];
  assign t[91] = t[124] & t[125];
  assign t[92] = ~(t[90] ^ t[126]);
  assign t[93] = t[127] ^ t[128];
  assign t[94] = t[97] ? x[64] : x[63];
  assign t[95] = t[174] ^ t[129];
  assign t[96] = t[97] ? x[66] : x[65];
  assign t[97] = ~(t[49]);
  assign t[98] = ~(t[130]);
  assign t[99] = ~(t[40]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind125(x, y);
 input [111:0] x;
 output y;

 wire [192:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[116] ^ t[117];
  assign t[101] = t[117] ^ t[24];
  assign t[102] = ~(t[119] & t[120]);
  assign t[103] = t[121] ^ t[158];
  assign t[104] = ~(t[155]);
  assign t[105] = t[122] & t[121];
  assign t[106] = t[27] ? x[69] : x[68];
  assign t[107] = t[7] ? t[123] : t[159];
  assign t[108] = t[7] ? t[124] : t[160];
  assign t[109] = ~(t[49]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[109] ? x[77] : x[76];
  assign t[111] = t[92] ^ t[113];
  assign t[112] = t[125];
  assign t[113] = ~t[126];
  assign t[114] = t[26] ? t[127] : t[161];
  assign t[115] = t[99] ^ t[117];
  assign t[116] = t[43] ? t[128] : t[162];
  assign t[117] = t[43] ? t[129] : t[163];
  assign t[118] = t[157] ^ t[130];
  assign t[119] = ~(t[122] | t[121]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = ~(t[131] | t[104]);
  assign t[121] = ~(t[164]);
  assign t[122] = ~(t[158]);
  assign t[123] = t[159] ^ t[132];
  assign t[124] = t[160] ^ t[133];
  assign t[125] = t[43] ? t[134] : t[165];
  assign t[126] = t[43] ? t[135] : t[166];
  assign t[127] = t[161] ^ t[136];
  assign t[128] = t[162] ^ t[137];
  assign t[129] = t[163] ^ t[138];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[95] ? x[97] : x[96];
  assign t[131] = ~(t[151]);
  assign t[132] = t[27] ? x[99] : x[98];
  assign t[133] = t[27] ? x[101] : x[100];
  assign t[134] = t[165] ^ t[139];
  assign t[135] = t[166] ^ t[140];
  assign t[136] = t[95] ? x[103] : x[102];
  assign t[137] = t[95] ? x[105] : x[104];
  assign t[138] = t[95] ? x[107] : x[106];
  assign t[139] = t[95] ? x[109] : x[108];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[95] ? x[111] : x[110];
  assign t[141] = t[167] ^ x[4];
  assign t[142] = t[168] ^ x[9];
  assign t[143] = t[169] ^ x[12];
  assign t[144] = t[170] ^ x[15];
  assign t[145] = t[171] ^ x[18];
  assign t[146] = t[172] ^ x[21];
  assign t[147] = t[173] ^ x[24];
  assign t[148] = t[174] ^ x[27];
  assign t[149] = t[175] ^ x[30];
  assign t[14] = ~(t[26]);
  assign t[150] = t[176] ^ x[33];
  assign t[151] = t[177] ^ x[36];
  assign t[152] = t[178] ^ x[39];
  assign t[153] = t[179] ^ x[42];
  assign t[154] = t[180] ^ x[45];
  assign t[155] = t[181] ^ x[50];
  assign t[156] = t[182] ^ x[53];
  assign t[157] = t[183] ^ x[64];
  assign t[158] = t[184] ^ x[67];
  assign t[159] = t[185] ^ x[72];
  assign t[15] = t[27] ? x[6] : x[5];
  assign t[160] = t[186] ^ x[75];
  assign t[161] = t[187] ^ x[80];
  assign t[162] = t[188] ^ x[83];
  assign t[163] = t[189] ^ x[86];
  assign t[164] = t[190] ^ x[89];
  assign t[165] = t[191] ^ x[92];
  assign t[166] = t[192] ^ x[95];
  assign t[167] = (x[2] & x[3]);
  assign t[168] = (x[7] & x[8]);
  assign t[169] = (x[10] & x[11]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[170] = (x[13] & x[14]);
  assign t[171] = (x[16] & x[17]);
  assign t[172] = (x[19] & x[20]);
  assign t[173] = (x[22] & x[23]);
  assign t[174] = (x[25] & x[26]);
  assign t[175] = (x[28] & x[29]);
  assign t[176] = (x[31] & x[32]);
  assign t[177] = (x[34] & x[35]);
  assign t[178] = (x[37] & x[38]);
  assign t[179] = (x[40] & x[41]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[180] = (x[43] & x[44]);
  assign t[181] = (x[48] & x[49]);
  assign t[182] = (x[51] & x[52]);
  assign t[183] = (x[62] & x[63]);
  assign t[184] = (x[65] & x[66]);
  assign t[185] = (x[70] & x[71]);
  assign t[186] = (x[73] & x[74]);
  assign t[187] = (x[78] & x[79]);
  assign t[188] = (x[81] & x[82]);
  assign t[189] = (x[84] & x[85]);
  assign t[18] = t[32] ^ t[33];
  assign t[190] = (x[87] & x[88]);
  assign t[191] = (x[90] & x[91]);
  assign t[192] = (x[93] & x[94]);
  assign t[19] = t[34] ^ t[35];
  assign t[1] = ~(t[4]);
  assign t[20] = t[36] ^ t[37];
  assign t[21] = t[38] & t[39];
  assign t[22] = ~t[40];
  assign t[23] = t[41] ^ t[42];
  assign t[24] = t[43] ? t[44] : t[142];
  assign t[25] = t[45] ^ t[46];
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49]);
  assign t[28] = ~(t[143]);
  assign t[29] = ~(t[144]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[145]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = t[143] ^ t[52];
  assign t[33] = t[146] ^ t[3];
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[55] & t[56];
  assign t[36] = t[26] ? t[57] : t[147];
  assign t[37] = t[26] ? t[58] : t[148];
  assign t[38] = ~(t[59]);
  assign t[39] = t[26] ? t[60] : t[149];
  assign t[3] = t[7] ? t[8] : t[141];
  assign t[40] = t[43] ? t[61] : t[150];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] & t[65];
  assign t[43] = ~(t[14]);
  assign t[44] = t[142] ^ t[66];
  assign t[45] = t[67] ^ t[68];
  assign t[46] = t[69] & t[70];
  assign t[47] = ~(t[71] & t[72]);
  assign t[48] = t[151] | t[73];
  assign t[49] = ~(t[74]);
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[152]);
  assign t[51] = ~(t[75] & t[146]);
  assign t[52] = t[7] ? t[76] : t[153];
  assign t[53] = t[77] & t[78];
  assign t[54] = t[79] & t[80];
  assign t[55] = ~(t[53] ^ t[81]);
  assign t[56] = t[82] ^ t[83];
  assign t[57] = t[147] ^ t[84];
  assign t[58] = t[148] ^ t[85];
  assign t[59] = t[26] ? t[86] : t[154];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[149] ^ t[87];
  assign t[61] = t[150] ^ t[88];
  assign t[62] = t[89] & t[90];
  assign t[63] = t[91] & t[92];
  assign t[64] = ~(t[93] ^ t[41]);
  assign t[65] = t[94] ^ t[92];
  assign t[66] = t[95] ? x[47] : x[46];
  assign t[67] = t[96] & t[97];
  assign t[68] = t[98] & t[99];
  assign t[69] = ~(t[100] ^ t[45]);
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[101] ^ t[99];
  assign t[71] = ~(t[73] & t[102]);
  assign t[72] = ~(t[155] ^ t[103]);
  assign t[73] = ~(t[104] & t[105]);
  assign t[74] = ~(t[48]);
  assign t[75] = ~(t[156]);
  assign t[76] = t[153] ^ t[106];
  assign t[77] = ~(t[83]);
  assign t[78] = ~(t[107]);
  assign t[79] = ~(t[32]);
  assign t[7] = ~(t[14]);
  assign t[80] = t[144] ^ t[108];
  assign t[81] = t[18] ^ t[107];
  assign t[82] = t[107] ^ t[33];
  assign t[83] = t[80] ^ t[32];
  assign t[84] = t[109] ? x[55] : x[54];
  assign t[85] = t[74] ? x[57] : x[56];
  assign t[86] = t[154] ^ t[110];
  assign t[87] = t[74] ? x[59] : x[58];
  assign t[88] = t[95] ? x[61] : x[60];
  assign t[89] = ~(t[111]);
  assign t[8] = t[141] ^ t[15];
  assign t[90] = ~(t[112]);
  assign t[91] = ~(t[113]);
  assign t[92] = t[114];
  assign t[93] = t[112] ^ t[113];
  assign t[94] = t[113] ^ t[22];
  assign t[95] = ~(t[49]);
  assign t[96] = ~(t[115]);
  assign t[97] = ~(t[116]);
  assign t[98] = ~(t[117]);
  assign t[99] = t[43] ? t[118] : t[157];
  assign t[9] = ~(t[16] | t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind126(x, y);
 input [111:0] x;
 output y;

 wire [202:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[43] ? t[126] : t[170];
  assign t[101] = t[166] ^ t[127];
  assign t[102] = ~(t[152]);
  assign t[103] = t[128] ? x[69] : x[68];
  assign t[104] = t[128] ? x[71] : x[70];
  assign t[105] = ~(t[111]);
  assign t[106] = ~(t[129]);
  assign t[107] = ~(t[56]);
  assign t[108] = t[43] ? t[130] : t[171];
  assign t[109] = t[35] ^ t[129];
  assign t[10] = t[19] ^ t[20];
  assign t[110] = t[129] ^ t[57];
  assign t[111] = t[108] ^ t[56];
  assign t[112] = t[131] ? x[76] : x[75];
  assign t[113] = ~(t[132]);
  assign t[114] = ~(t[133]);
  assign t[115] = ~(t[134]);
  assign t[116] = t[168] ^ t[135];
  assign t[117] = t[133] ^ t[134];
  assign t[118] = t[134] ^ t[37];
  assign t[119] = t[131] ? x[78] : x[77];
  assign t[11] = t[21] ^ t[22];
  assign t[120] = ~(t[136]);
  assign t[121] = ~(t[39]);
  assign t[122] = ~(t[40]);
  assign t[123] = t[7] ? t[137] : t[172];
  assign t[124] = t[169] ^ t[138];
  assign t[125] = ~(t[30]);
  assign t[126] = t[170] ^ t[139];
  assign t[127] = t[99] ? x[83] : x[82];
  assign t[128] = ~(t[125]);
  assign t[129] = t[43] ? t[140] : t[173];
  assign t[12] = t[23] ^ t[24];
  assign t[130] = t[171] ^ t[141];
  assign t[131] = ~(t[125]);
  assign t[132] = t[116] ^ t[134];
  assign t[133] = t[7] ? t[142] : t[174];
  assign t[134] = t[158] ^ t[143];
  assign t[135] = t[7] ? t[144] : t[175];
  assign t[136] = t[66] ^ t[40];
  assign t[137] = t[172] ^ t[145];
  assign t[138] = t[131] ? x[94] : x[93];
  assign t[139] = t[99] ? x[96] : x[95];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[173] ^ t[146];
  assign t[141] = t[128] ? x[98] : x[97];
  assign t[142] = t[174] ^ t[147];
  assign t[143] = t[7] ? t[148] : t[176];
  assign t[144] = t[175] ^ t[149];
  assign t[145] = t[30] ? x[103] : x[102];
  assign t[146] = t[128] ? x[105] : x[104];
  assign t[147] = t[99] ? x[107] : x[106];
  assign t[148] = t[176] ^ t[150];
  assign t[149] = t[30] ? x[109] : x[108];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[99] ? x[111] : x[110];
  assign t[151] = t[177] ^ x[4];
  assign t[152] = t[178] ^ x[7];
  assign t[153] = t[179] ^ x[12];
  assign t[154] = t[180] ^ x[15];
  assign t[155] = t[181] ^ x[18];
  assign t[156] = t[182] ^ x[21];
  assign t[157] = t[183] ^ x[24];
  assign t[158] = t[184] ^ x[27];
  assign t[159] = t[185] ^ x[30];
  assign t[15] = t[152] | t[29];
  assign t[160] = t[186] ^ x[33];
  assign t[161] = t[187] ^ x[36];
  assign t[162] = t[188] ^ x[39];
  assign t[163] = t[189] ^ x[42];
  assign t[164] = t[190] ^ x[45];
  assign t[165] = t[191] ^ x[48];
  assign t[166] = t[192] ^ x[55];
  assign t[167] = t[193] ^ x[58];
  assign t[168] = t[194] ^ x[61];
  assign t[169] = t[195] ^ x[64];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[196] ^ x[67];
  assign t[171] = t[197] ^ x[74];
  assign t[172] = t[198] ^ x[81];
  assign t[173] = t[199] ^ x[86];
  assign t[174] = t[200] ^ x[89];
  assign t[175] = t[201] ^ x[92];
  assign t[176] = t[202] ^ x[101];
  assign t[177] = (x[2] & x[3]);
  assign t[178] = (x[5] & x[6]);
  assign t[179] = (x[10] & x[11]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = (x[13] & x[14]);
  assign t[181] = (x[16] & x[17]);
  assign t[182] = (x[19] & x[20]);
  assign t[183] = (x[22] & x[23]);
  assign t[184] = (x[25] & x[26]);
  assign t[185] = (x[28] & x[29]);
  assign t[186] = (x[31] & x[32]);
  assign t[187] = (x[34] & x[35]);
  assign t[188] = (x[37] & x[38]);
  assign t[189] = (x[40] & x[41]);
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = (x[43] & x[44]);
  assign t[191] = (x[46] & x[47]);
  assign t[192] = (x[53] & x[54]);
  assign t[193] = (x[56] & x[57]);
  assign t[194] = (x[59] & x[60]);
  assign t[195] = (x[62] & x[63]);
  assign t[196] = (x[65] & x[66]);
  assign t[197] = (x[72] & x[73]);
  assign t[198] = (x[79] & x[80]);
  assign t[199] = (x[84] & x[85]);
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[87] & x[88]);
  assign t[201] = (x[90] & x[91]);
  assign t[202] = (x[99] & x[100]);
  assign t[20] = t[37] ^ t[38];
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[41] & t[42];
  assign t[23] = t[43] ? t[44] : t[153];
  assign t[24] = t[43] ? t[45] : t[154];
  assign t[25] = t[46] ^ t[47];
  assign t[26] = t[48] & t[49];
  assign t[27] = ~(t[29] & t[50]);
  assign t[28] = ~(t[155] ^ t[51]);
  assign t[29] = ~(t[52] & t[53]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[15]);
  assign t[31] = ~(t[156]);
  assign t[32] = ~(t[157]);
  assign t[33] = ~(t[158]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = t[56] ^ t[57];
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[159] ^ t[60];
  assign t[38] = t[61] ^ t[62];
  assign t[39] = ~t[3];
  assign t[3] = t[7] ? t[8] : t[151];
  assign t[40] = t[63];
  assign t[41] = ~(t[21] ^ t[64]);
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[67]);
  assign t[44] = t[153] ^ t[68];
  assign t[45] = t[154] ^ t[69];
  assign t[46] = t[70] & t[71];
  assign t[47] = t[72] & t[73];
  assign t[48] = ~(t[46] ^ t[74]);
  assign t[49] = t[75] ^ t[76];
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[77] & t[78]);
  assign t[51] = t[79] ^ t[160];
  assign t[52] = ~(t[155]);
  assign t[53] = t[80] & t[79];
  assign t[54] = ~(t[159]);
  assign t[55] = ~(t[81] & t[161]);
  assign t[56] = t[43] ? t[82] : t[162];
  assign t[57] = t[43] ? t[83] : t[163];
  assign t[58] = t[84] ^ t[85];
  assign t[59] = t[86] & t[87];
  assign t[5] = ~(t[10] ^ t[11]);
  assign t[60] = t[88] ? t[89] : t[164];
  assign t[61] = t[90] ^ t[91];
  assign t[62] = t[92] & t[93];
  assign t[63] = t[7] ? t[94] : t[165];
  assign t[64] = t[95] ^ t[96];
  assign t[65] = t[40] ^ t[97];
  assign t[66] = t[98];
  assign t[67] = ~(t[7]);
  assign t[68] = t[99] ? x[50] : x[49];
  assign t[69] = t[99] ? x[52] : x[51];
  assign t[6] = t[12] ^ t[13];
  assign t[70] = ~(t[76]);
  assign t[71] = ~(t[100]);
  assign t[72] = ~(t[23]);
  assign t[73] = t[43] ? t[101] : t[166];
  assign t[74] = t[12] ^ t[100];
  assign t[75] = t[100] ^ t[24];
  assign t[76] = t[73] ^ t[23];
  assign t[77] = ~(t[80] | t[79]);
  assign t[78] = ~(t[102] | t[52]);
  assign t[79] = ~(t[167]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[160]);
  assign t[81] = ~(t[168]);
  assign t[82] = t[162] ^ t[103];
  assign t[83] = t[163] ^ t[104];
  assign t[84] = t[105] & t[106];
  assign t[85] = t[107] & t[108];
  assign t[86] = ~(t[84] ^ t[109]);
  assign t[87] = t[110] ^ t[111];
  assign t[88] = ~(t[67]);
  assign t[89] = t[164] ^ t[112];
  assign t[8] = t[151] ^ t[16];
  assign t[90] = t[113] & t[114];
  assign t[91] = t[115] & t[116];
  assign t[92] = ~(t[117] ^ t[61]);
  assign t[93] = t[118] ^ t[116];
  assign t[94] = t[165] ^ t[119];
  assign t[95] = t[120] & t[121];
  assign t[96] = t[122] & t[66];
  assign t[97] = t[123];
  assign t[98] = t[7] ? t[124] : t[169];
  assign t[99] = ~(t[125]);
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind127(x, y);
 input [111:0] x;
 output y;

 wire [203:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[69] ^ t[130];
  assign t[101] = t[58] ? t[131] : t[174];
  assign t[102] = t[80] ? x[78] : x[77];
  assign t[103] = ~(t[132]);
  assign t[104] = ~(t[35]);
  assign t[105] = t[35] ^ t[57];
  assign t[106] = t[57] ^ t[25];
  assign t[107] = ~(t[153]);
  assign t[108] = t[80] ? x[80] : x[79];
  assign t[109] = t[170] ^ t[133];
  assign t[10] = t[19] ^ t[20];
  assign t[110] = ~(t[53]);
  assign t[111] = ~(t[134]);
  assign t[112] = ~(t[38]);
  assign t[113] = ~(t[39]);
  assign t[114] = t[171] ^ t[135];
  assign t[115] = t[110] ? x[82] : x[81];
  assign t[116] = t[172] ^ t[136];
  assign t[117] = ~(t[84]);
  assign t[118] = t[173] ^ t[137];
  assign t[119] = ~(t[125]);
  assign t[11] = t[21] ^ t[22];
  assign t[120] = ~(t[138]);
  assign t[121] = ~(t[64]);
  assign t[122] = t[169] ^ t[139];
  assign t[123] = t[42] ^ t[138];
  assign t[124] = t[138] ^ t[65];
  assign t[125] = t[122] ^ t[64];
  assign t[126] = t[140] ? x[84] : x[83];
  assign t[127] = t[140] ? x[86] : x[85];
  assign t[128] = t[141] & t[142];
  assign t[129] = t[143] & t[101];
  assign t[12] = t[23] ^ t[24];
  assign t[130] = t[58] ? t[144] : t[175];
  assign t[131] = t[174] ^ t[145];
  assign t[132] = t[37] ^ t[57];
  assign t[133] = t[30] ? x[91] : x[90];
  assign t[134] = t[63] ^ t[39];
  assign t[135] = t[110] ? x[93] : x[92];
  assign t[136] = t[110] ? x[95] : x[94];
  assign t[137] = t[30] ? x[97] : x[96];
  assign t[138] = t[7] ? t[146] : t[176];
  assign t[139] = t[7] ? t[147] : t[177];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = ~(t[53]);
  assign t[141] = ~(t[148]);
  assign t[142] = ~(t[68]);
  assign t[143] = ~(t[69]);
  assign t[144] = t[175] ^ t[149];
  assign t[145] = t[140] ? x[105] : x[104];
  assign t[146] = t[176] ^ t[150];
  assign t[147] = t[177] ^ t[151];
  assign t[148] = t[101] ^ t[69];
  assign t[149] = t[140] ? x[107] : x[106];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[110] ? x[109] : x[108];
  assign t[151] = t[80] ? x[111] : x[110];
  assign t[152] = t[178] ^ x[4];
  assign t[153] = t[179] ^ x[7];
  assign t[154] = t[180] ^ x[12];
  assign t[155] = t[181] ^ x[15];
  assign t[156] = t[182] ^ x[18];
  assign t[157] = t[183] ^ x[21];
  assign t[158] = t[184] ^ x[24];
  assign t[159] = t[185] ^ x[27];
  assign t[15] = t[153] | t[29];
  assign t[160] = t[186] ^ x[30];
  assign t[161] = t[187] ^ x[33];
  assign t[162] = t[188] ^ x[36];
  assign t[163] = t[189] ^ x[39];
  assign t[164] = t[190] ^ x[42];
  assign t[165] = t[191] ^ x[45];
  assign t[166] = t[192] ^ x[48];
  assign t[167] = t[193] ^ x[51];
  assign t[168] = t[194] ^ x[54];
  assign t[169] = t[195] ^ x[57];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[196] ^ x[60];
  assign t[171] = t[197] ^ x[67];
  assign t[172] = t[198] ^ x[70];
  assign t[173] = t[199] ^ x[73];
  assign t[174] = t[200] ^ x[76];
  assign t[175] = t[201] ^ x[89];
  assign t[176] = t[202] ^ x[100];
  assign t[177] = t[203] ^ x[103];
  assign t[178] = (x[2] & x[3]);
  assign t[179] = (x[5] & x[6]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = (x[10] & x[11]);
  assign t[181] = (x[13] & x[14]);
  assign t[182] = (x[16] & x[17]);
  assign t[183] = (x[19] & x[20]);
  assign t[184] = (x[22] & x[23]);
  assign t[185] = (x[25] & x[26]);
  assign t[186] = (x[28] & x[29]);
  assign t[187] = (x[31] & x[32]);
  assign t[188] = (x[34] & x[35]);
  assign t[189] = (x[37] & x[38]);
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = (x[40] & x[41]);
  assign t[191] = (x[43] & x[44]);
  assign t[192] = (x[46] & x[47]);
  assign t[193] = (x[49] & x[50]);
  assign t[194] = (x[52] & x[53]);
  assign t[195] = (x[55] & x[56]);
  assign t[196] = (x[58] & x[59]);
  assign t[197] = (x[65] & x[66]);
  assign t[198] = (x[68] & x[69]);
  assign t[199] = (x[71] & x[72]);
  assign t[19] = t[35] ^ t[25];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[74] & x[75]);
  assign t[201] = (x[87] & x[88]);
  assign t[202] = (x[98] & x[99]);
  assign t[203] = (x[101] & x[102]);
  assign t[20] = t[36] & t[37];
  assign t[21] = t[38] ^ t[39];
  assign t[22] = t[40] & t[41];
  assign t[23] = t[42] ^ t[43];
  assign t[24] = t[44] ^ t[45];
  assign t[25] = t[46];
  assign t[26] = t[47] ^ t[48];
  assign t[27] = ~(t[29] & t[49]);
  assign t[28] = ~(t[154] ^ t[50]);
  assign t[29] = ~(t[51] & t[52]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[53]);
  assign t[31] = ~(t[155]);
  assign t[32] = ~(t[156]);
  assign t[33] = ~(t[157]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = ~t[56];
  assign t[36] = ~(t[57]);
  assign t[37] = t[3];
  assign t[38] = t[58] ? t[59] : t[158];
  assign t[39] = t[58] ? t[60] : t[159];
  assign t[3] = t[7] ? t[8] : t[152];
  assign t[40] = ~(t[21] ^ t[61]);
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] ^ t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] & t[71];
  assign t[46] = t[7] ? t[72] : t[160];
  assign t[47] = t[73] ^ t[20];
  assign t[48] = t[74] & t[75];
  assign t[49] = ~(t[76] & t[77]);
  assign t[4] = ~(t[9]);
  assign t[50] = t[78] ^ t[161];
  assign t[51] = ~(t[154]);
  assign t[52] = t[79] & t[78];
  assign t[53] = ~(t[80]);
  assign t[54] = ~(t[162]);
  assign t[55] = ~(t[81] & t[163]);
  assign t[56] = t[7] ? t[82] : t[164];
  assign t[57] = t[83];
  assign t[58] = ~(t[84]);
  assign t[59] = t[158] ^ t[85];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[159] ^ t[86];
  assign t[61] = t[87] ^ t[88];
  assign t[62] = t[39] ^ t[89];
  assign t[63] = t[58] ? t[90] : t[165];
  assign t[64] = t[157] ^ t[91];
  assign t[65] = t[162] ^ t[92];
  assign t[66] = t[93] ^ t[94];
  assign t[67] = t[95] & t[96];
  assign t[68] = t[58] ? t[97] : t[166];
  assign t[69] = t[58] ? t[98] : t[167];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = ~(t[44] ^ t[99]);
  assign t[71] = t[100] ^ t[101];
  assign t[72] = t[160] ^ t[102];
  assign t[73] = t[103] & t[104];
  assign t[74] = ~(t[105] ^ t[47]);
  assign t[75] = t[106] ^ t[37];
  assign t[76] = ~(t[79] | t[78]);
  assign t[77] = ~(t[107] | t[51]);
  assign t[78] = ~(t[168]);
  assign t[79] = ~(t[161]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[15]);
  assign t[81] = ~(t[169]);
  assign t[82] = t[164] ^ t[108];
  assign t[83] = t[7] ? t[109] : t[170];
  assign t[84] = ~(t[7]);
  assign t[85] = t[110] ? x[62] : x[61];
  assign t[86] = t[110] ? x[64] : x[63];
  assign t[87] = t[111] & t[112];
  assign t[88] = t[113] & t[63];
  assign t[89] = t[58] ? t[114] : t[171];
  assign t[8] = t[152] ^ t[16];
  assign t[90] = t[165] ^ t[115];
  assign t[91] = t[7] ? t[116] : t[172];
  assign t[92] = t[117] ? t[118] : t[173];
  assign t[93] = t[119] & t[120];
  assign t[94] = t[121] & t[122];
  assign t[95] = ~(t[93] ^ t[123]);
  assign t[96] = t[124] ^ t[125];
  assign t[97] = t[166] ^ t[126];
  assign t[98] = t[167] ^ t[127];
  assign t[99] = t[128] ^ t[129];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind128(x, y);
 input [111:0] x;
 output y;

 wire [214:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[131] ^ t[132];
  assign t[101] = t[104] ? x[72] : x[71];
  assign t[102] = t[178] ^ t[133];
  assign t[103] = t[104] ? x[74] : x[73];
  assign t[104] = ~(t[54]);
  assign t[105] = ~(t[134]);
  assign t[106] = ~(t[43]);
  assign t[107] = t[43] ^ t[71];
  assign t[108] = t[71] ^ t[25];
  assign t[109] = ~(t[164]);
  assign t[10] = t[19] ^ t[20];
  assign t[110] = ~(t[54]);
  assign t[111] = ~(t[135]);
  assign t[112] = ~(t[60]);
  assign t[113] = t[60] ^ t[89];
  assign t[114] = t[89] ^ t[35];
  assign t[115] = t[110] ? x[76] : x[75];
  assign t[116] = t[181] ^ t[136];
  assign t[117] = t[110] ? x[78] : x[77];
  assign t[118] = t[182] ^ t[137];
  assign t[119] = t[7] ? t[138] : t[184];
  assign t[11] = ~(t[21] ^ t[22]);
  assign t[120] = t[139] ^ t[140];
  assign t[121] = t[92] ^ t[141];
  assign t[122] = t[180] ^ t[142];
  assign t[123] = t[183] ^ t[143];
  assign t[124] = ~(t[144] ^ t[68]);
  assign t[125] = t[41] ^ t[129];
  assign t[126] = ~(t[132]);
  assign t[127] = ~(t[145]);
  assign t[128] = ~(t[67]);
  assign t[129] = t[146];
  assign t[12] = t[23] ^ t[24];
  assign t[130] = t[41] ^ t[145];
  assign t[131] = t[145] ^ t[65];
  assign t[132] = t[129] ^ t[67];
  assign t[133] = t[104] ? x[83] : x[82];
  assign t[134] = t[45] ^ t[71];
  assign t[135] = t[62] ^ t[89];
  assign t[136] = t[110] ? x[85] : x[84];
  assign t[137] = t[110] ? x[87] : x[86];
  assign t[138] = t[184] ^ t[147];
  assign t[139] = t[148] & t[149];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[150] & t[122];
  assign t[141] = t[174] ^ t[151];
  assign t[142] = t[7] ? t[152] : t[185];
  assign t[143] = t[82] ? x[92] : x[91];
  assign t[144] = t[145] ^ t[67];
  assign t[145] = ~t[153];
  assign t[146] = t[7] ? t[154] : t[186];
  assign t[147] = t[110] ? x[97] : x[96];
  assign t[148] = ~(t[155]);
  assign t[149] = ~(t[91]);
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = ~(t[92]);
  assign t[151] = t[156] ? t[157] : t[187];
  assign t[152] = t[185] ^ t[158];
  assign t[153] = t[7] ? t[159] : t[188];
  assign t[154] = t[186] ^ t[160];
  assign t[155] = t[122] ^ t[92];
  assign t[156] = ~(t[73]);
  assign t[157] = t[187] ^ t[161];
  assign t[158] = t[82] ? x[105] : x[104];
  assign t[159] = t[188] ^ t[162];
  assign t[15] = t[164] | t[29];
  assign t[160] = t[30] ? x[107] : x[106];
  assign t[161] = t[30] ? x[109] : x[108];
  assign t[162] = t[82] ? x[111] : x[110];
  assign t[163] = t[189] ^ x[4];
  assign t[164] = t[190] ^ x[7];
  assign t[165] = t[191] ^ x[12];
  assign t[166] = t[192] ^ x[15];
  assign t[167] = t[193] ^ x[18];
  assign t[168] = t[194] ^ x[21];
  assign t[169] = t[195] ^ x[24];
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = t[196] ^ x[27];
  assign t[171] = t[197] ^ x[30];
  assign t[172] = t[198] ^ x[33];
  assign t[173] = t[199] ^ x[36];
  assign t[174] = t[200] ^ x[39];
  assign t[175] = t[201] ^ x[42];
  assign t[176] = t[202] ^ x[45];
  assign t[177] = t[203] ^ x[48];
  assign t[178] = t[204] ^ x[51];
  assign t[179] = t[205] ^ x[56];
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = t[206] ^ x[59];
  assign t[181] = t[207] ^ x[64];
  assign t[182] = t[208] ^ x[67];
  assign t[183] = t[209] ^ x[70];
  assign t[184] = t[210] ^ x[81];
  assign t[185] = t[211] ^ x[90];
  assign t[186] = t[212] ^ x[95];
  assign t[187] = t[213] ^ x[100];
  assign t[188] = t[214] ^ x[103];
  assign t[189] = (x[2] & x[3]);
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = (x[5] & x[6]);
  assign t[191] = (x[10] & x[11]);
  assign t[192] = (x[13] & x[14]);
  assign t[193] = (x[16] & x[17]);
  assign t[194] = (x[19] & x[20]);
  assign t[195] = (x[22] & x[23]);
  assign t[196] = (x[25] & x[26]);
  assign t[197] = (x[28] & x[29]);
  assign t[198] = (x[31] & x[32]);
  assign t[199] = (x[34] & x[35]);
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[200] = (x[37] & x[38]);
  assign t[201] = (x[40] & x[41]);
  assign t[202] = (x[43] & x[44]);
  assign t[203] = (x[46] & x[47]);
  assign t[204] = (x[49] & x[50]);
  assign t[205] = (x[54] & x[55]);
  assign t[206] = (x[57] & x[58]);
  assign t[207] = (x[62] & x[63]);
  assign t[208] = (x[65] & x[66]);
  assign t[209] = (x[68] & x[69]);
  assign t[20] = t[37] ^ t[38];
  assign t[210] = (x[79] & x[80]);
  assign t[211] = (x[88] & x[89]);
  assign t[212] = (x[93] & x[94]);
  assign t[213] = (x[98] & x[99]);
  assign t[214] = (x[101] & x[102]);
  assign t[21] = ~(t[39] ^ t[40]);
  assign t[22] = t[41] ^ t[42];
  assign t[23] = t[43] ^ t[25];
  assign t[24] = t[44] & t[45];
  assign t[25] = t[46] ? t[47] : t[165];
  assign t[26] = t[48] ^ t[49];
  assign t[27] = ~(t[29] & t[50]);
  assign t[28] = ~(t[166] ^ t[51]);
  assign t[29] = ~(t[52] & t[53]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[54]);
  assign t[31] = ~(t[167]);
  assign t[32] = ~(t[168]);
  assign t[33] = ~(t[169]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = t[46] ? t[57] : t[170];
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[60] ^ t[35];
  assign t[38] = t[61] & t[62];
  assign t[39] = t[63] ^ t[64];
  assign t[3] = t[7] ? t[8] : t[163];
  assign t[40] = t[65] ^ t[66];
  assign t[41] = t[67] ^ t[65];
  assign t[42] = t[68] ^ t[69];
  assign t[43] = t[46] ? t[70] : t[171];
  assign t[44] = ~(t[71]);
  assign t[45] = t[46] ? t[72] : t[172];
  assign t[46] = ~(t[73]);
  assign t[47] = t[165] ^ t[74];
  assign t[48] = t[75] ^ t[24];
  assign t[49] = t[76] & t[77];
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[78] & t[79]);
  assign t[51] = t[80] ^ t[173];
  assign t[52] = ~(t[166]);
  assign t[53] = t[81] & t[80];
  assign t[54] = ~(t[82]);
  assign t[55] = ~(t[174]);
  assign t[56] = ~(t[83] & t[175]);
  assign t[57] = t[170] ^ t[84];
  assign t[58] = t[85] ^ t[38];
  assign t[59] = t[86] & t[87];
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[46] ? t[88] : t[176];
  assign t[61] = ~(t[89]);
  assign t[62] = t[46] ? t[90] : t[177];
  assign t[63] = t[91] ^ t[92];
  assign t[64] = t[93] & t[94];
  assign t[65] = t[95];
  assign t[66] = t[68] ^ t[96];
  assign t[67] = t[3];
  assign t[68] = t[97] ^ t[98];
  assign t[69] = t[99] & t[100];
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[171] ^ t[101];
  assign t[71] = t[46] ? t[102] : t[178];
  assign t[72] = t[172] ^ t[103];
  assign t[73] = ~(t[7]);
  assign t[74] = t[104] ? x[53] : x[52];
  assign t[75] = t[105] & t[106];
  assign t[76] = ~(t[107] ^ t[48]);
  assign t[77] = t[108] ^ t[45];
  assign t[78] = ~(t[81] | t[80]);
  assign t[79] = ~(t[109] | t[52]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[179]);
  assign t[81] = ~(t[173]);
  assign t[82] = ~(t[15]);
  assign t[83] = ~(t[180]);
  assign t[84] = t[110] ? x[61] : x[60];
  assign t[85] = t[111] & t[112];
  assign t[86] = ~(t[113] ^ t[58]);
  assign t[87] = t[114] ^ t[62];
  assign t[88] = t[176] ^ t[115];
  assign t[89] = t[46] ? t[116] : t[181];
  assign t[8] = t[163] ^ t[16];
  assign t[90] = t[177] ^ t[117];
  assign t[91] = t[7] ? t[118] : t[182];
  assign t[92] = t[169] ^ t[119];
  assign t[93] = ~(t[63] ^ t[120]);
  assign t[94] = t[121] ^ t[122];
  assign t[95] = t[7] ? t[123] : t[183];
  assign t[96] = t[124] & t[125];
  assign t[97] = t[126] & t[127];
  assign t[98] = t[128] & t[129];
  assign t[99] = ~(t[97] ^ t[130]);
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind129(x, y);
 input [111:0] x;
 output y;

 wire [192:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[100] = t[118] ^ t[23];
  assign t[101] = ~(t[115]);
  assign t[102] = ~(t[120]);
  assign t[103] = ~(t[121]);
  assign t[104] = ~(t[122]);
  assign t[105] = t[43] ? t[123] : t[160];
  assign t[106] = t[121] ^ t[122];
  assign t[107] = t[122] ^ t[25];
  assign t[108] = ~(t[142]);
  assign t[109] = t[124] ? x[71] : x[70];
  assign t[10] = t[19] ^ t[20];
  assign t[110] = ~t[125];
  assign t[111] = t[7] ? t[126] : t[161];
  assign t[112] = t[124] ? x[76] : x[75];
  assign t[113] = t[158] ^ t[127];
  assign t[114] = t[30] ? x[78] : x[77];
  assign t[115] = ~(t[30]);
  assign t[116] = t[98] ^ t[118];
  assign t[117] = t[43] ? t[128] : t[162];
  assign t[118] = t[43] ? t[129] : t[163];
  assign t[119] = t[159] ^ t[130];
  assign t[11] = t[21] ^ t[22];
  assign t[120] = t[105] ^ t[122];
  assign t[121] = t[43] ? t[131] : t[164];
  assign t[122] = t[43] ? t[132] : t[165];
  assign t[123] = t[160] ^ t[133];
  assign t[124] = ~(t[115]);
  assign t[125] = t[7] ? t[134] : t[166];
  assign t[126] = t[161] ^ t[135];
  assign t[127] = t[94] ? x[95] : x[94];
  assign t[128] = t[162] ^ t[136];
  assign t[129] = t[163] ^ t[137];
  assign t[12] = t[23] ^ t[24];
  assign t[130] = t[94] ? x[97] : x[96];
  assign t[131] = t[164] ^ t[138];
  assign t[132] = t[165] ^ t[139];
  assign t[133] = t[101] ? x[99] : x[98];
  assign t[134] = t[166] ^ t[140];
  assign t[135] = t[124] ? x[101] : x[100];
  assign t[136] = t[94] ? x[103] : x[102];
  assign t[137] = t[94] ? x[105] : x[104];
  assign t[138] = t[101] ? x[107] : x[106];
  assign t[139] = t[101] ? x[109] : x[108];
  assign t[13] = t[25] ^ t[26];
  assign t[140] = t[30] ? x[111] : x[110];
  assign t[141] = t[167] ^ x[4];
  assign t[142] = t[168] ^ x[7];
  assign t[143] = t[169] ^ x[12];
  assign t[144] = t[170] ^ x[15];
  assign t[145] = t[171] ^ x[18];
  assign t[146] = t[172] ^ x[21];
  assign t[147] = t[173] ^ x[24];
  assign t[148] = t[174] ^ x[27];
  assign t[149] = t[175] ^ x[30];
  assign t[14] = ~(t[27] & t[28]);
  assign t[150] = t[176] ^ x[33];
  assign t[151] = t[177] ^ x[36];
  assign t[152] = t[178] ^ x[39];
  assign t[153] = t[179] ^ x[42];
  assign t[154] = t[180] ^ x[45];
  assign t[155] = t[181] ^ x[48];
  assign t[156] = t[182] ^ x[51];
  assign t[157] = t[183] ^ x[58];
  assign t[158] = t[184] ^ x[63];
  assign t[159] = t[185] ^ x[66];
  assign t[15] = t[142] | t[29];
  assign t[160] = t[186] ^ x[69];
  assign t[161] = t[187] ^ x[74];
  assign t[162] = t[188] ^ x[81];
  assign t[163] = t[189] ^ x[84];
  assign t[164] = t[190] ^ x[87];
  assign t[165] = t[191] ^ x[90];
  assign t[166] = t[192] ^ x[93];
  assign t[167] = (x[2] & x[3]);
  assign t[168] = (x[5] & x[6]);
  assign t[169] = (x[10] & x[11]);
  assign t[16] = t[30] ? x[9] : x[8];
  assign t[170] = (x[13] & x[14]);
  assign t[171] = (x[16] & x[17]);
  assign t[172] = (x[19] & x[20]);
  assign t[173] = (x[22] & x[23]);
  assign t[174] = (x[25] & x[26]);
  assign t[175] = (x[28] & x[29]);
  assign t[176] = (x[31] & x[32]);
  assign t[177] = (x[34] & x[35]);
  assign t[178] = (x[37] & x[38]);
  assign t[179] = (x[40] & x[41]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[180] = (x[43] & x[44]);
  assign t[181] = (x[46] & x[47]);
  assign t[182] = (x[49] & x[50]);
  assign t[183] = (x[56] & x[57]);
  assign t[184] = (x[61] & x[62]);
  assign t[185] = (x[64] & x[65]);
  assign t[186] = (x[67] & x[68]);
  assign t[187] = (x[72] & x[73]);
  assign t[188] = (x[79] & x[80]);
  assign t[189] = (x[82] & x[83]);
  assign t[18] = ~(t[33] & t[34]);
  assign t[190] = (x[85] & x[86]);
  assign t[191] = (x[88] & x[89]);
  assign t[192] = (x[91] & x[92]);
  assign t[19] = t[35] ^ t[36];
  assign t[1] = ~(t[4]);
  assign t[20] = t[37] ^ t[38];
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[41] & t[42];
  assign t[23] = t[43] ? t[44] : t[143];
  assign t[24] = t[45] ^ t[46];
  assign t[25] = t[43] ? t[47] : t[144];
  assign t[26] = t[48] ^ t[49];
  assign t[27] = ~(t[29] & t[50]);
  assign t[28] = ~(t[145] ^ t[51]);
  assign t[29] = ~(t[52] & t[53]);
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = ~(t[15]);
  assign t[31] = ~(t[146]);
  assign t[32] = ~(t[147]);
  assign t[33] = ~(t[148]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = t[56];
  assign t[36] = t[3];
  assign t[37] = t[57] ^ t[58];
  assign t[38] = t[59] & t[60];
  assign t[39] = t[7] ? t[61] : t[149];
  assign t[3] = t[7] ? t[8] : t[141];
  assign t[40] = t[150] ^ t[62];
  assign t[41] = ~(t[63]);
  assign t[42] = t[151] ^ t[64];
  assign t[43] = ~(t[65]);
  assign t[44] = t[143] ^ t[66];
  assign t[45] = t[67] ^ t[68];
  assign t[46] = t[69] & t[70];
  assign t[47] = t[144] ^ t[71];
  assign t[48] = t[72] ^ t[73];
  assign t[49] = t[74] & t[75];
  assign t[4] = ~(t[9]);
  assign t[50] = ~(t[76] & t[77]);
  assign t[51] = t[78] ^ t[152];
  assign t[52] = ~(t[145]);
  assign t[53] = t[79] & t[78];
  assign t[54] = ~(t[150]);
  assign t[55] = ~(t[80] & t[153]);
  assign t[56] = t[7] ? t[81] : t[154];
  assign t[57] = t[82] & t[83];
  assign t[58] = t[84] & t[85];
  assign t[59] = ~(t[57] ^ t[86]);
  assign t[5] = t[10] ^ t[11];
  assign t[60] = t[87] ^ t[88];
  assign t[61] = t[149] ^ t[89];
  assign t[62] = t[90] ? t[91] : t[155];
  assign t[63] = t[148] ^ t[92];
  assign t[64] = t[7] ? t[93] : t[156];
  assign t[65] = ~(t[7]);
  assign t[66] = t[94] ? x[53] : x[52];
  assign t[67] = t[95] & t[96];
  assign t[68] = t[97] & t[98];
  assign t[69] = ~(t[99] ^ t[45]);
  assign t[6] = ~(t[12] ^ t[13]);
  assign t[70] = t[100] ^ t[98];
  assign t[71] = t[101] ? x[55] : x[54];
  assign t[72] = t[102] & t[103];
  assign t[73] = t[104] & t[105];
  assign t[74] = ~(t[106] ^ t[48]);
  assign t[75] = t[107] ^ t[105];
  assign t[76] = ~(t[79] | t[78]);
  assign t[77] = ~(t[108] | t[52]);
  assign t[78] = ~(t[157]);
  assign t[79] = ~(t[152]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[80] = ~(t[151]);
  assign t[81] = t[154] ^ t[109];
  assign t[82] = ~(t[88]);
  assign t[83] = ~(t[110]);
  assign t[84] = ~(t[35]);
  assign t[85] = t[111];
  assign t[86] = t[19] ^ t[110];
  assign t[87] = t[110] ^ t[36];
  assign t[88] = t[85] ^ t[35];
  assign t[89] = t[94] ? x[60] : x[59];
  assign t[8] = t[141] ^ t[16];
  assign t[90] = ~(t[65]);
  assign t[91] = t[155] ^ t[112];
  assign t[92] = t[7] ? t[113] : t[158];
  assign t[93] = t[156] ^ t[114];
  assign t[94] = ~(t[115]);
  assign t[95] = ~(t[116]);
  assign t[96] = ~(t[117]);
  assign t[97] = ~(t[118]);
  assign t[98] = t[43] ? t[119] : t[159];
  assign t[99] = t[117] ^ t[118];
  assign t[9] = ~(t[17] | t[18]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind130(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = t[2] ^ x[3];
  assign t[2] = (x[1] & x[2]);
  assign y = ~(t[0] | x[0]);
endmodule

module R1ind131(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = t[2] ^ x[3];
  assign t[2] = (x[1] & x[2]);
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind132(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = t[2] ^ x[3];
  assign t[2] = (x[1] & x[2]);
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind133(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = t[2] ^ x[3];
  assign t[2] = (x[1] & x[2]);
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind134(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = t[2] ^ x[3];
  assign t[2] = (x[1] & x[2]);
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind135(x, y);
 input [6:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[1] = ~(t[3]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[3];
  assign t[4] = t[6] ^ x[6];
  assign t[5] = (x[1] & x[2]);
  assign t[6] = (x[4] & x[5]);
  assign y = x[0] | t[0];
endmodule

module R1ind136(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = t[2] ^ x[3];
  assign t[2] = (x[1] & x[2]);
  assign y = ~(t[0] | x[0]);
endmodule

module R1ind137(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = t[2] ^ x[3];
  assign t[2] = (x[1] & x[2]);
  assign y = ~(t[0] | x[0]);
endmodule

module R1ind138(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = t[2] ^ x[3];
  assign t[2] = (x[1] & x[2]);
  assign y = ~(t[0] | x[0]);
endmodule

module R1ind139(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0] | x[3]);
endmodule

module R1_ind(x, y);
 input [417:0] x;
 output [139:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[8], x[7], x[6]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[11], x[10], x[9]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[14], x[13], x[12]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[17], x[16], x[15]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[20], x[19], x[18]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[23], x[22], x[21]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[26], x[25], x[24]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[29], x[28], x[27]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[32], x[31], x[30]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[35], x[34], x[33]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[38], x[37], x[36]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[41], x[40], x[39]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[44], x[43], x[42]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[47], x[46], x[45]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[50], x[49], x[48]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[53], x[52], x[51]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[56], x[55], x[54]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[59], x[58], x[57]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[62], x[61], x[60]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[65], x[64], x[63]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[68], x[67], x[66]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[71], x[70], x[69]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[74], x[73], x[72]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[77], x[76], x[75]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[80], x[79], x[78]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[83], x[82], x[81]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[86], x[85], x[84]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[89], x[88], x[87]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[92], x[91], x[90]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[95], x[94], x[93]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[98], x[97], x[96]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[101], x[100], x[99]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[104], x[103], x[102]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[107], x[106], x[105]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[110], x[109], x[108]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[113], x[112], x[111]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[116], x[115], x[114]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[119], x[118], x[117]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[122], x[121], x[120]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[125], x[124], x[123]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[128], x[127], x[126]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[131], x[130], x[129]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[134], x[133], x[132]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[137], x[136], x[135]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[140], x[139], x[138]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[143], x[142], x[141]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[146], x[145], x[144]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[149], x[148], x[147]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[152], x[151], x[150]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[155], x[154], x[153]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[158], x[157], x[156]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[161], x[160], x[159]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[164], x[163], x[162]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[167], x[166], x[165]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[170], x[169], x[168]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[173], x[172], x[171]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[176], x[175], x[174]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[179], x[178], x[177]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[182], x[181], x[180]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[185], x[184], x[183]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[188], x[187], x[186]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[191], x[190], x[189]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[194], x[193], x[192]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[2], x[1], x[0], x[195]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[260], x[259], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[119], x[118], x[117], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[116], x[115], x[114], x[56], x[55], x[54], x[113], x[112], x[111], x[122], x[121], x[120], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[47], x[46], x[45], x[59], x[58], x[57], x[62], x[61], x[60], x[53], x[52], x[51], x[41], x[40], x[39], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[44], x[43], x[42], x[50], x[49], x[48], x[198], x[197], x[196], x[222], x[221], x[220], x[179], x[178], x[177], x[173], x[172], x[171], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[176], x[175], x[174], x[182], x[181], x[180], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[216], x[215], x[194], x[193], x[192], x[214], x[195]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[248], x[247], x[246], x[245], x[260], x[259], x[256], x[255], x[258], x[257], x[59], x[58], x[57], x[252], x[251], x[233], x[232], x[240], x[239], x[62], x[61], x[60], x[231], x[230], x[119], x[118], x[117], x[254], x[253], x[244], x[243], x[56], x[55], x[54], x[226], x[225], x[224], x[223], x[250], x[249], x[238], x[237], x[236], x[235], x[234], x[116], x[115], x[114], x[242], x[241], x[122], x[121], x[120], x[179], x[178], x[177], x[44], x[43], x[42], x[229], x[228], x[227], x[173], x[172], x[171], x[113], x[112], x[111], x[53], x[52], x[51], x[176], x[175], x[174], x[182], x[181], x[180], x[47], x[46], x[45], x[50], x[49], x[48], x[198], x[197], x[196], x[222], x[221], x[220], x[41], x[40], x[39], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[263], x[262], x[191], x[190], x[189], x[261], x[195]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[248], x[247], x[250], x[249], x[238], x[237], x[240], x[239], x[258], x[257], x[246], x[245], x[242], x[241], x[244], x[243], x[256], x[255], x[260], x[259], x[233], x[232], x[224], x[223], x[254], x[253], x[59], x[58], x[57], x[47], x[46], x[45], x[50], x[49], x[48], x[252], x[251], x[44], x[43], x[42], x[226], x[225], x[116], x[115], x[114], x[236], x[235], x[234], x[62], x[61], x[60], x[41], x[40], x[39], x[53], x[52], x[51], x[56], x[55], x[54], x[119], x[118], x[117], x[179], x[178], x[177], x[182], x[181], x[180], x[229], x[228], x[227], x[113], x[112], x[111], x[122], x[121], x[120], x[231], x[230], x[176], x[175], x[174], x[198], x[197], x[196], x[222], x[221], x[220], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[173], x[172], x[171], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[266], x[265], x[188], x[187], x[186], x[264], x[195]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[260], x[259], x[258], x[257], x[224], x[223], x[238], x[237], x[250], x[249], x[252], x[251], x[233], x[232], x[256], x[255], x[119], x[118], x[117], x[248], x[247], x[244], x[243], x[246], x[245], x[116], x[115], x[114], x[182], x[181], x[180], x[50], x[49], x[48], x[236], x[235], x[234], x[254], x[253], x[47], x[46], x[45], x[242], x[241], x[240], x[239], x[122], x[121], x[120], x[179], x[178], x[177], x[226], x[225], x[56], x[55], x[54], x[229], x[228], x[227], x[231], x[230], x[59], x[58], x[57], x[53], x[52], x[51], x[62], x[61], x[60], x[198], x[197], x[196], x[222], x[221], x[220], x[113], x[112], x[111], x[41], x[40], x[39], x[44], x[43], x[42], x[176], x[175], x[174], x[207], x[206], x[205], x[219], x[218], x[217], x[201], x[200], x[199], x[173], x[172], x[171], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[269], x[268], x[185], x[184], x[183], x[267], x[195]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[107], x[106], x[105], x[110], x[109], x[108], x[290], x[289], x[288], x[287], x[286], x[285], x[284], x[283], x[282], x[281], x[104], x[103], x[102], x[280], x[279], x[278], x[277], x[101], x[100], x[99], x[276], x[275], x[236], x[235], x[234], x[274], x[273], x[35], x[34], x[33], x[92], x[91], x[90], x[29], x[28], x[27], x[229], x[228], x[227], x[167], x[166], x[165], x[272], x[271], x[161], x[160], x[159], x[32], x[31], x[30], x[38], x[37], x[36], x[95], x[94], x[93], x[98], x[97], x[96], x[89], x[88], x[87], x[222], x[221], x[220], x[198], x[197], x[196], x[164], x[163], x[162], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[170], x[169], x[168], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[224], x[223], x[182], x[181], x[180], x[270], x[195]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[302], x[301], x[280], x[279], x[300], x[299], x[288], x[287], x[278], x[277], x[286], x[285], x[298], x[297], x[292], x[291], x[274], x[273], x[284], x[283], x[107], x[106], x[105], x[296], x[295], x[95], x[94], x[93], x[110], x[109], x[108], x[167], x[166], x[165], x[272], x[271], x[294], x[293], x[282], x[281], x[236], x[235], x[234], x[98], x[97], x[96], x[161], x[160], x[159], x[104], x[103], x[102], x[276], x[275], x[290], x[289], x[92], x[91], x[90], x[164], x[163], x[162], x[32], x[31], x[30], x[229], x[228], x[227], x[101], x[100], x[99], x[170], x[169], x[168], x[35], x[34], x[33], x[38], x[37], x[36], x[198], x[197], x[196], x[222], x[221], x[220], x[89], x[88], x[87], x[29], x[28], x[27], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[233], x[232], x[179], x[178], x[177], x[303], x[195]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[294], x[293], x[282], x[281], x[284], x[283], x[298], x[297], x[288], x[287], x[280], x[279], x[290], x[289], x[302], x[301], x[300], x[299], x[274], x[273], x[272], x[271], x[296], x[295], x[278], x[277], x[35], x[34], x[33], x[38], x[37], x[36], x[276], x[275], x[292], x[291], x[32], x[31], x[30], x[104], x[103], x[102], x[167], x[166], x[165], x[236], x[235], x[234], x[95], x[94], x[93], x[29], x[28], x[27], x[107], x[106], x[105], x[110], x[109], x[108], x[286], x[285], x[164], x[163], x[162], x[170], x[169], x[168], x[229], x[228], x[227], x[101], x[100], x[99], x[98], x[97], x[96], x[89], x[88], x[87], x[92], x[91], x[90], x[198], x[197], x[196], x[222], x[221], x[220], x[161], x[160], x[159], x[201], x[200], x[199], x[219], x[218], x[217], x[207], x[206], x[205], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[226], x[225], x[176], x[175], x[174], x[304], x[195]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[302], x[301], x[298], x[297], x[300], x[299], x[288], x[287], x[272], x[271], x[282], x[281], x[294], x[293], x[107], x[106], x[105], x[104], x[103], x[102], x[110], x[109], x[108], x[167], x[166], x[165], x[274], x[273], x[292], x[291], x[170], x[169], x[168], x[38], x[37], x[36], x[236], x[235], x[234], x[296], x[295], x[286], x[285], x[280], x[279], x[276], x[275], x[278], x[277], x[35], x[34], x[33], x[290], x[289], x[284], x[283], x[229], x[228], x[227], x[164], x[163], x[162], x[92], x[91], x[90], x[198], x[197], x[196], x[222], x[221], x[220], x[101], x[100], x[99], x[161], x[160], x[159], x[95], x[94], x[93], x[89], x[88], x[87], x[98], x[97], x[96], x[29], x[28], x[27], x[32], x[31], x[30], x[201], x[200], x[199], x[219], x[218], x[217], x[207], x[206], x[205], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[231], x[230], x[173], x[172], x[171], x[305], x[195]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[338], x[337], x[336], x[335], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[322], x[321], x[320], x[319], x[23], x[22], x[21], x[318], x[317], x[316], x[315], x[314], x[313], x[143], x[142], x[141], x[146], x[145], x[144], x[312], x[311], x[17], x[16], x[15], x[236], x[235], x[234], x[310], x[309], x[308], x[307], x[20], x[19], x[18], x[140], x[139], x[138], x[80], x[79], x[78], x[137], x[136], x[135], x[229], x[228], x[227], x[155], x[154], x[153], x[149], x[148], x[147], x[26], x[25], x[24], x[83], x[82], x[81], x[86], x[85], x[84], x[77], x[76], x[75], x[198], x[197], x[196], x[222], x[221], x[220], x[152], x[151], x[150], x[158], x[157], x[156], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[272], x[271], x[170], x[169], x[168], x[306], x[195]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[316], x[315], x[322], x[321], x[330], x[329], x[314], x[313], x[320], x[319], x[336], x[335], x[334], x[333], x[326], x[325], x[310], x[309], x[308], x[307], x[338], x[337], x[328], x[327], x[83], x[82], x[81], x[332], x[331], x[155], x[154], x[153], x[20], x[19], x[18], x[318], x[317], x[236], x[235], x[234], x[86], x[85], x[84], x[149], x[148], x[147], x[143], x[142], x[141], x[324], x[323], x[312], x[311], x[146], x[145], x[144], x[80], x[79], x[78], x[152], x[151], x[150], x[158], x[157], x[156], x[23], x[22], x[21], x[229], x[228], x[227], x[140], x[139], x[138], x[17], x[16], x[15], x[26], x[25], x[24], x[198], x[197], x[196], x[222], x[221], x[220], x[137], x[136], x[135], x[77], x[76], x[75], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[288], x[287], x[167], x[166], x[165], x[339], x[195]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[338], x[337], x[330], x[329], x[332], x[331], x[318], x[317], x[322], x[321], x[308], x[307], x[316], x[315], x[23], x[22], x[21], x[20], x[19], x[18], x[310], x[309], x[328], x[327], x[314], x[313], x[17], x[16], x[15], x[26], x[25], x[24], x[312], x[311], x[326], x[325], x[336], x[335], x[334], x[333], x[155], x[154], x[153], x[158], x[157], x[156], x[236], x[235], x[234], x[324], x[323], x[83], x[82], x[81], x[320], x[319], x[152], x[151], x[150], x[140], x[139], x[138], x[229], x[228], x[227], x[86], x[85], x[84], x[77], x[76], x[75], x[80], x[79], x[78], x[143], x[142], x[141], x[146], x[145], x[144], x[222], x[221], x[220], x[137], x[136], x[135], x[149], x[148], x[147], x[219], x[218], x[217], x[198], x[197], x[196], x[201], x[200], x[199], x[207], x[206], x[205], x[274], x[273], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[164], x[163], x[162], x[340], x[195]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[308], x[307], x[338], x[337], x[322], x[321], x[318], x[317], x[336], x[335], x[328], x[327], x[334], x[333], x[158], x[157], x[156], x[23], x[22], x[21], x[332], x[331], x[330], x[329], x[155], x[154], x[153], x[310], x[309], x[326], x[325], x[26], x[25], x[24], x[236], x[235], x[234], x[143], x[142], x[141], x[320], x[319], x[316], x[315], x[312], x[311], x[314], x[313], x[140], x[139], x[138], x[146], x[145], x[144], x[229], x[228], x[227], x[324], x[323], x[17], x[16], x[15], x[20], x[19], x[18], x[152], x[151], x[150], x[80], x[79], x[78], x[222], x[221], x[220], x[149], x[148], x[147], x[83], x[82], x[81], x[77], x[76], x[75], x[86], x[85], x[84], x[219], x[218], x[217], x[137], x[136], x[135], x[198], x[197], x[196], x[201], x[200], x[199], x[207], x[206], x[205], x[286], x[285], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[161], x[160], x[159], x[341], x[195]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[366], x[365], x[364], x[363], x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[352], x[351], x[350], x[349], x[348], x[347], x[346], x[345], x[11], x[10], x[9], x[68], x[67], x[66], x[344], x[343], x[131], x[130], x[129], x[134], x[133], x[132], x[5], x[4], x[3], x[236], x[235], x[234], x[263], x[262], x[269], x[268], x[8], x[7], x[6], x[14], x[13], x[12], x[128], x[127], x[126], x[71], x[70], x[69], x[125], x[124], x[123], x[65], x[64], x[63], x[229], x[228], x[227], x[266], x[265], x[216], x[215], x[74], x[73], x[72], x[222], x[221], x[220], x[191], x[190], x[189], x[185], x[184], x[183], x[219], x[218], x[217], x[188], x[187], x[186], x[194], x[193], x[192], x[198], x[197], x[196], x[201], x[200], x[199], x[207], x[206], x[205], x[308], x[307], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[158], x[157], x[156], x[342], x[195]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[350], x[349], x[364], x[363], x[356], x[355], x[344], x[343], x[362], x[361], x[71], x[70], x[69], x[360], x[359], x[263], x[262], x[366], x[365], x[354], x[353], x[269], x[268], x[352], x[351], x[346], x[345], x[358], x[357], x[68], x[67], x[66], x[266], x[265], x[216], x[215], x[8], x[7], x[6], x[74], x[73], x[72], x[131], x[130], x[129], x[348], x[347], x[134], x[133], x[132], x[191], x[190], x[189], x[11], x[10], x[9], x[14], x[13], x[12], x[185], x[184], x[183], x[128], x[127], x[126], x[65], x[64], x[63], x[5], x[4], x[3], x[188], x[187], x[186], x[194], x[193], x[192], x[236], x[235], x[234], x[125], x[124], x[123], x[229], x[228], x[227], x[198], x[197], x[196], x[222], x[221], x[220], x[201], x[200], x[199], x[207], x[206], x[205], x[322], x[321], x[219], x[218], x[217], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[155], x[154], x[153], x[367], x[195]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[366], x[365], x[354], x[353], x[356], x[355], x[350], x[349], x[358], x[357], x[11], x[10], x[9], x[14], x[13], x[12], x[346], x[345], x[364], x[363], x[8], x[7], x[6], x[352], x[351], x[263], x[262], x[216], x[215], x[71], x[70], x[69], x[344], x[343], x[5], x[4], x[3], x[362], x[361], x[360], x[359], x[266], x[265], x[236], x[235], x[234], x[348], x[347], x[65], x[64], x[63], x[68], x[67], x[66], x[128], x[127], x[126], x[191], x[190], x[189], x[194], x[193], x[192], x[229], x[228], x[227], x[74], x[73], x[72], x[131], x[130], x[129], x[134], x[133], x[132], x[269], x[268], x[188], x[187], x[186], x[222], x[221], x[220], x[125], x[124], x[123], x[219], x[218], x[217], x[185], x[184], x[183], x[198], x[197], x[196], x[201], x[200], x[199], x[207], x[206], x[205], x[310], x[309], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[152], x[151], x[150], x[368], x[195]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[354], x[353], x[366], x[365], x[216], x[215], x[362], x[361], x[352], x[351], x[360], x[359], x[263], x[262], x[364], x[363], x[14], x[13], x[12], x[350], x[349], x[346], x[345], x[11], x[10], x[9], x[358], x[357], x[356], x[355], x[194], x[193], x[192], x[236], x[235], x[234], x[131], x[130], x[129], x[344], x[343], x[128], x[127], x[126], x[134], x[133], x[132], x[191], x[190], x[189], x[266], x[265], x[68], x[67], x[66], x[229], x[228], x[227], x[348], x[347], x[269], x[268], x[71], x[70], x[69], x[65], x[64], x[63], x[5], x[4], x[3], x[8], x[7], x[6], x[222], x[221], x[220], x[74], x[73], x[72], x[188], x[187], x[186], x[219], x[218], x[217], x[125], x[124], x[123], x[185], x[184], x[183], x[198], x[197], x[196], x[201], x[200], x[199], x[207], x[206], x[205], x[320], x[319], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[149], x[148], x[147], x[369], x[195]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[256], x[255], x[254], x[253], x[240], x[239], x[248], x[247], x[244], x[243], x[246], x[245], x[260], x[259], x[233], x[232], x[250], x[249], x[238], x[237], x[226], x[225], x[224], x[223], x[56], x[55], x[54], x[236], x[235], x[234], x[113], x[112], x[111], x[258], x[257], x[242], x[241], x[44], x[43], x[42], x[59], x[58], x[57], x[53], x[52], x[51], x[62], x[61], x[60], x[229], x[228], x[227], x[119], x[118], x[117], x[252], x[251], x[179], x[178], x[177], x[47], x[46], x[45], x[50], x[49], x[48], x[176], x[175], x[174], x[182], x[181], x[180], x[222], x[221], x[220], x[116], x[115], x[114], x[231], x[230], x[41], x[40], x[39], x[219], x[218], x[217], x[122], x[121], x[120], x[198], x[197], x[196], x[173], x[172], x[171], x[201], x[200], x[199], x[207], x[206], x[205], x[334], x[333], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[146], x[145], x[144], x[370], x[195]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[260], x[259], x[248], x[247], x[254], x[253], x[238], x[237], x[258], x[257], x[250], x[249], x[256], x[255], x[246], x[245], x[224], x[223], x[119], x[118], x[117], x[252], x[251], x[59], x[58], x[57], x[233], x[232], x[236], x[235], x[234], x[113], x[112], x[111], x[50], x[49], x[48], x[116], x[115], x[114], x[244], x[243], x[47], x[46], x[45], x[240], x[239], x[242], x[241], x[56], x[55], x[54], x[62], x[61], x[60], x[182], x[181], x[180], x[229], x[228], x[227], x[122], x[121], x[120], x[179], x[178], x[177], x[231], x[230], x[226], x[225], x[198], x[197], x[196], x[222], x[221], x[220], x[53], x[52], x[51], x[44], x[43], x[42], x[41], x[40], x[39], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[173], x[172], x[171], x[176], x[175], x[174], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[336], x[335], x[143], x[142], x[141], x[371], x[195]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[248], x[247], x[250], x[249], x[240], x[239], x[238], x[237], x[246], x[245], x[242], x[241], x[244], x[243], x[256], x[255], x[260], x[259], x[59], x[58], x[57], x[47], x[46], x[45], x[252], x[251], x[258], x[257], x[233], x[232], x[44], x[43], x[42], x[50], x[49], x[48], x[236], x[235], x[234], x[62], x[61], x[60], x[41], x[40], x[39], x[231], x[230], x[53], x[52], x[51], x[56], x[55], x[54], x[119], x[118], x[117], x[254], x[253], x[226], x[225], x[224], x[223], x[229], x[228], x[227], x[122], x[121], x[120], x[116], x[115], x[114], x[179], x[178], x[177], x[198], x[197], x[196], x[222], x[221], x[220], x[173], x[172], x[171], x[113], x[112], x[111], x[176], x[175], x[174], x[182], x[181], x[180], x[207], x[206], x[205], x[219], x[218], x[217], x[201], x[200], x[199], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[328], x[327], x[140], x[139], x[138], x[372], x[195]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[248], x[247], x[250], x[249], x[244], x[243], x[260], x[259], x[252], x[251], x[256], x[255], x[246], x[245], x[242], x[241], x[240], x[239], x[238], x[237], x[59], x[58], x[57], x[236], x[235], x[234], x[47], x[46], x[45], x[53], x[52], x[51], x[119], x[118], x[117], x[122], x[121], x[120], x[254], x[253], x[258], x[257], x[56], x[55], x[54], x[62], x[61], x[60], x[41], x[40], x[39], x[226], x[225], x[229], x[228], x[227], x[44], x[43], x[42], x[50], x[49], x[48], x[233], x[232], x[231], x[230], x[224], x[223], x[198], x[197], x[196], x[222], x[221], x[220], x[113], x[112], x[111], x[116], x[115], x[114], x[176], x[175], x[174], x[207], x[206], x[205], x[219], x[218], x[217], x[201], x[200], x[199], x[179], x[178], x[177], x[173], x[172], x[171], x[182], x[181], x[180], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[324], x[323], x[137], x[136], x[135], x[373], x[195]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[296], x[295], x[288], x[287], x[284], x[283], x[274], x[273], x[292], x[291], x[302], x[301], x[294], x[293], x[282], x[281], x[272], x[271], x[280], x[279], x[276], x[275], x[278], x[277], x[236], x[235], x[234], x[101], x[100], x[99], x[298], x[297], x[300], x[299], x[167], x[166], x[165], x[290], x[289], x[32], x[31], x[30], x[164], x[163], x[162], x[92], x[91], x[90], x[229], x[228], x[227], x[107], x[106], x[105], x[286], x[285], x[35], x[34], x[33], x[38], x[37], x[36], x[170], x[169], x[168], x[95], x[94], x[93], x[89], x[88], x[87], x[98], x[97], x[96], x[222], x[221], x[220], x[104], x[103], x[102], x[110], x[109], x[108], x[29], x[28], x[27], x[219], x[218], x[217], x[161], x[160], x[159], x[198], x[197], x[196], x[201], x[200], x[199], x[207], x[206], x[205], x[360], x[359], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[134], x[133], x[132], x[374], x[195]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[302], x[301], x[296], x[295], x[282], x[281], x[298], x[297], x[300], x[299], x[294], x[293], x[280], x[279], x[288], x[287], x[272], x[271], x[107], x[106], x[105], x[292], x[291], x[278], x[277], x[236], x[235], x[234], x[101], x[100], x[99], x[38], x[37], x[36], x[104], x[103], x[102], x[110], x[109], x[108], x[35], x[34], x[33], x[284], x[283], x[290], x[289], x[95], x[94], x[93], x[167], x[166], x[165], x[170], x[169], x[168], x[286], x[285], x[274], x[273], x[229], x[228], x[227], x[276], x[275], x[92], x[91], x[90], x[98], x[97], x[96], x[198], x[197], x[196], x[222], x[221], x[220], x[32], x[31], x[30], x[29], x[28], x[27], x[161], x[160], x[159], x[164], x[163], x[162], x[201], x[200], x[199], x[219], x[218], x[217], x[89], x[88], x[87], x[207], x[206], x[205], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[362], x[361], x[131], x[130], x[129], x[375], x[195]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[294], x[293], x[284], x[283], x[282], x[281], x[280], x[279], x[290], x[289], x[302], x[301], x[300], x[299], x[288], x[287], x[278], x[277], x[35], x[34], x[33], x[286], x[285], x[276], x[275], x[292], x[291], x[298], x[297], x[274], x[273], x[32], x[31], x[30], x[38], x[37], x[36], x[236], x[235], x[234], x[95], x[94], x[93], x[29], x[28], x[27], x[107], x[106], x[105], x[110], x[109], x[108], x[296], x[295], x[167], x[166], x[165], x[272], x[271], x[229], x[228], x[227], x[98], x[97], x[96], x[161], x[160], x[159], x[89], x[88], x[87], x[92], x[91], x[90], x[104], x[103], x[102], x[164], x[163], x[162], x[198], x[197], x[196], x[222], x[221], x[220], x[101], x[100], x[99], x[170], x[169], x[168], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[352], x[351], x[128], x[127], x[126], x[376], x[195]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[300], x[299], x[294], x[293], x[302], x[301], x[280], x[279], x[290], x[289], x[284], x[283], x[282], x[281], x[276], x[275], x[110], x[109], x[108], x[292], x[291], x[278], x[277], x[274], x[273], x[236], x[235], x[234], x[35], x[34], x[33], x[107], x[106], x[105], x[296], x[295], x[298], x[297], x[95], x[94], x[93], x[29], x[28], x[27], x[288], x[287], x[286], x[285], x[229], x[228], x[227], x[32], x[31], x[30], x[38], x[37], x[36], x[89], x[88], x[87], x[92], x[91], x[90], x[98], x[97], x[96], x[164], x[163], x[162], x[272], x[271], x[222], x[221], x[220], x[101], x[100], x[99], x[104], x[103], x[102], x[167], x[166], x[165], x[161], x[160], x[159], x[201], x[200], x[199], x[219], x[218], x[217], x[198], x[197], x[196], x[207], x[206], x[205], x[170], x[169], x[168], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[348], x[347], x[125], x[124], x[123], x[377], x[195]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[330], x[329], x[322], x[321], x[338], x[337], x[310], x[309], x[308], x[307], x[326], x[325], x[324], x[323], x[332], x[331], x[20], x[19], x[18], x[318], x[317], x[316], x[315], x[312], x[311], x[314], x[313], x[236], x[235], x[234], x[336], x[335], x[155], x[154], x[153], x[23], x[22], x[21], x[152], x[151], x[150], x[158], x[157], x[156], x[80], x[79], x[78], x[229], x[228], x[227], x[137], x[136], x[135], x[328], x[327], x[334], x[333], x[320], x[319], x[17], x[16], x[15], x[26], x[25], x[24], x[83], x[82], x[81], x[77], x[76], x[75], x[86], x[85], x[84], x[198], x[197], x[196], x[222], x[221], x[220], x[143], x[142], x[141], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[140], x[139], x[138], x[146], x[145], x[144], x[149], x[148], x[147], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[252], x[251], x[122], x[121], x[120], x[378], x[195]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[338], x[337], x[308], x[307], x[318], x[317], x[336], x[335], x[316], x[315], x[322], x[321], x[324], x[323], x[328], x[327], x[334], x[333], x[23], x[22], x[21], x[330], x[329], x[332], x[331], x[326], x[325], x[314], x[313], x[158], x[157], x[156], x[236], x[235], x[234], x[26], x[25], x[24], x[143], x[142], x[141], x[83], x[82], x[81], x[155], x[154], x[153], x[320], x[319], x[310], x[309], x[229], x[228], x[227], x[137], x[136], x[135], x[140], x[139], x[138], x[146], x[145], x[144], x[312], x[311], x[20], x[19], x[18], x[17], x[16], x[15], x[80], x[79], x[78], x[86], x[85], x[84], x[198], x[197], x[196], x[222], x[221], x[220], x[149], x[148], x[147], x[152], x[151], x[150], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[77], x[76], x[75], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[260], x[259], x[119], x[118], x[117], x[379], x[195]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[338], x[337], x[330], x[329], x[332], x[331], x[318], x[317], x[316], x[315], x[23], x[22], x[21], x[322], x[321], x[20], x[19], x[18], x[314], x[313], x[17], x[16], x[15], x[320], x[319], x[312], x[311], x[326], x[325], x[336], x[335], x[334], x[333], x[310], x[309], x[308], x[307], x[26], x[25], x[24], x[83], x[82], x[81], x[328], x[327], x[155], x[154], x[153], x[86], x[85], x[84], x[149], x[148], x[147], x[77], x[76], x[75], x[80], x[79], x[78], x[143], x[142], x[141], x[146], x[145], x[144], x[324], x[323], x[152], x[151], x[150], x[158], x[157], x[156], x[198], x[197], x[196], x[236], x[235], x[234], x[140], x[139], x[138], x[201], x[200], x[199], x[207], x[206], x[205], x[229], x[228], x[227], x[137], x[136], x[135], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[258], x[257], x[219], x[218], x[217], x[116], x[115], x[114], x[380], x[195]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[338], x[337], x[332], x[331], x[330], x[329], x[334], x[333], x[316], x[315], x[23], x[22], x[21], x[318], x[317], x[312], x[311], x[336], x[335], x[326], x[325], x[314], x[313], x[17], x[16], x[15], x[310], x[309], x[236], x[235], x[234], x[20], x[19], x[18], x[146], x[145], x[144], x[83], x[82], x[81], x[322], x[321], x[320], x[319], x[308], x[307], x[229], x[228], x[227], x[26], x[25], x[24], x[77], x[76], x[75], x[143], x[142], x[141], x[324], x[323], x[328], x[327], x[80], x[79], x[78], x[86], x[85], x[84], x[152], x[151], x[150], x[198], x[197], x[196], x[222], x[221], x[220], x[155], x[154], x[153], x[149], x[148], x[147], x[158], x[157], x[156], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[137], x[136], x[135], x[140], x[139], x[138], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[254], x[253], x[113], x[112], x[111], x[381], x[195]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[356], x[355], x[364], x[363], x[366], x[365], x[354], x[353], x[350], x[349], x[346], x[345], x[348], x[347], x[263], x[262], x[358], x[357], x[8], x[7], x[6], x[266], x[265], x[216], x[215], x[68], x[67], x[66], x[344], x[343], x[236], x[235], x[234], x[362], x[361], x[11], x[10], x[9], x[14], x[13], x[12], x[71], x[70], x[69], x[65], x[64], x[63], x[229], x[228], x[227], x[125], x[124], x[123], x[352], x[351], x[360], x[359], x[191], x[190], x[189], x[5], x[4], x[3], x[188], x[187], x[186], x[194], x[193], x[192], x[74], x[73], x[72], x[198], x[197], x[196], x[222], x[221], x[220], x[131], x[130], x[129], x[269], x[268], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[128], x[127], x[126], x[134], x[133], x[132], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[185], x[184], x[183], x[300], x[299], x[110], x[109], x[108], x[382], x[195]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[354], x[353], x[366], x[365], x[350], x[349], x[362], x[361], x[364], x[363], x[216], x[215], x[348], x[347], x[14], x[13], x[12], x[352], x[351], x[360], x[359], x[11], x[10], x[9], x[356], x[355], x[358], x[357], x[71], x[70], x[69], x[344], x[343], x[263], x[262], x[236], x[235], x[234], x[131], x[130], x[129], x[346], x[345], x[68], x[67], x[66], x[194], x[193], x[192], x[229], x[228], x[227], x[125], x[124], x[123], x[128], x[127], x[126], x[134], x[133], x[132], x[8], x[7], x[6], x[5], x[4], x[3], x[74], x[73], x[72], x[191], x[190], x[189], x[269], x[268], x[266], x[265], x[198], x[197], x[196], x[222], x[221], x[220], x[65], x[64], x[63], x[201], x[200], x[199], x[219], x[218], x[217], x[207], x[206], x[205], x[185], x[184], x[183], x[188], x[187], x[186], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[302], x[301], x[107], x[106], x[105], x[383], x[195]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[366], x[365], x[356], x[355], x[354], x[353], x[350], x[349], x[358], x[357], x[11], x[10], x[9], x[346], x[345], x[364], x[363], x[8], x[7], x[6], x[14], x[13], x[12], x[71], x[70], x[69], x[344], x[343], x[5], x[4], x[3], x[362], x[361], x[360], x[359], x[263], x[262], x[236], x[235], x[234], x[269], x[268], x[65], x[64], x[63], x[68], x[67], x[66], x[352], x[351], x[266], x[265], x[216], x[215], x[229], x[228], x[227], x[74], x[73], x[72], x[131], x[130], x[129], x[134], x[133], x[132], x[348], x[347], x[191], x[190], x[189], x[198], x[197], x[196], x[222], x[221], x[220], x[185], x[184], x[183], x[128], x[127], x[126], x[188], x[187], x[186], x[194], x[193], x[192], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[125], x[124], x[123], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[298], x[297], x[104], x[103], x[102], x[384], x[195]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[366], x[365], x[350], x[349], x[358], x[357], x[356], x[355], x[354], x[353], x[346], x[345], x[360], x[359], x[364], x[363], x[11], x[10], x[9], x[362], x[361], x[71], x[70], x[69], x[344], x[343], x[5], x[4], x[3], x[236], x[235], x[234], x[8], x[7], x[6], x[14], x[13], x[12], x[65], x[64], x[63], x[134], x[133], x[132], x[68], x[67], x[66], x[266], x[265], x[229], x[228], x[227], x[131], x[130], x[129], x[348], x[347], x[352], x[351], x[74], x[73], x[72], x[263], x[262], x[269], x[268], x[216], x[215], x[198], x[197], x[196], x[222], x[221], x[220], x[188], x[187], x[186], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[125], x[124], x[123], x[128], x[127], x[126], x[191], x[190], x[189], x[185], x[184], x[183], x[194], x[193], x[192], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[296], x[295], x[101], x[100], x[99], x[385], x[195]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[258], x[257], x[260], x[259], x[244], x[243], x[252], x[251], x[240], x[239], x[233], x[232], x[248], x[247], x[116], x[115], x[114], x[224], x[223], x[250], x[249], x[238], x[237], x[236], x[235], x[234], x[119], x[118], x[117], x[53], x[52], x[51], x[256], x[255], x[246], x[245], x[242], x[241], x[122], x[121], x[120], x[44], x[43], x[42], x[229], x[228], x[227], x[254], x[253], x[179], x[178], x[177], x[231], x[230], x[226], x[225], x[59], x[58], x[57], x[182], x[181], x[180], x[47], x[46], x[45], x[50], x[49], x[48], x[198], x[197], x[196], x[222], x[221], x[220], x[56], x[55], x[54], x[62], x[61], x[60], x[41], x[40], x[39], x[207], x[206], x[205], x[219], x[218], x[217], x[113], x[112], x[111], x[173], x[172], x[171], x[176], x[175], x[174], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[201], x[200], x[199], x[278], x[277], x[98], x[97], x[96], x[386], x[195]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[238], x[237], x[250], x[249], x[50], x[49], x[48], x[260], x[259], x[47], x[46], x[45], x[240], x[239], x[242], x[241], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[231], x[230], x[236], x[235], x[234], x[233], x[232], x[248], x[247], x[244], x[243], x[246], x[245], x[119], x[118], x[117], x[44], x[43], x[42], x[41], x[40], x[39], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[116], x[115], x[114], x[56], x[55], x[54], x[113], x[112], x[111], x[122], x[121], x[120], x[173], x[172], x[171], x[198], x[197], x[196], x[222], x[221], x[220], x[179], x[178], x[177], x[59], x[58], x[57], x[53], x[52], x[51], x[62], x[61], x[60], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[176], x[175], x[174], x[182], x[181], x[180], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[280], x[279], x[95], x[94], x[93], x[387], x[195]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[246], x[245], x[250], x[249], x[260], x[259], x[248], x[247], x[254], x[253], x[242], x[241], x[240], x[239], x[238], x[237], x[258], x[257], x[256], x[255], x[62], x[61], x[60], x[47], x[46], x[45], x[119], x[118], x[117], x[252], x[251], x[59], x[58], x[57], x[236], x[235], x[234], x[113], x[112], x[111], x[41], x[40], x[39], x[44], x[43], x[42], x[50], x[49], x[48], x[116], x[115], x[114], x[56], x[55], x[54], x[244], x[243], x[226], x[225], x[229], x[228], x[227], x[122], x[121], x[120], x[233], x[232], x[224], x[223], x[198], x[197], x[196], x[222], x[221], x[220], x[53], x[52], x[51], x[176], x[175], x[174], x[231], x[230], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[179], x[178], x[177], x[182], x[181], x[180], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[173], x[172], x[171], x[292], x[291], x[92], x[91], x[90], x[388], x[195]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[242], x[241], x[246], x[245], x[224], x[223], x[250], x[249], x[248], x[247], x[233], x[232], x[41], x[40], x[39], x[240], x[239], x[238], x[237], x[62], x[61], x[60], x[258], x[257], x[236], x[235], x[234], x[182], x[181], x[180], x[226], x[225], x[47], x[46], x[45], x[59], x[58], x[57], x[244], x[243], x[256], x[255], x[260], x[259], x[254], x[253], x[229], x[228], x[227], x[179], x[178], x[177], x[44], x[43], x[42], x[50], x[49], x[48], x[116], x[115], x[114], x[252], x[251], x[198], x[197], x[196], x[222], x[221], x[220], x[231], x[230], x[176], x[175], x[174], x[53], x[52], x[51], x[56], x[55], x[54], x[119], x[118], x[117], x[113], x[112], x[111], x[207], x[206], x[205], x[219], x[218], x[217], x[201], x[200], x[199], x[122], x[121], x[120], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[173], x[172], x[171], x[276], x[275], x[89], x[88], x[87], x[389], x[195]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[298], x[297], x[300], x[299], x[302], x[301], x[288], x[287], x[284], x[283], x[276], x[275], x[104], x[103], x[102], x[110], x[109], x[108], x[272], x[271], x[294], x[293], x[282], x[281], x[107], x[106], x[105], x[167], x[166], x[165], x[286], x[285], x[274], x[273], x[280], x[279], x[290], x[289], x[32], x[31], x[30], x[296], x[295], x[89], x[88], x[87], x[292], x[291], x[278], x[277], x[170], x[169], x[168], x[35], x[34], x[33], x[38], x[37], x[36], x[198], x[197], x[196], x[236], x[235], x[234], x[161], x[160], x[159], x[164], x[163], x[162], x[95], x[94], x[93], x[29], x[28], x[27], x[201], x[200], x[199], x[229], x[228], x[227], x[101], x[100], x[99], x[207], x[206], x[205], x[92], x[91], x[90], x[98], x[97], x[96], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[314], x[313], x[219], x[218], x[217], x[86], x[85], x[84], x[390], x[195]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[282], x[281], x[294], x[293], x[38], x[37], x[36], x[302], x[301], x[300], x[299], x[35], x[34], x[33], x[284], x[283], x[290], x[289], x[286], x[285], x[288], x[287], x[298], x[297], x[296], x[295], x[274], x[273], x[292], x[291], x[107], x[106], x[105], x[110], x[109], x[108], x[32], x[31], x[30], x[29], x[28], x[27], x[161], x[160], x[159], x[167], x[166], x[165], x[272], x[271], x[104], x[103], x[102], x[280], x[279], x[276], x[275], x[278], x[277], x[101], x[100], x[99], x[236], x[235], x[234], x[198], x[197], x[196], x[164], x[163], x[162], x[92], x[91], x[90], x[201], x[200], x[199], x[207], x[206], x[205], x[229], x[228], x[227], x[170], x[169], x[168], x[95], x[94], x[93], x[89], x[88], x[87], x[98], x[97], x[96], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[316], x[315], x[219], x[218], x[217], x[83], x[82], x[81], x[391], x[195]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[294], x[293], x[302], x[301], x[296], x[295], x[278], x[277], x[290], x[289], x[284], x[283], x[282], x[281], x[298], x[297], x[300], x[299], x[280], x[279], x[35], x[34], x[33], x[107], x[106], x[105], x[292], x[291], x[274], x[273], x[101], x[100], x[99], x[98], x[97], x[96], x[29], x[28], x[27], x[32], x[31], x[30], x[38], x[37], x[36], x[104], x[103], x[102], x[110], x[109], x[108], x[95], x[94], x[93], x[288], x[287], x[92], x[91], x[90], x[276], x[275], x[164], x[163], x[162], x[272], x[271], x[286], x[285], x[236], x[235], x[234], x[167], x[166], x[165], x[201], x[200], x[199], x[229], x[228], x[227], x[89], x[88], x[87], x[198], x[197], x[196], x[170], x[169], x[168], x[161], x[160], x[159], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[207], x[206], x[205], x[326], x[325], x[219], x[218], x[217], x[80], x[79], x[78], x[392], x[195]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[290], x[289], x[288], x[287], x[272], x[271], x[294], x[293], x[278], x[277], x[274], x[273], x[29], x[28], x[27], x[284], x[283], x[282], x[281], x[280], x[279], x[298], x[297], x[167], x[166], x[165], x[170], x[169], x[168], x[35], x[34], x[33], x[98], x[97], x[96], x[302], x[301], x[296], x[295], x[300], x[299], x[286], x[285], x[164], x[163], x[162], x[32], x[31], x[30], x[38], x[37], x[36], x[95], x[94], x[93], x[276], x[275], x[292], x[291], x[104], x[103], x[102], x[198], x[197], x[196], x[236], x[235], x[234], x[107], x[106], x[105], x[101], x[100], x[99], x[110], x[109], x[108], x[201], x[200], x[199], x[229], x[228], x[227], x[161], x[160], x[159], x[89], x[88], x[87], x[92], x[91], x[90], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[207], x[206], x[205], x[312], x[311], x[219], x[218], x[217], x[77], x[76], x[75], x[393], x[195]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[330], x[329], x[322], x[321], x[328], x[327], x[334], x[333], x[308], x[307], x[338], x[337], x[336], x[335], x[312], x[311], x[332], x[331], x[20], x[19], x[18], x[318], x[317], x[155], x[154], x[153], x[320], x[319], x[310], x[309], x[316], x[315], x[140], x[139], x[138], x[146], x[145], x[144], x[158], x[157], x[156], x[23], x[22], x[21], x[143], x[142], x[141], x[77], x[76], x[75], x[326], x[325], x[314], x[313], x[17], x[16], x[15], x[26], x[25], x[24], x[198], x[197], x[196], x[236], x[235], x[234], x[324], x[323], x[149], x[148], x[147], x[152], x[151], x[150], x[83], x[82], x[81], x[201], x[200], x[199], x[207], x[206], x[205], x[229], x[228], x[227], x[80], x[79], x[78], x[86], x[85], x[84], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[137], x[136], x[135], x[344], x[343], x[219], x[218], x[217], x[74], x[73], x[72], x[394], x[195]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[338], x[337], x[318], x[317], x[23], x[22], x[21], x[26], x[25], x[24], x[330], x[329], x[332], x[331], x[320], x[319], x[322], x[321], x[336], x[335], x[334], x[333], x[20], x[19], x[18], x[17], x[16], x[15], x[310], x[309], x[308], x[307], x[328], x[327], x[326], x[325], x[324], x[323], x[149], x[148], x[147], x[155], x[154], x[153], x[316], x[315], x[312], x[311], x[314], x[313], x[143], x[142], x[141], x[146], x[145], x[144], x[198], x[197], x[196], x[236], x[235], x[234], x[152], x[151], x[150], x[158], x[157], x[156], x[140], x[139], x[138], x[80], x[79], x[78], x[137], x[136], x[135], x[201], x[200], x[199], x[207], x[206], x[205], x[229], x[228], x[227], x[83], x[82], x[81], x[77], x[76], x[75], x[86], x[85], x[84], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[350], x[349], x[219], x[218], x[217], x[71], x[70], x[69], x[395], x[195]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[338], x[337], x[332], x[331], x[330], x[329], x[314], x[313], x[23], x[22], x[21], x[318], x[317], x[336], x[335], x[316], x[315], x[324], x[323], x[17], x[16], x[15], x[20], x[19], x[18], x[328], x[327], x[334], x[333], x[326], x[325], x[310], x[309], x[86], x[85], x[84], x[26], x[25], x[24], x[143], x[142], x[141], x[83], x[82], x[81], x[322], x[321], x[308], x[307], x[137], x[136], x[135], x[140], x[139], x[138], x[146], x[145], x[144], x[80], x[79], x[78], x[312], x[311], x[152], x[151], x[150], x[320], x[319], x[198], x[197], x[196], x[236], x[235], x[234], x[155], x[154], x[153], x[158], x[157], x[156], x[201], x[200], x[199], x[207], x[206], x[205], x[229], x[228], x[227], x[77], x[76], x[75], x[149], x[148], x[147], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[364], x[363], x[219], x[218], x[217], x[68], x[67], x[66], x[396], x[195]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[332], x[331], x[308], x[307], x[338], x[337], x[322], x[321], x[17], x[16], x[15], x[330], x[329], x[314], x[313], x[158], x[157], x[156], x[310], x[309], x[23], x[22], x[21], x[318], x[317], x[316], x[315], x[236], x[235], x[234], x[155], x[154], x[153], x[20], x[19], x[18], x[86], x[85], x[84], x[328], x[327], x[229], x[228], x[227], x[320], x[319], x[152], x[151], x[150], x[26], x[25], x[24], x[83], x[82], x[81], x[312], x[311], x[326], x[325], x[336], x[335], x[324], x[323], x[334], x[333], x[198], x[197], x[196], x[222], x[221], x[220], x[140], x[139], x[138], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[149], x[148], x[147], x[77], x[76], x[75], x[80], x[79], x[78], x[143], x[142], x[141], x[137], x[136], x[135], x[146], x[145], x[144], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[346], x[345], x[65], x[64], x[63], x[397], x[195]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[356], x[355], x[346], x[345], x[352], x[351], x[360], x[359], x[366], x[365], x[354], x[353], x[362], x[361], x[263], x[262], x[350], x[349], x[358], x[357], x[216], x[215], x[8], x[7], x[6], x[65], x[64], x[63], x[364], x[363], x[128], x[127], x[126], x[134], x[133], x[132], x[11], x[10], x[9], x[14], x[13], x[12], x[131], x[130], x[129], x[191], x[190], x[189], x[269], x[268], x[266], x[265], x[71], x[70], x[69], x[344], x[343], x[5], x[4], x[3], x[194], x[193], x[192], x[236], x[235], x[234], x[348], x[347], x[198], x[197], x[196], x[68], x[67], x[66], x[201], x[200], x[199], x[207], x[206], x[205], x[229], x[228], x[227], x[185], x[184], x[183], x[188], x[187], x[186], x[74], x[73], x[72], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[125], x[124], x[123], x[246], x[245], x[219], x[218], x[217], x[62], x[61], x[60], x[398], x[195]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[354], x[353], x[366], x[365], x[14], x[13], x[12], x[11], x[10], x[9], x[356], x[355], x[358], x[357], x[364], x[363], x[362], x[361], x[360], x[359], x[8], x[7], x[6], x[5], x[4], x[3], x[269], x[268], x[263], x[262], x[352], x[351], x[350], x[349], x[346], x[345], x[348], x[347], x[266], x[265], x[216], x[215], x[68], x[67], x[66], x[344], x[343], x[131], x[130], x[129], x[134], x[133], x[132], x[185], x[184], x[183], x[236], x[235], x[234], x[191], x[190], x[189], x[128], x[127], x[126], x[71], x[70], x[69], x[65], x[64], x[63], x[125], x[124], x[123], x[201], x[200], x[199], x[229], x[228], x[227], x[188], x[187], x[186], x[194], x[193], x[192], x[198], x[197], x[196], x[207], x[206], x[205], x[74], x[73], x[72], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[248], x[247], x[219], x[218], x[217], x[59], x[58], x[57], x[399], x[195]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[366], x[365], x[358], x[357], x[356], x[355], x[354], x[353], x[350], x[349], x[344], x[343], x[11], x[10], x[9], x[362], x[361], x[364], x[363], x[348], x[347], x[5], x[4], x[3], x[8], x[7], x[6], x[14], x[13], x[12], x[352], x[351], x[360], x[359], x[71], x[70], x[69], x[74], x[73], x[72], x[131], x[130], x[129], x[68], x[67], x[66], x[346], x[345], x[266], x[265], x[125], x[124], x[123], x[128], x[127], x[126], x[134], x[133], x[132], x[263], x[262], x[216], x[215], x[198], x[197], x[196], x[236], x[235], x[234], x[65], x[64], x[63], x[188], x[187], x[186], x[269], x[268], x[201], x[200], x[199], x[229], x[228], x[227], x[207], x[206], x[205], x[191], x[190], x[189], x[194], x[193], x[192], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[185], x[184], x[183], x[256], x[255], x[219], x[218], x[217], x[56], x[55], x[54], x[400], x[195]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[358], x[357], x[366], x[365], x[216], x[215], x[5], x[4], x[3], x[356], x[355], x[354], x[353], x[350], x[349], x[344], x[343], x[263], x[262], x[11], x[10], x[9], x[194], x[193], x[192], x[266], x[265], x[8], x[7], x[6], x[14], x[13], x[12], x[71], x[70], x[69], x[74], x[73], x[72], x[346], x[345], x[364], x[363], x[352], x[351], x[191], x[190], x[189], x[362], x[361], x[348], x[347], x[360], x[359], x[198], x[197], x[196], x[236], x[235], x[234], x[269], x[268], x[188], x[187], x[186], x[65], x[64], x[63], x[68], x[67], x[66], x[128], x[127], x[126], x[201], x[200], x[199], x[229], x[228], x[227], x[207], x[206], x[205], x[131], x[130], x[129], x[125], x[124], x[123], x[134], x[133], x[132], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[185], x[184], x[183], x[244], x[243], x[219], x[218], x[217], x[53], x[52], x[51], x[401], x[195]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[256], x[255], x[246], x[245], x[248], x[247], x[260], x[259], x[252], x[251], x[56], x[55], x[54], x[62], x[61], x[60], x[224], x[223], x[242], x[241], x[59], x[58], x[57], x[119], x[118], x[117], x[122], x[121], x[120], x[254], x[253], x[258], x[257], x[236], x[235], x[234], x[233], x[232], x[250], x[249], x[244], x[243], x[229], x[228], x[227], x[182], x[181], x[180], x[41], x[40], x[39], x[240], x[239], x[113], x[112], x[111], x[116], x[115], x[114], x[198], x[197], x[196], x[222], x[221], x[220], x[179], x[178], x[177], x[231], x[230], x[226], x[225], x[47], x[46], x[45], x[53], x[52], x[51], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[44], x[43], x[42], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[173], x[172], x[171], x[176], x[175], x[174], x[238], x[237], x[50], x[49], x[48], x[402], x[195]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[246], x[245], x[254], x[253], x[248], x[247], x[260], x[259], x[62], x[61], x[60], x[113], x[112], x[111], x[258], x[257], x[59], x[58], x[57], x[244], x[243], x[256], x[255], x[231], x[230], x[236], x[235], x[234], x[119], x[118], x[117], x[252], x[251], x[233], x[232], x[240], x[239], x[229], x[228], x[227], x[116], x[115], x[114], x[53], x[52], x[51], x[56], x[55], x[54], x[173], x[172], x[171], x[226], x[225], x[224], x[223], x[238], x[237], x[198], x[197], x[196], x[222], x[221], x[220], x[242], x[241], x[122], x[121], x[120], x[179], x[178], x[177], x[44], x[43], x[42], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[176], x[175], x[174], x[182], x[181], x[180], x[50], x[49], x[48], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[41], x[40], x[39], x[250], x[249], x[47], x[46], x[45], x[403], x[195]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[244], x[243], x[238], x[237], x[248], x[247], x[250], x[249], x[53], x[52], x[51], x[256], x[255], x[246], x[245], x[258], x[257], x[50], x[49], x[48], x[59], x[58], x[57], x[226], x[225], x[236], x[235], x[234], x[260], x[259], x[47], x[46], x[45], x[242], x[241], x[56], x[55], x[54], x[62], x[61], x[60], x[233], x[232], x[224], x[223], x[229], x[228], x[227], x[254], x[253], x[116], x[115], x[114], x[252], x[251], x[176], x[175], x[174], x[231], x[230], x[198], x[197], x[196], x[222], x[221], x[220], x[119], x[118], x[117], x[41], x[40], x[39], x[179], x[178], x[177], x[182], x[181], x[180], x[207], x[206], x[205], x[219], x[218], x[217], x[113], x[112], x[111], x[122], x[121], x[120], x[173], x[172], x[171], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[201], x[200], x[199], x[240], x[239], x[44], x[43], x[42], x[404], x[195]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[258], x[257], x[260], x[259], x[252], x[251], x[226], x[225], x[224], x[223], x[238], x[237], x[116], x[115], x[114], x[233], x[232], x[256], x[255], x[250], x[249], x[236], x[235], x[234], x[119], x[118], x[117], x[122], x[121], x[120], x[176], x[175], x[174], x[182], x[181], x[180], x[248], x[247], x[244], x[243], x[246], x[245], x[50], x[49], x[48], x[229], x[228], x[227], x[254], x[253], x[179], x[178], x[177], x[56], x[55], x[54], x[47], x[46], x[45], x[240], x[239], x[198], x[197], x[196], x[222], x[221], x[220], x[231], x[230], x[59], x[58], x[57], x[53], x[52], x[51], x[62], x[61], x[60], x[207], x[206], x[205], x[219], x[218], x[217], x[113], x[112], x[111], x[44], x[43], x[42], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[201], x[200], x[199], x[173], x[172], x[171], x[242], x[241], x[41], x[40], x[39], x[405], x[195]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[300], x[299], x[292], x[291], x[278], x[277], x[302], x[301], x[280], x[279], x[110], x[109], x[108], x[288], x[287], x[272], x[271], x[290], x[289], x[92], x[91], x[90], x[98], x[97], x[96], x[107], x[106], x[105], x[296], x[295], x[298], x[297], x[236], x[235], x[234], x[294], x[293], x[95], x[94], x[93], x[229], x[228], x[227], x[167], x[166], x[165], x[170], x[169], x[168], x[286], x[285], x[274], x[273], x[29], x[28], x[27], x[284], x[283], x[276], x[275], x[101], x[100], x[99], x[104], x[103], x[102], x[222], x[221], x[220], x[198], x[197], x[196], x[35], x[34], x[33], x[201], x[200], x[199], x[219], x[218], x[217], x[161], x[160], x[159], x[164], x[163], x[162], x[32], x[31], x[30], x[89], x[88], x[87], x[204], x[203], x[202], x[210], x[209], x[208], x[207], x[206], x[205], x[213], x[212], x[211], x[282], x[281], x[38], x[37], x[36], x[406], x[195]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[296], x[295], x[278], x[277], x[302], x[301], x[280], x[279], x[286], x[285], x[101], x[100], x[99], x[298], x[297], x[300], x[299], x[98], x[97], x[96], x[288], x[287], x[236], x[235], x[234], x[107], x[106], x[105], x[95], x[94], x[93], x[276], x[275], x[292], x[291], x[161], x[160], x[159], x[274], x[273], x[284], x[283], x[229], x[228], x[227], x[104], x[103], x[102], x[110], x[109], x[108], x[167], x[166], x[165], x[272], x[271], x[282], x[281], x[222], x[221], x[220], x[290], x[289], x[89], x[88], x[87], x[92], x[91], x[90], x[198], x[197], x[196], x[164], x[163], x[162], x[32], x[31], x[30], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[170], x[169], x[168], x[38], x[37], x[36], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[29], x[28], x[27], x[294], x[293], x[35], x[34], x[33], x[407], x[195]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[282], x[281], x[276], x[275], x[294], x[293], x[280], x[279], x[274], x[273], x[298], x[297], x[38], x[37], x[36], x[89], x[88], x[87], x[292], x[291], x[278], x[277], x[288], x[287], x[236], x[235], x[234], x[302], x[301], x[300], x[299], x[35], x[34], x[33], x[290], x[289], x[95], x[94], x[93], x[164], x[163], x[162], x[272], x[271], x[286], x[285], x[229], x[228], x[227], x[296], x[295], x[104], x[103], x[102], x[92], x[91], x[90], x[98], x[97], x[96], x[167], x[166], x[165], x[222], x[221], x[220], x[107], x[106], x[105], x[110], x[109], x[108], x[29], x[28], x[27], x[198], x[197], x[196], x[170], x[169], x[168], x[161], x[160], x[159], x[201], x[200], x[199], x[219], x[218], x[217], x[101], x[100], x[99], x[207], x[206], x[205], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[284], x[283], x[32], x[31], x[30], x[408], x[195]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[298], x[297], x[300], x[299], x[274], x[273], x[302], x[301], x[288], x[287], x[272], x[271], x[282], x[281], x[104], x[103], x[102], x[110], x[109], x[108], x[164], x[163], x[162], x[294], x[293], x[236], x[235], x[234], x[107], x[106], x[105], x[167], x[166], x[165], x[170], x[169], x[168], x[292], x[291], x[38], x[37], x[36], x[229], x[228], x[227], x[296], x[295], x[286], x[285], x[280], x[279], x[276], x[275], x[278], x[277], x[35], x[34], x[33], x[284], x[283], x[198], x[197], x[196], x[222], x[221], x[220], x[92], x[91], x[90], x[201], x[200], x[199], x[219], x[218], x[217], x[101], x[100], x[99], x[161], x[160], x[159], x[95], x[94], x[93], x[89], x[88], x[87], x[98], x[97], x[96], x[32], x[31], x[30], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[207], x[206], x[205], x[290], x[289], x[29], x[28], x[27], x[409], x[195]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[326], x[325], x[314], x[313], x[334], x[333], x[308], x[307], x[332], x[331], x[316], x[315], x[336], x[335], x[322], x[321], x[338], x[337], x[80], x[79], x[78], x[86], x[85], x[84], x[146], x[145], x[144], x[236], x[235], x[234], x[158], x[157], x[156], x[17], x[16], x[15], x[330], x[329], x[83], x[82], x[81], x[143], x[142], x[141], x[324], x[323], x[328], x[327], x[229], x[228], x[227], x[155], x[154], x[153], x[320], x[319], x[310], x[309], x[23], x[22], x[21], x[312], x[311], x[198], x[197], x[196], x[222], x[221], x[220], x[20], x[19], x[18], x[137], x[136], x[135], x[140], x[139], x[138], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[149], x[148], x[147], x[152], x[151], x[150], x[77], x[76], x[75], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[318], x[317], x[26], x[25], x[24], x[410], x[195]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[314], x[313], x[324], x[323], x[316], x[315], x[320], x[319], x[336], x[335], x[86], x[85], x[84], x[322], x[321], x[330], x[329], x[236], x[235], x[234], x[137], x[136], x[135], x[328], x[327], x[334], x[333], x[83], x[82], x[81], x[312], x[311], x[326], x[325], x[149], x[148], x[147], x[310], x[309], x[308], x[307], x[229], x[228], x[227], x[332], x[331], x[143], x[142], x[141], x[155], x[154], x[153], x[20], x[19], x[18], x[318], x[317], x[198], x[197], x[196], x[222], x[221], x[220], x[140], x[139], x[138], x[146], x[145], x[144], x[77], x[76], x[75], x[80], x[79], x[78], x[152], x[151], x[150], x[158], x[157], x[156], x[207], x[206], x[205], x[219], x[218], x[217], x[17], x[16], x[15], x[26], x[25], x[24], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[201], x[200], x[199], x[338], x[337], x[23], x[22], x[21], x[411], x[195]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[338], x[337], x[318], x[317], x[312], x[311], x[316], x[315], x[310], x[309], x[23], x[22], x[21], x[26], x[25], x[24], x[332], x[331], x[77], x[76], x[75], x[326], x[325], x[314], x[313], x[322], x[321], x[308], x[307], x[236], x[235], x[234], x[328], x[327], x[83], x[82], x[81], x[152], x[151], x[150], x[320], x[319], x[229], x[228], x[227], x[336], x[335], x[334], x[333], x[17], x[16], x[15], x[80], x[79], x[78], x[86], x[85], x[84], x[155], x[154], x[153], x[158], x[157], x[156], x[198], x[197], x[196], x[222], x[221], x[220], x[324], x[323], x[140], x[139], x[138], x[149], x[148], x[147], x[201], x[200], x[199], x[207], x[206], x[205], x[219], x[218], x[217], x[143], x[142], x[141], x[146], x[145], x[144], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[137], x[136], x[135], x[330], x[329], x[20], x[19], x[18], x[412], x[195]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[310], x[309], x[308], x[307], x[328], x[327], x[334], x[333], x[322], x[321], x[338], x[337], x[318], x[317], x[336], x[335], x[152], x[151], x[150], x[158], x[157], x[156], x[236], x[235], x[234], x[140], x[139], x[138], x[146], x[145], x[144], x[155], x[154], x[153], x[326], x[325], x[23], x[22], x[21], x[26], x[25], x[24], x[330], x[329], x[229], x[228], x[227], x[143], x[142], x[141], x[320], x[319], x[316], x[315], x[312], x[311], x[314], x[313], x[198], x[197], x[196], x[222], x[221], x[220], x[324], x[323], x[80], x[79], x[78], x[20], x[19], x[18], x[207], x[206], x[205], x[219], x[218], x[217], x[149], x[148], x[147], x[83], x[82], x[81], x[77], x[76], x[75], x[86], x[85], x[84], x[201], x[200], x[199], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[137], x[136], x[135], x[332], x[331], x[17], x[16], x[15], x[413], x[195]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[364], x[363], x[350], x[349], x[344], x[343], x[360], x[359], x[358], x[357], x[68], x[67], x[66], x[362], x[361], x[216], x[215], x[366], x[365], x[71], x[70], x[69], x[74], x[73], x[72], x[134], x[133], x[132], x[263], x[262], x[5], x[4], x[3], x[356], x[355], x[346], x[345], x[131], x[130], x[129], x[348], x[347], x[352], x[351], x[194], x[193], x[192], x[11], x[10], x[9], x[198], x[197], x[196], x[236], x[235], x[234], x[191], x[190], x[189], x[269], x[268], x[266], x[265], x[8], x[7], x[6], x[65], x[64], x[63], x[125], x[124], x[123], x[128], x[127], x[126], x[201], x[200], x[199], x[229], x[228], x[227], x[207], x[206], x[205], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[185], x[184], x[183], x[188], x[187], x[186], x[354], x[353], x[219], x[218], x[217], x[14], x[13], x[12], x[414], x[195]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[350], x[349], x[344], x[343], x[348], x[347], x[362], x[361], x[71], x[70], x[69], x[74], x[73], x[72], x[346], x[345], x[364], x[363], x[269], x[268], x[356], x[355], x[125], x[124], x[123], x[352], x[351], x[360], x[359], x[263], x[262], x[354], x[353], x[358], x[357], x[131], x[130], x[129], x[65], x[64], x[63], x[68], x[67], x[66], x[185], x[184], x[183], x[266], x[265], x[216], x[215], x[8], x[7], x[6], x[198], x[197], x[196], x[236], x[235], x[234], x[128], x[127], x[126], x[134], x[133], x[132], x[191], x[190], x[189], x[14], x[13], x[12], x[201], x[200], x[199], x[207], x[206], x[205], x[229], x[228], x[227], x[5], x[4], x[3], x[188], x[187], x[186], x[194], x[193], x[192], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[366], x[365], x[219], x[218], x[217], x[11], x[10], x[9], x[415], x[195]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[354], x[353], x[346], x[345], x[366], x[365], x[350], x[349], x[14], x[13], x[12], x[65], x[64], x[63], x[364], x[363], x[11], x[10], x[9], x[358], x[357], x[71], x[70], x[69], x[344], x[343], x[266], x[265], x[352], x[351], x[68], x[67], x[66], x[263], x[262], x[216], x[215], x[362], x[361], x[360], x[359], x[5], x[4], x[3], x[74], x[73], x[72], x[188], x[187], x[186], x[269], x[268], x[198], x[197], x[196], x[236], x[235], x[234], x[348], x[347], x[128], x[127], x[126], x[191], x[190], x[189], x[194], x[193], x[192], x[201], x[200], x[199], x[207], x[206], x[205], x[229], x[228], x[227], x[131], x[130], x[129], x[134], x[133], x[132], x[185], x[184], x[183], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[125], x[124], x[123], x[356], x[355], x[219], x[218], x[217], x[8], x[7], x[6], x[416], x[195]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[354], x[353], x[352], x[351], x[360], x[359], x[266], x[265], x[216], x[215], x[366], x[365], x[362], x[361], x[263], x[262], x[364], x[363], x[14], x[13], x[12], x[128], x[127], x[126], x[134], x[133], x[132], x[188], x[187], x[186], x[194], x[193], x[192], x[350], x[349], x[346], x[345], x[11], x[10], x[9], x[356], x[355], x[131], x[130], x[129], x[191], x[190], x[189], x[68], x[67], x[66], x[344], x[343], x[236], x[235], x[234], x[348], x[347], x[269], x[268], x[71], x[70], x[69], x[65], x[64], x[63], x[8], x[7], x[6], x[201], x[200], x[199], x[229], x[228], x[227], x[198], x[197], x[196], x[207], x[206], x[205], x[74], x[73], x[72], x[213], x[212], x[211], x[204], x[203], x[202], x[210], x[209], x[208], x[222], x[221], x[220], x[125], x[124], x[123], x[185], x[184], x[183], x[358], x[357], x[219], x[218], x[217], x[5], x[4], x[3], x[417], x[195]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[210], x[209], x[208], x[195]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[201], x[200], x[199], x[195]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[198], x[197], x[196], x[195]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[213], x[212], x[211], x[195]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[207], x[206], x[205], x[195]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[204], x[203], x[202], x[210], x[209], x[208], x[195]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[222], x[221], x[220], x[195]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[229], x[228], x[227], x[195]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[236], x[235], x[234], x[195]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[195], x[219], x[218], x[217]}), .y(y[139]));
endmodule

module R2ind0(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (t[2] & ~t[3]);
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[1];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [21:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = t[21] ^ x[3];
  assign t[15] = t[22] ^ x[6];
  assign t[16] = t[23] ^ x[9];
  assign t[17] = t[24] ^ x[12];
  assign t[18] = t[25] ^ x[15];
  assign t[19] = t[26] ^ x[18];
  assign t[1] = ~(t[7] | t[2]);
  assign t[20] = t[27] ^ x[21];
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = (t[34] & ~t[35]);
  assign t[25] = (t[36] & ~t[37]);
  assign t[26] = (t[38] & ~t[39]);
  assign t[27] = (t[40] & ~t[41]);
  assign t[28] = t[42] ^ x[3];
  assign t[29] = t[43] ^ x[2];
  assign t[2] = ~(t[8] | t[3]);
  assign t[30] = t[44] ^ x[6];
  assign t[31] = t[45] ^ x[5];
  assign t[32] = t[46] ^ x[9];
  assign t[33] = t[47] ^ x[8];
  assign t[34] = t[48] ^ x[12];
  assign t[35] = t[49] ^ x[11];
  assign t[36] = t[50] ^ x[15];
  assign t[37] = t[51] ^ x[14];
  assign t[38] = t[52] ^ x[18];
  assign t[39] = t[53] ^ x[17];
  assign t[3] = ~(t[9] & t[4]);
  assign t[40] = t[54] ^ x[21];
  assign t[41] = t[55] ^ x[20];
  assign t[42] = (x[1]);
  assign t[43] = (x[1]);
  assign t[44] = (x[4]);
  assign t[45] = (x[4]);
  assign t[46] = (x[7]);
  assign t[47] = (x[7]);
  assign t[48] = (x[10]);
  assign t[49] = (x[10]);
  assign t[4] = ~(t[10] | t[5]);
  assign t[50] = (x[13]);
  assign t[51] = (x[13]);
  assign t[52] = (x[16]);
  assign t[53] = (x[16]);
  assign t[54] = (x[19]);
  assign t[55] = (x[19]);
  assign t[5] = ~(t[11] & t[6]);
  assign t[6] = ~(t[12] | t[13]);
  assign t[7] = (t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind3(x, y);
 input [21:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = t[21] ^ x[3];
  assign t[15] = t[22] ^ x[6];
  assign t[16] = t[23] ^ x[9];
  assign t[17] = t[24] ^ x[12];
  assign t[18] = t[25] ^ x[15];
  assign t[19] = t[26] ^ x[18];
  assign t[1] = ~(t[7] | t[2]);
  assign t[20] = t[27] ^ x[21];
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = (t[34] & ~t[35]);
  assign t[25] = (t[36] & ~t[37]);
  assign t[26] = (t[38] & ~t[39]);
  assign t[27] = (t[40] & ~t[41]);
  assign t[28] = t[42] ^ x[3];
  assign t[29] = t[43] ^ x[2];
  assign t[2] = ~(t[8] | t[3]);
  assign t[30] = t[44] ^ x[6];
  assign t[31] = t[45] ^ x[5];
  assign t[32] = t[46] ^ x[9];
  assign t[33] = t[47] ^ x[8];
  assign t[34] = t[48] ^ x[12];
  assign t[35] = t[49] ^ x[11];
  assign t[36] = t[50] ^ x[15];
  assign t[37] = t[51] ^ x[14];
  assign t[38] = t[52] ^ x[18];
  assign t[39] = t[53] ^ x[17];
  assign t[3] = ~(t[9] & t[4]);
  assign t[40] = t[54] ^ x[21];
  assign t[41] = t[55] ^ x[20];
  assign t[42] = (x[1]);
  assign t[43] = (x[1]);
  assign t[44] = (x[4]);
  assign t[45] = (x[4]);
  assign t[46] = (x[7]);
  assign t[47] = (x[7]);
  assign t[48] = (x[10]);
  assign t[49] = (x[10]);
  assign t[4] = ~(t[10] | t[5]);
  assign t[50] = (x[13]);
  assign t[51] = (x[13]);
  assign t[52] = (x[16]);
  assign t[53] = (x[16]);
  assign t[54] = (x[19]);
  assign t[55] = (x[19]);
  assign t[5] = ~(t[11] & t[6]);
  assign t[6] = ~(t[12] | t[13]);
  assign t[7] = (t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind4(x, y);
 input [6:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = x[0] | t[1];
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[2];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[5];
  assign t[14] = (x[1]);
  assign t[15] = (x[1]);
  assign t[16] = (x[4]);
  assign t[17] = (x[4]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[3];
  assign t[7] = t[9] ^ x[6];
  assign t[8] = (t[10] & ~t[11]);
  assign t[9] = (t[12] & ~t[13]);
  assign y = (t[0]);
endmodule

module R2ind5(x, y);
 input [6:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = x[0] | t[1];
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[2];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[5];
  assign t[14] = (x[1]);
  assign t[15] = (x[1]);
  assign t[16] = (x[4]);
  assign t[17] = (x[4]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[3];
  assign t[7] = t[9] ^ x[6];
  assign t[8] = (t[10] & ~t[11]);
  assign t[9] = (t[12] & ~t[13]);
  assign y = (t[0]);
endmodule

module R2ind6(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind7(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind8(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind9(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind11(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind12(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind13(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind14(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1] | x[0]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1] | x[0]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind16(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1] | x[3]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind17(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1] | x[3]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind18(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1] | x[0]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind19(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1] | x[0]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1] | x[0]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind21(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1] | x[0]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind22(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1] | x[0]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind23(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1] | x[0]);
  assign t[1] = ~(t[2]);
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind24(x, y);
 input [111:0] x;
 output y;

 wire [323:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[118] ^ t[119];
  assign t[101] = t[119] ^ t[24];
  assign t[102] = ~(t[116]);
  assign t[103] = ~(t[121]);
  assign t[104] = ~(t[122]);
  assign t[105] = ~(t[123]);
  assign t[106] = t[44] ? t[124] : t[161];
  assign t[107] = t[122] ^ t[123];
  assign t[108] = t[123] ^ t[26];
  assign t[109] = ~(t[143]);
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[125] ? x[71] : x[70];
  assign t[111] = ~t[126];
  assign t[112] = t[8] ? t[127] : t[162];
  assign t[113] = t[125] ? x[76] : x[75];
  assign t[114] = t[159] ^ t[128];
  assign t[115] = t[31] ? x[78] : x[77];
  assign t[116] = ~(t[31]);
  assign t[117] = t[99] ^ t[119];
  assign t[118] = t[44] ? t[129] : t[163];
  assign t[119] = t[44] ? t[130] : t[164];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[160] ^ t[131];
  assign t[121] = t[106] ^ t[123];
  assign t[122] = t[44] ? t[132] : t[165];
  assign t[123] = t[44] ? t[133] : t[166];
  assign t[124] = t[161] ^ t[134];
  assign t[125] = ~(t[116]);
  assign t[126] = t[8] ? t[135] : t[167];
  assign t[127] = t[162] ^ t[136];
  assign t[128] = t[95] ? x[95] : x[94];
  assign t[129] = t[163] ^ t[137];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[164] ^ t[138];
  assign t[131] = t[95] ? x[97] : x[96];
  assign t[132] = t[165] ^ t[139];
  assign t[133] = t[166] ^ t[140];
  assign t[134] = t[102] ? x[99] : x[98];
  assign t[135] = t[167] ^ t[141];
  assign t[136] = t[125] ? x[101] : x[100];
  assign t[137] = t[95] ? x[103] : x[102];
  assign t[138] = t[95] ? x[105] : x[104];
  assign t[139] = t[102] ? x[107] : x[106];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[102] ? x[109] : x[108];
  assign t[141] = t[31] ? x[111] : x[110];
  assign t[142] = (t[168]);
  assign t[143] = (t[169]);
  assign t[144] = (t[170]);
  assign t[145] = (t[171]);
  assign t[146] = (t[172]);
  assign t[147] = (t[173]);
  assign t[148] = (t[174]);
  assign t[149] = (t[175]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = (t[176]);
  assign t[151] = (t[177]);
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = t[194] ^ x[4];
  assign t[169] = t[195] ^ x[7];
  assign t[16] = t[143] | t[30];
  assign t[170] = t[196] ^ x[12];
  assign t[171] = t[197] ^ x[15];
  assign t[172] = t[198] ^ x[18];
  assign t[173] = t[199] ^ x[21];
  assign t[174] = t[200] ^ x[24];
  assign t[175] = t[201] ^ x[27];
  assign t[176] = t[202] ^ x[30];
  assign t[177] = t[203] ^ x[33];
  assign t[178] = t[204] ^ x[36];
  assign t[179] = t[205] ^ x[39];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[206] ^ x[42];
  assign t[181] = t[207] ^ x[45];
  assign t[182] = t[208] ^ x[48];
  assign t[183] = t[209] ^ x[51];
  assign t[184] = t[210] ^ x[58];
  assign t[185] = t[211] ^ x[63];
  assign t[186] = t[212] ^ x[66];
  assign t[187] = t[213] ^ x[69];
  assign t[188] = t[214] ^ x[74];
  assign t[189] = t[215] ^ x[81];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[216] ^ x[84];
  assign t[191] = t[217] ^ x[87];
  assign t[192] = t[218] ^ x[90];
  assign t[193] = t[219] ^ x[93];
  assign t[194] = (t[220] & ~t[221]);
  assign t[195] = (t[222] & ~t[223]);
  assign t[196] = (t[224] & ~t[225]);
  assign t[197] = (t[226] & ~t[227]);
  assign t[198] = (t[228] & ~t[229]);
  assign t[199] = (t[230] & ~t[231]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[232] & ~t[233]);
  assign t[201] = (t[234] & ~t[235]);
  assign t[202] = (t[236] & ~t[237]);
  assign t[203] = (t[238] & ~t[239]);
  assign t[204] = (t[240] & ~t[241]);
  assign t[205] = (t[242] & ~t[243]);
  assign t[206] = (t[244] & ~t[245]);
  assign t[207] = (t[246] & ~t[247]);
  assign t[208] = (t[248] & ~t[249]);
  assign t[209] = (t[250] & ~t[251]);
  assign t[20] = t[36] ^ t[37];
  assign t[210] = (t[252] & ~t[253]);
  assign t[211] = (t[254] & ~t[255]);
  assign t[212] = (t[256] & ~t[257]);
  assign t[213] = (t[258] & ~t[259]);
  assign t[214] = (t[260] & ~t[261]);
  assign t[215] = (t[262] & ~t[263]);
  assign t[216] = (t[264] & ~t[265]);
  assign t[217] = (t[266] & ~t[267]);
  assign t[218] = (t[268] & ~t[269]);
  assign t[219] = (t[270] & ~t[271]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[272] ^ x[4];
  assign t[221] = t[273] ^ x[3];
  assign t[222] = t[274] ^ x[7];
  assign t[223] = t[275] ^ x[6];
  assign t[224] = t[276] ^ x[12];
  assign t[225] = t[277] ^ x[11];
  assign t[226] = t[278] ^ x[15];
  assign t[227] = t[279] ^ x[14];
  assign t[228] = t[280] ^ x[18];
  assign t[229] = t[281] ^ x[17];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[282] ^ x[21];
  assign t[231] = t[283] ^ x[20];
  assign t[232] = t[284] ^ x[24];
  assign t[233] = t[285] ^ x[23];
  assign t[234] = t[286] ^ x[27];
  assign t[235] = t[287] ^ x[26];
  assign t[236] = t[288] ^ x[30];
  assign t[237] = t[289] ^ x[29];
  assign t[238] = t[290] ^ x[33];
  assign t[239] = t[291] ^ x[32];
  assign t[23] = t[42] & t[43];
  assign t[240] = t[292] ^ x[36];
  assign t[241] = t[293] ^ x[35];
  assign t[242] = t[294] ^ x[39];
  assign t[243] = t[295] ^ x[38];
  assign t[244] = t[296] ^ x[42];
  assign t[245] = t[297] ^ x[41];
  assign t[246] = t[298] ^ x[45];
  assign t[247] = t[299] ^ x[44];
  assign t[248] = t[300] ^ x[48];
  assign t[249] = t[301] ^ x[47];
  assign t[24] = t[44] ? t[45] : t[144];
  assign t[250] = t[302] ^ x[51];
  assign t[251] = t[303] ^ x[50];
  assign t[252] = t[304] ^ x[58];
  assign t[253] = t[305] ^ x[57];
  assign t[254] = t[306] ^ x[63];
  assign t[255] = t[307] ^ x[62];
  assign t[256] = t[308] ^ x[66];
  assign t[257] = t[309] ^ x[65];
  assign t[258] = t[310] ^ x[69];
  assign t[259] = t[311] ^ x[68];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[312] ^ x[74];
  assign t[261] = t[313] ^ x[73];
  assign t[262] = t[314] ^ x[81];
  assign t[263] = t[315] ^ x[80];
  assign t[264] = t[316] ^ x[84];
  assign t[265] = t[317] ^ x[83];
  assign t[266] = t[318] ^ x[87];
  assign t[267] = t[319] ^ x[86];
  assign t[268] = t[320] ^ x[90];
  assign t[269] = t[321] ^ x[89];
  assign t[26] = t[44] ? t[48] : t[145];
  assign t[270] = t[322] ^ x[93];
  assign t[271] = t[323] ^ x[92];
  assign t[272] = (x[2]);
  assign t[273] = (x[2]);
  assign t[274] = (x[5]);
  assign t[275] = (x[5]);
  assign t[276] = (x[10]);
  assign t[277] = (x[10]);
  assign t[278] = (x[13]);
  assign t[279] = (x[13]);
  assign t[27] = t[49] ^ t[50];
  assign t[280] = (x[16]);
  assign t[281] = (x[16]);
  assign t[282] = (x[19]);
  assign t[283] = (x[19]);
  assign t[284] = (x[22]);
  assign t[285] = (x[22]);
  assign t[286] = (x[25]);
  assign t[287] = (x[25]);
  assign t[288] = (x[28]);
  assign t[289] = (x[28]);
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = (x[31]);
  assign t[291] = (x[31]);
  assign t[292] = (x[34]);
  assign t[293] = (x[34]);
  assign t[294] = (x[37]);
  assign t[295] = (x[37]);
  assign t[296] = (x[40]);
  assign t[297] = (x[40]);
  assign t[298] = (x[43]);
  assign t[299] = (x[43]);
  assign t[29] = ~(t[146] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[46]);
  assign t[301] = (x[46]);
  assign t[302] = (x[49]);
  assign t[303] = (x[49]);
  assign t[304] = (x[56]);
  assign t[305] = (x[56]);
  assign t[306] = (x[61]);
  assign t[307] = (x[61]);
  assign t[308] = (x[64]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = (x[67]);
  assign t[311] = (x[67]);
  assign t[312] = (x[72]);
  assign t[313] = (x[72]);
  assign t[314] = (x[79]);
  assign t[315] = (x[79]);
  assign t[316] = (x[82]);
  assign t[317] = (x[82]);
  assign t[318] = (x[85]);
  assign t[319] = (x[85]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[88]);
  assign t[321] = (x[88]);
  assign t[322] = (x[91]);
  assign t[323] = (x[91]);
  assign t[32] = ~(t[147]);
  assign t[33] = ~(t[148]);
  assign t[34] = ~(t[149]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = t[57];
  assign t[37] = t[4];
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[60] & t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[62] : t[150];
  assign t[41] = t[151] ^ t[63];
  assign t[42] = ~(t[64]);
  assign t[43] = t[152] ^ t[65];
  assign t[44] = ~(t[66]);
  assign t[45] = t[144] ^ t[67];
  assign t[46] = t[68] ^ t[69];
  assign t[47] = t[70] & t[71];
  assign t[48] = t[145] ^ t[72];
  assign t[49] = t[73] ^ t[74];
  assign t[4] = t[8] ? t[9] : t[142];
  assign t[50] = t[75] & t[76];
  assign t[51] = ~(t[77] & t[78]);
  assign t[52] = t[79] ^ t[153];
  assign t[53] = ~(t[146]);
  assign t[54] = t[80] & t[79];
  assign t[55] = ~(t[151]);
  assign t[56] = ~(t[81] & t[154]);
  assign t[57] = t[8] ? t[82] : t[155];
  assign t[58] = t[83] & t[84];
  assign t[59] = t[85] & t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = ~(t[58] ^ t[87]);
  assign t[61] = t[88] ^ t[89];
  assign t[62] = t[150] ^ t[90];
  assign t[63] = t[91] ? t[92] : t[156];
  assign t[64] = t[149] ^ t[93];
  assign t[65] = t[8] ? t[94] : t[157];
  assign t[66] = ~(t[8]);
  assign t[67] = t[95] ? x[53] : x[52];
  assign t[68] = t[96] & t[97];
  assign t[69] = t[98] & t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[100] ^ t[46]);
  assign t[71] = t[101] ^ t[99];
  assign t[72] = t[102] ? x[55] : x[54];
  assign t[73] = t[103] & t[104];
  assign t[74] = t[105] & t[106];
  assign t[75] = ~(t[107] ^ t[49]);
  assign t[76] = t[108] ^ t[106];
  assign t[77] = ~(t[80] | t[79]);
  assign t[78] = ~(t[109] | t[53]);
  assign t[79] = ~(t[158]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[153]);
  assign t[81] = ~(t[152]);
  assign t[82] = t[155] ^ t[110];
  assign t[83] = ~(t[89]);
  assign t[84] = ~(t[111]);
  assign t[85] = ~(t[36]);
  assign t[86] = t[112];
  assign t[87] = t[20] ^ t[111];
  assign t[88] = t[111] ^ t[37];
  assign t[89] = t[86] ^ t[36];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[95] ? x[60] : x[59];
  assign t[91] = ~(t[66]);
  assign t[92] = t[156] ^ t[113];
  assign t[93] = t[8] ? t[114] : t[159];
  assign t[94] = t[157] ^ t[115];
  assign t[95] = ~(t[116]);
  assign t[96] = ~(t[117]);
  assign t[97] = ~(t[118]);
  assign t[98] = ~(t[119]);
  assign t[99] = t[44] ? t[120] : t[160];
  assign t[9] = t[142] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [111:0] x;
 output y;

 wire [323:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[118] ^ t[119];
  assign t[101] = t[119] ^ t[24];
  assign t[102] = ~(t[116]);
  assign t[103] = ~(t[121]);
  assign t[104] = ~(t[122]);
  assign t[105] = ~(t[123]);
  assign t[106] = t[44] ? t[124] : t[161];
  assign t[107] = t[122] ^ t[123];
  assign t[108] = t[123] ^ t[26];
  assign t[109] = ~(t[143]);
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[125] ? x[71] : x[70];
  assign t[111] = ~t[126];
  assign t[112] = t[8] ? t[127] : t[162];
  assign t[113] = t[125] ? x[76] : x[75];
  assign t[114] = t[159] ^ t[128];
  assign t[115] = t[31] ? x[78] : x[77];
  assign t[116] = ~(t[31]);
  assign t[117] = t[99] ^ t[119];
  assign t[118] = t[44] ? t[129] : t[163];
  assign t[119] = t[44] ? t[130] : t[164];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[160] ^ t[131];
  assign t[121] = t[106] ^ t[123];
  assign t[122] = t[44] ? t[132] : t[165];
  assign t[123] = t[44] ? t[133] : t[166];
  assign t[124] = t[161] ^ t[134];
  assign t[125] = ~(t[116]);
  assign t[126] = t[8] ? t[135] : t[167];
  assign t[127] = t[162] ^ t[136];
  assign t[128] = t[95] ? x[95] : x[94];
  assign t[129] = t[163] ^ t[137];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[164] ^ t[138];
  assign t[131] = t[95] ? x[97] : x[96];
  assign t[132] = t[165] ^ t[139];
  assign t[133] = t[166] ^ t[140];
  assign t[134] = t[102] ? x[99] : x[98];
  assign t[135] = t[167] ^ t[141];
  assign t[136] = t[125] ? x[101] : x[100];
  assign t[137] = t[95] ? x[103] : x[102];
  assign t[138] = t[95] ? x[105] : x[104];
  assign t[139] = t[102] ? x[107] : x[106];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[102] ? x[109] : x[108];
  assign t[141] = t[31] ? x[111] : x[110];
  assign t[142] = (t[168]);
  assign t[143] = (t[169]);
  assign t[144] = (t[170]);
  assign t[145] = (t[171]);
  assign t[146] = (t[172]);
  assign t[147] = (t[173]);
  assign t[148] = (t[174]);
  assign t[149] = (t[175]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = (t[176]);
  assign t[151] = (t[177]);
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = t[194] ^ x[4];
  assign t[169] = t[195] ^ x[7];
  assign t[16] = t[143] | t[30];
  assign t[170] = t[196] ^ x[12];
  assign t[171] = t[197] ^ x[15];
  assign t[172] = t[198] ^ x[18];
  assign t[173] = t[199] ^ x[21];
  assign t[174] = t[200] ^ x[24];
  assign t[175] = t[201] ^ x[27];
  assign t[176] = t[202] ^ x[30];
  assign t[177] = t[203] ^ x[33];
  assign t[178] = t[204] ^ x[36];
  assign t[179] = t[205] ^ x[39];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[206] ^ x[42];
  assign t[181] = t[207] ^ x[45];
  assign t[182] = t[208] ^ x[48];
  assign t[183] = t[209] ^ x[51];
  assign t[184] = t[210] ^ x[58];
  assign t[185] = t[211] ^ x[63];
  assign t[186] = t[212] ^ x[66];
  assign t[187] = t[213] ^ x[69];
  assign t[188] = t[214] ^ x[74];
  assign t[189] = t[215] ^ x[81];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[216] ^ x[84];
  assign t[191] = t[217] ^ x[87];
  assign t[192] = t[218] ^ x[90];
  assign t[193] = t[219] ^ x[93];
  assign t[194] = (t[220] & ~t[221]);
  assign t[195] = (t[222] & ~t[223]);
  assign t[196] = (t[224] & ~t[225]);
  assign t[197] = (t[226] & ~t[227]);
  assign t[198] = (t[228] & ~t[229]);
  assign t[199] = (t[230] & ~t[231]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[232] & ~t[233]);
  assign t[201] = (t[234] & ~t[235]);
  assign t[202] = (t[236] & ~t[237]);
  assign t[203] = (t[238] & ~t[239]);
  assign t[204] = (t[240] & ~t[241]);
  assign t[205] = (t[242] & ~t[243]);
  assign t[206] = (t[244] & ~t[245]);
  assign t[207] = (t[246] & ~t[247]);
  assign t[208] = (t[248] & ~t[249]);
  assign t[209] = (t[250] & ~t[251]);
  assign t[20] = t[36] ^ t[37];
  assign t[210] = (t[252] & ~t[253]);
  assign t[211] = (t[254] & ~t[255]);
  assign t[212] = (t[256] & ~t[257]);
  assign t[213] = (t[258] & ~t[259]);
  assign t[214] = (t[260] & ~t[261]);
  assign t[215] = (t[262] & ~t[263]);
  assign t[216] = (t[264] & ~t[265]);
  assign t[217] = (t[266] & ~t[267]);
  assign t[218] = (t[268] & ~t[269]);
  assign t[219] = (t[270] & ~t[271]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[272] ^ x[4];
  assign t[221] = t[273] ^ x[3];
  assign t[222] = t[274] ^ x[7];
  assign t[223] = t[275] ^ x[6];
  assign t[224] = t[276] ^ x[12];
  assign t[225] = t[277] ^ x[11];
  assign t[226] = t[278] ^ x[15];
  assign t[227] = t[279] ^ x[14];
  assign t[228] = t[280] ^ x[18];
  assign t[229] = t[281] ^ x[17];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[282] ^ x[21];
  assign t[231] = t[283] ^ x[20];
  assign t[232] = t[284] ^ x[24];
  assign t[233] = t[285] ^ x[23];
  assign t[234] = t[286] ^ x[27];
  assign t[235] = t[287] ^ x[26];
  assign t[236] = t[288] ^ x[30];
  assign t[237] = t[289] ^ x[29];
  assign t[238] = t[290] ^ x[33];
  assign t[239] = t[291] ^ x[32];
  assign t[23] = t[42] & t[43];
  assign t[240] = t[292] ^ x[36];
  assign t[241] = t[293] ^ x[35];
  assign t[242] = t[294] ^ x[39];
  assign t[243] = t[295] ^ x[38];
  assign t[244] = t[296] ^ x[42];
  assign t[245] = t[297] ^ x[41];
  assign t[246] = t[298] ^ x[45];
  assign t[247] = t[299] ^ x[44];
  assign t[248] = t[300] ^ x[48];
  assign t[249] = t[301] ^ x[47];
  assign t[24] = t[44] ? t[45] : t[144];
  assign t[250] = t[302] ^ x[51];
  assign t[251] = t[303] ^ x[50];
  assign t[252] = t[304] ^ x[58];
  assign t[253] = t[305] ^ x[57];
  assign t[254] = t[306] ^ x[63];
  assign t[255] = t[307] ^ x[62];
  assign t[256] = t[308] ^ x[66];
  assign t[257] = t[309] ^ x[65];
  assign t[258] = t[310] ^ x[69];
  assign t[259] = t[311] ^ x[68];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[312] ^ x[74];
  assign t[261] = t[313] ^ x[73];
  assign t[262] = t[314] ^ x[81];
  assign t[263] = t[315] ^ x[80];
  assign t[264] = t[316] ^ x[84];
  assign t[265] = t[317] ^ x[83];
  assign t[266] = t[318] ^ x[87];
  assign t[267] = t[319] ^ x[86];
  assign t[268] = t[320] ^ x[90];
  assign t[269] = t[321] ^ x[89];
  assign t[26] = t[44] ? t[48] : t[145];
  assign t[270] = t[322] ^ x[93];
  assign t[271] = t[323] ^ x[92];
  assign t[272] = (x[2]);
  assign t[273] = (x[2]);
  assign t[274] = (x[5]);
  assign t[275] = (x[5]);
  assign t[276] = (x[10]);
  assign t[277] = (x[10]);
  assign t[278] = (x[13]);
  assign t[279] = (x[13]);
  assign t[27] = t[49] ^ t[50];
  assign t[280] = (x[16]);
  assign t[281] = (x[16]);
  assign t[282] = (x[19]);
  assign t[283] = (x[19]);
  assign t[284] = (x[22]);
  assign t[285] = (x[22]);
  assign t[286] = (x[25]);
  assign t[287] = (x[25]);
  assign t[288] = (x[28]);
  assign t[289] = (x[28]);
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = (x[31]);
  assign t[291] = (x[31]);
  assign t[292] = (x[34]);
  assign t[293] = (x[34]);
  assign t[294] = (x[37]);
  assign t[295] = (x[37]);
  assign t[296] = (x[40]);
  assign t[297] = (x[40]);
  assign t[298] = (x[43]);
  assign t[299] = (x[43]);
  assign t[29] = ~(t[146] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[46]);
  assign t[301] = (x[46]);
  assign t[302] = (x[49]);
  assign t[303] = (x[49]);
  assign t[304] = (x[56]);
  assign t[305] = (x[56]);
  assign t[306] = (x[61]);
  assign t[307] = (x[61]);
  assign t[308] = (x[64]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = (x[67]);
  assign t[311] = (x[67]);
  assign t[312] = (x[72]);
  assign t[313] = (x[72]);
  assign t[314] = (x[79]);
  assign t[315] = (x[79]);
  assign t[316] = (x[82]);
  assign t[317] = (x[82]);
  assign t[318] = (x[85]);
  assign t[319] = (x[85]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[88]);
  assign t[321] = (x[88]);
  assign t[322] = (x[91]);
  assign t[323] = (x[91]);
  assign t[32] = ~(t[147]);
  assign t[33] = ~(t[148]);
  assign t[34] = ~(t[149]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = t[57];
  assign t[37] = t[4];
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[60] & t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[62] : t[150];
  assign t[41] = t[151] ^ t[63];
  assign t[42] = ~(t[64]);
  assign t[43] = t[152] ^ t[65];
  assign t[44] = ~(t[66]);
  assign t[45] = t[144] ^ t[67];
  assign t[46] = t[68] ^ t[69];
  assign t[47] = t[70] & t[71];
  assign t[48] = t[145] ^ t[72];
  assign t[49] = t[73] ^ t[74];
  assign t[4] = t[8] ? t[9] : t[142];
  assign t[50] = t[75] & t[76];
  assign t[51] = ~(t[77] & t[78]);
  assign t[52] = t[79] ^ t[153];
  assign t[53] = ~(t[146]);
  assign t[54] = t[80] & t[79];
  assign t[55] = ~(t[151]);
  assign t[56] = ~(t[81] & t[154]);
  assign t[57] = t[8] ? t[82] : t[155];
  assign t[58] = t[83] & t[84];
  assign t[59] = t[85] & t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = ~(t[58] ^ t[87]);
  assign t[61] = t[88] ^ t[89];
  assign t[62] = t[150] ^ t[90];
  assign t[63] = t[91] ? t[92] : t[156];
  assign t[64] = t[149] ^ t[93];
  assign t[65] = t[8] ? t[94] : t[157];
  assign t[66] = ~(t[8]);
  assign t[67] = t[95] ? x[53] : x[52];
  assign t[68] = t[96] & t[97];
  assign t[69] = t[98] & t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[100] ^ t[46]);
  assign t[71] = t[101] ^ t[99];
  assign t[72] = t[102] ? x[55] : x[54];
  assign t[73] = t[103] & t[104];
  assign t[74] = t[105] & t[106];
  assign t[75] = ~(t[107] ^ t[49]);
  assign t[76] = t[108] ^ t[106];
  assign t[77] = ~(t[80] | t[79]);
  assign t[78] = ~(t[109] | t[53]);
  assign t[79] = ~(t[158]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[153]);
  assign t[81] = ~(t[152]);
  assign t[82] = t[155] ^ t[110];
  assign t[83] = ~(t[89]);
  assign t[84] = ~(t[111]);
  assign t[85] = ~(t[36]);
  assign t[86] = t[112];
  assign t[87] = t[20] ^ t[111];
  assign t[88] = t[111] ^ t[37];
  assign t[89] = t[86] ^ t[36];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[95] ? x[60] : x[59];
  assign t[91] = ~(t[66]);
  assign t[92] = t[156] ^ t[113];
  assign t[93] = t[8] ? t[114] : t[159];
  assign t[94] = t[157] ^ t[115];
  assign t[95] = ~(t[116]);
  assign t[96] = ~(t[117]);
  assign t[97] = ~(t[118]);
  assign t[98] = ~(t[119]);
  assign t[99] = t[44] ? t[120] : t[160];
  assign t[9] = t[142] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind26(x, y);
 input [111:0] x;
 output y;

 wire [345:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[98] ^ t[131]);
  assign t[101] = t[132] ^ t[133];
  assign t[102] = t[105] ? x[72] : x[71];
  assign t[103] = t[179] ^ t[134];
  assign t[104] = t[105] ? x[74] : x[73];
  assign t[105] = ~(t[55]);
  assign t[106] = ~(t[135]);
  assign t[107] = ~(t[44]);
  assign t[108] = t[44] ^ t[72];
  assign t[109] = t[72] ^ t[26];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[165]);
  assign t[111] = ~(t[55]);
  assign t[112] = ~(t[136]);
  assign t[113] = ~(t[61]);
  assign t[114] = t[61] ^ t[90];
  assign t[115] = t[90] ^ t[36];
  assign t[116] = t[111] ? x[76] : x[75];
  assign t[117] = t[182] ^ t[137];
  assign t[118] = t[111] ? x[78] : x[77];
  assign t[119] = t[183] ^ t[138];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[8] ? t[139] : t[185];
  assign t[121] = t[140] ^ t[141];
  assign t[122] = t[93] ^ t[142];
  assign t[123] = t[181] ^ t[143];
  assign t[124] = t[184] ^ t[144];
  assign t[125] = ~(t[145] ^ t[69]);
  assign t[126] = t[42] ^ t[130];
  assign t[127] = ~(t[133]);
  assign t[128] = ~(t[146]);
  assign t[129] = ~(t[68]);
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[147];
  assign t[131] = t[42] ^ t[146];
  assign t[132] = t[146] ^ t[66];
  assign t[133] = t[130] ^ t[68];
  assign t[134] = t[105] ? x[83] : x[82];
  assign t[135] = t[46] ^ t[72];
  assign t[136] = t[63] ^ t[90];
  assign t[137] = t[111] ? x[85] : x[84];
  assign t[138] = t[111] ? x[87] : x[86];
  assign t[139] = t[185] ^ t[148];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[149] & t[150];
  assign t[141] = t[151] & t[123];
  assign t[142] = t[175] ^ t[152];
  assign t[143] = t[8] ? t[153] : t[186];
  assign t[144] = t[83] ? x[92] : x[91];
  assign t[145] = t[146] ^ t[68];
  assign t[146] = ~t[154];
  assign t[147] = t[8] ? t[155] : t[187];
  assign t[148] = t[111] ? x[97] : x[96];
  assign t[149] = ~(t[156]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = ~(t[92]);
  assign t[151] = ~(t[93]);
  assign t[152] = t[157] ? t[158] : t[188];
  assign t[153] = t[186] ^ t[159];
  assign t[154] = t[8] ? t[160] : t[189];
  assign t[155] = t[187] ^ t[161];
  assign t[156] = t[123] ^ t[93];
  assign t[157] = ~(t[74]);
  assign t[158] = t[188] ^ t[162];
  assign t[159] = t[83] ? x[105] : x[104];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[189] ^ t[163];
  assign t[161] = t[31] ? x[107] : x[106];
  assign t[162] = t[31] ? x[109] : x[108];
  assign t[163] = t[83] ? x[111] : x[110];
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[165] | t[30];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = (t[205]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[206]);
  assign t[181] = (t[207]);
  assign t[182] = (t[208]);
  assign t[183] = (t[209]);
  assign t[184] = (t[210]);
  assign t[185] = (t[211]);
  assign t[186] = (t[212]);
  assign t[187] = (t[213]);
  assign t[188] = (t[214]);
  assign t[189] = (t[215]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[216] ^ x[4];
  assign t[191] = t[217] ^ x[7];
  assign t[192] = t[218] ^ x[12];
  assign t[193] = t[219] ^ x[15];
  assign t[194] = t[220] ^ x[18];
  assign t[195] = t[221] ^ x[21];
  assign t[196] = t[222] ^ x[24];
  assign t[197] = t[223] ^ x[27];
  assign t[198] = t[224] ^ x[30];
  assign t[199] = t[225] ^ x[33];
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[36];
  assign t[201] = t[227] ^ x[39];
  assign t[202] = t[228] ^ x[42];
  assign t[203] = t[229] ^ x[45];
  assign t[204] = t[230] ^ x[48];
  assign t[205] = t[231] ^ x[51];
  assign t[206] = t[232] ^ x[56];
  assign t[207] = t[233] ^ x[59];
  assign t[208] = t[234] ^ x[64];
  assign t[209] = t[235] ^ x[67];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[236] ^ x[70];
  assign t[211] = t[237] ^ x[81];
  assign t[212] = t[238] ^ x[90];
  assign t[213] = t[239] ^ x[95];
  assign t[214] = t[240] ^ x[100];
  assign t[215] = t[241] ^ x[103];
  assign t[216] = (t[242] & ~t[243]);
  assign t[217] = (t[244] & ~t[245]);
  assign t[218] = (t[246] & ~t[247]);
  assign t[219] = (t[248] & ~t[249]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = (t[250] & ~t[251]);
  assign t[221] = (t[252] & ~t[253]);
  assign t[222] = (t[254] & ~t[255]);
  assign t[223] = (t[256] & ~t[257]);
  assign t[224] = (t[258] & ~t[259]);
  assign t[225] = (t[260] & ~t[261]);
  assign t[226] = (t[262] & ~t[263]);
  assign t[227] = (t[264] & ~t[265]);
  assign t[228] = (t[266] & ~t[267]);
  assign t[229] = (t[268] & ~t[269]);
  assign t[22] = ~(t[40] ^ t[41]);
  assign t[230] = (t[270] & ~t[271]);
  assign t[231] = (t[272] & ~t[273]);
  assign t[232] = (t[274] & ~t[275]);
  assign t[233] = (t[276] & ~t[277]);
  assign t[234] = (t[278] & ~t[279]);
  assign t[235] = (t[280] & ~t[281]);
  assign t[236] = (t[282] & ~t[283]);
  assign t[237] = (t[284] & ~t[285]);
  assign t[238] = (t[286] & ~t[287]);
  assign t[239] = (t[288] & ~t[289]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (t[290] & ~t[291]);
  assign t[241] = (t[292] & ~t[293]);
  assign t[242] = t[294] ^ x[4];
  assign t[243] = t[295] ^ x[3];
  assign t[244] = t[296] ^ x[7];
  assign t[245] = t[297] ^ x[6];
  assign t[246] = t[298] ^ x[12];
  assign t[247] = t[299] ^ x[11];
  assign t[248] = t[300] ^ x[15];
  assign t[249] = t[301] ^ x[14];
  assign t[24] = t[44] ^ t[26];
  assign t[250] = t[302] ^ x[18];
  assign t[251] = t[303] ^ x[17];
  assign t[252] = t[304] ^ x[21];
  assign t[253] = t[305] ^ x[20];
  assign t[254] = t[306] ^ x[24];
  assign t[255] = t[307] ^ x[23];
  assign t[256] = t[308] ^ x[27];
  assign t[257] = t[309] ^ x[26];
  assign t[258] = t[310] ^ x[30];
  assign t[259] = t[311] ^ x[29];
  assign t[25] = t[45] & t[46];
  assign t[260] = t[312] ^ x[33];
  assign t[261] = t[313] ^ x[32];
  assign t[262] = t[314] ^ x[36];
  assign t[263] = t[315] ^ x[35];
  assign t[264] = t[316] ^ x[39];
  assign t[265] = t[317] ^ x[38];
  assign t[266] = t[318] ^ x[42];
  assign t[267] = t[319] ^ x[41];
  assign t[268] = t[320] ^ x[45];
  assign t[269] = t[321] ^ x[44];
  assign t[26] = t[47] ? t[48] : t[166];
  assign t[270] = t[322] ^ x[48];
  assign t[271] = t[323] ^ x[47];
  assign t[272] = t[324] ^ x[51];
  assign t[273] = t[325] ^ x[50];
  assign t[274] = t[326] ^ x[56];
  assign t[275] = t[327] ^ x[55];
  assign t[276] = t[328] ^ x[59];
  assign t[277] = t[329] ^ x[58];
  assign t[278] = t[330] ^ x[64];
  assign t[279] = t[331] ^ x[63];
  assign t[27] = t[49] ^ t[50];
  assign t[280] = t[332] ^ x[67];
  assign t[281] = t[333] ^ x[66];
  assign t[282] = t[334] ^ x[70];
  assign t[283] = t[335] ^ x[69];
  assign t[284] = t[336] ^ x[81];
  assign t[285] = t[337] ^ x[80];
  assign t[286] = t[338] ^ x[90];
  assign t[287] = t[339] ^ x[89];
  assign t[288] = t[340] ^ x[95];
  assign t[289] = t[341] ^ x[94];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[342] ^ x[100];
  assign t[291] = t[343] ^ x[99];
  assign t[292] = t[344] ^ x[103];
  assign t[293] = t[345] ^ x[102];
  assign t[294] = (x[2]);
  assign t[295] = (x[2]);
  assign t[296] = (x[5]);
  assign t[297] = (x[5]);
  assign t[298] = (x[10]);
  assign t[299] = (x[10]);
  assign t[29] = ~(t[167] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[13]);
  assign t[301] = (x[13]);
  assign t[302] = (x[16]);
  assign t[303] = (x[16]);
  assign t[304] = (x[19]);
  assign t[305] = (x[19]);
  assign t[306] = (x[22]);
  assign t[307] = (x[22]);
  assign t[308] = (x[25]);
  assign t[309] = (x[25]);
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = (x[28]);
  assign t[311] = (x[28]);
  assign t[312] = (x[31]);
  assign t[313] = (x[31]);
  assign t[314] = (x[34]);
  assign t[315] = (x[34]);
  assign t[316] = (x[37]);
  assign t[317] = (x[37]);
  assign t[318] = (x[40]);
  assign t[319] = (x[40]);
  assign t[31] = ~(t[55]);
  assign t[320] = (x[43]);
  assign t[321] = (x[43]);
  assign t[322] = (x[46]);
  assign t[323] = (x[46]);
  assign t[324] = (x[49]);
  assign t[325] = (x[49]);
  assign t[326] = (x[54]);
  assign t[327] = (x[54]);
  assign t[328] = (x[57]);
  assign t[329] = (x[57]);
  assign t[32] = ~(t[168]);
  assign t[330] = (x[62]);
  assign t[331] = (x[62]);
  assign t[332] = (x[65]);
  assign t[333] = (x[65]);
  assign t[334] = (x[68]);
  assign t[335] = (x[68]);
  assign t[336] = (x[79]);
  assign t[337] = (x[79]);
  assign t[338] = (x[88]);
  assign t[339] = (x[88]);
  assign t[33] = ~(t[169]);
  assign t[340] = (x[93]);
  assign t[341] = (x[93]);
  assign t[342] = (x[98]);
  assign t[343] = (x[98]);
  assign t[344] = (x[101]);
  assign t[345] = (x[101]);
  assign t[34] = ~(t[170]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[36] = t[47] ? t[58] : t[171];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[61] ^ t[36];
  assign t[39] = t[62] & t[63];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[66] ^ t[67];
  assign t[42] = t[68] ^ t[66];
  assign t[43] = t[69] ^ t[70];
  assign t[44] = t[47] ? t[71] : t[172];
  assign t[45] = ~(t[72]);
  assign t[46] = t[47] ? t[73] : t[173];
  assign t[47] = ~(t[74]);
  assign t[48] = t[166] ^ t[75];
  assign t[49] = t[76] ^ t[25];
  assign t[4] = t[8] ? t[9] : t[164];
  assign t[50] = t[77] & t[78];
  assign t[51] = ~(t[79] & t[80]);
  assign t[52] = t[81] ^ t[174];
  assign t[53] = ~(t[167]);
  assign t[54] = t[82] & t[81];
  assign t[55] = ~(t[83]);
  assign t[56] = ~(t[175]);
  assign t[57] = ~(t[84] & t[176]);
  assign t[58] = t[171] ^ t[85];
  assign t[59] = t[86] ^ t[39];
  assign t[5] = ~(t[10]);
  assign t[60] = t[87] & t[88];
  assign t[61] = t[47] ? t[89] : t[177];
  assign t[62] = ~(t[90]);
  assign t[63] = t[47] ? t[91] : t[178];
  assign t[64] = t[92] ^ t[93];
  assign t[65] = t[94] & t[95];
  assign t[66] = t[96];
  assign t[67] = t[69] ^ t[97];
  assign t[68] = t[4];
  assign t[69] = t[98] ^ t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[100] & t[101];
  assign t[71] = t[172] ^ t[102];
  assign t[72] = t[47] ? t[103] : t[179];
  assign t[73] = t[173] ^ t[104];
  assign t[74] = ~(t[8]);
  assign t[75] = t[105] ? x[53] : x[52];
  assign t[76] = t[106] & t[107];
  assign t[77] = ~(t[108] ^ t[49]);
  assign t[78] = t[109] ^ t[46];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[110] | t[53]);
  assign t[81] = ~(t[180]);
  assign t[82] = ~(t[174]);
  assign t[83] = ~(t[16]);
  assign t[84] = ~(t[181]);
  assign t[85] = t[111] ? x[61] : x[60];
  assign t[86] = t[112] & t[113];
  assign t[87] = ~(t[114] ^ t[59]);
  assign t[88] = t[115] ^ t[63];
  assign t[89] = t[177] ^ t[116];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[47] ? t[117] : t[182];
  assign t[91] = t[178] ^ t[118];
  assign t[92] = t[8] ? t[119] : t[183];
  assign t[93] = t[170] ^ t[120];
  assign t[94] = ~(t[64] ^ t[121]);
  assign t[95] = t[122] ^ t[123];
  assign t[96] = t[8] ? t[124] : t[184];
  assign t[97] = t[125] & t[126];
  assign t[98] = t[127] & t[128];
  assign t[99] = t[129] & t[130];
  assign t[9] = t[164] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind27(x, y);
 input [111:0] x;
 output y;

 wire [345:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[98] ^ t[131]);
  assign t[101] = t[132] ^ t[133];
  assign t[102] = t[105] ? x[72] : x[71];
  assign t[103] = t[179] ^ t[134];
  assign t[104] = t[105] ? x[74] : x[73];
  assign t[105] = ~(t[55]);
  assign t[106] = ~(t[135]);
  assign t[107] = ~(t[44]);
  assign t[108] = t[44] ^ t[72];
  assign t[109] = t[72] ^ t[26];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[165]);
  assign t[111] = ~(t[55]);
  assign t[112] = ~(t[136]);
  assign t[113] = ~(t[61]);
  assign t[114] = t[61] ^ t[90];
  assign t[115] = t[90] ^ t[36];
  assign t[116] = t[111] ? x[76] : x[75];
  assign t[117] = t[182] ^ t[137];
  assign t[118] = t[111] ? x[78] : x[77];
  assign t[119] = t[183] ^ t[138];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[8] ? t[139] : t[185];
  assign t[121] = t[140] ^ t[141];
  assign t[122] = t[93] ^ t[142];
  assign t[123] = t[181] ^ t[143];
  assign t[124] = t[184] ^ t[144];
  assign t[125] = ~(t[145] ^ t[69]);
  assign t[126] = t[42] ^ t[130];
  assign t[127] = ~(t[133]);
  assign t[128] = ~(t[146]);
  assign t[129] = ~(t[68]);
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[147];
  assign t[131] = t[42] ^ t[146];
  assign t[132] = t[146] ^ t[66];
  assign t[133] = t[130] ^ t[68];
  assign t[134] = t[105] ? x[83] : x[82];
  assign t[135] = t[46] ^ t[72];
  assign t[136] = t[63] ^ t[90];
  assign t[137] = t[111] ? x[85] : x[84];
  assign t[138] = t[111] ? x[87] : x[86];
  assign t[139] = t[185] ^ t[148];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[149] & t[150];
  assign t[141] = t[151] & t[123];
  assign t[142] = t[175] ^ t[152];
  assign t[143] = t[8] ? t[153] : t[186];
  assign t[144] = t[83] ? x[92] : x[91];
  assign t[145] = t[146] ^ t[68];
  assign t[146] = ~t[154];
  assign t[147] = t[8] ? t[155] : t[187];
  assign t[148] = t[111] ? x[97] : x[96];
  assign t[149] = ~(t[156]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = ~(t[92]);
  assign t[151] = ~(t[93]);
  assign t[152] = t[157] ? t[158] : t[188];
  assign t[153] = t[186] ^ t[159];
  assign t[154] = t[8] ? t[160] : t[189];
  assign t[155] = t[187] ^ t[161];
  assign t[156] = t[123] ^ t[93];
  assign t[157] = ~(t[74]);
  assign t[158] = t[188] ^ t[162];
  assign t[159] = t[83] ? x[105] : x[104];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[189] ^ t[163];
  assign t[161] = t[31] ? x[107] : x[106];
  assign t[162] = t[31] ? x[109] : x[108];
  assign t[163] = t[83] ? x[111] : x[110];
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[165] | t[30];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = (t[205]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[206]);
  assign t[181] = (t[207]);
  assign t[182] = (t[208]);
  assign t[183] = (t[209]);
  assign t[184] = (t[210]);
  assign t[185] = (t[211]);
  assign t[186] = (t[212]);
  assign t[187] = (t[213]);
  assign t[188] = (t[214]);
  assign t[189] = (t[215]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[216] ^ x[4];
  assign t[191] = t[217] ^ x[7];
  assign t[192] = t[218] ^ x[12];
  assign t[193] = t[219] ^ x[15];
  assign t[194] = t[220] ^ x[18];
  assign t[195] = t[221] ^ x[21];
  assign t[196] = t[222] ^ x[24];
  assign t[197] = t[223] ^ x[27];
  assign t[198] = t[224] ^ x[30];
  assign t[199] = t[225] ^ x[33];
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[36];
  assign t[201] = t[227] ^ x[39];
  assign t[202] = t[228] ^ x[42];
  assign t[203] = t[229] ^ x[45];
  assign t[204] = t[230] ^ x[48];
  assign t[205] = t[231] ^ x[51];
  assign t[206] = t[232] ^ x[56];
  assign t[207] = t[233] ^ x[59];
  assign t[208] = t[234] ^ x[64];
  assign t[209] = t[235] ^ x[67];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[236] ^ x[70];
  assign t[211] = t[237] ^ x[81];
  assign t[212] = t[238] ^ x[90];
  assign t[213] = t[239] ^ x[95];
  assign t[214] = t[240] ^ x[100];
  assign t[215] = t[241] ^ x[103];
  assign t[216] = (t[242] & ~t[243]);
  assign t[217] = (t[244] & ~t[245]);
  assign t[218] = (t[246] & ~t[247]);
  assign t[219] = (t[248] & ~t[249]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = (t[250] & ~t[251]);
  assign t[221] = (t[252] & ~t[253]);
  assign t[222] = (t[254] & ~t[255]);
  assign t[223] = (t[256] & ~t[257]);
  assign t[224] = (t[258] & ~t[259]);
  assign t[225] = (t[260] & ~t[261]);
  assign t[226] = (t[262] & ~t[263]);
  assign t[227] = (t[264] & ~t[265]);
  assign t[228] = (t[266] & ~t[267]);
  assign t[229] = (t[268] & ~t[269]);
  assign t[22] = ~(t[40] ^ t[41]);
  assign t[230] = (t[270] & ~t[271]);
  assign t[231] = (t[272] & ~t[273]);
  assign t[232] = (t[274] & ~t[275]);
  assign t[233] = (t[276] & ~t[277]);
  assign t[234] = (t[278] & ~t[279]);
  assign t[235] = (t[280] & ~t[281]);
  assign t[236] = (t[282] & ~t[283]);
  assign t[237] = (t[284] & ~t[285]);
  assign t[238] = (t[286] & ~t[287]);
  assign t[239] = (t[288] & ~t[289]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (t[290] & ~t[291]);
  assign t[241] = (t[292] & ~t[293]);
  assign t[242] = t[294] ^ x[4];
  assign t[243] = t[295] ^ x[3];
  assign t[244] = t[296] ^ x[7];
  assign t[245] = t[297] ^ x[6];
  assign t[246] = t[298] ^ x[12];
  assign t[247] = t[299] ^ x[11];
  assign t[248] = t[300] ^ x[15];
  assign t[249] = t[301] ^ x[14];
  assign t[24] = t[44] ^ t[26];
  assign t[250] = t[302] ^ x[18];
  assign t[251] = t[303] ^ x[17];
  assign t[252] = t[304] ^ x[21];
  assign t[253] = t[305] ^ x[20];
  assign t[254] = t[306] ^ x[24];
  assign t[255] = t[307] ^ x[23];
  assign t[256] = t[308] ^ x[27];
  assign t[257] = t[309] ^ x[26];
  assign t[258] = t[310] ^ x[30];
  assign t[259] = t[311] ^ x[29];
  assign t[25] = t[45] & t[46];
  assign t[260] = t[312] ^ x[33];
  assign t[261] = t[313] ^ x[32];
  assign t[262] = t[314] ^ x[36];
  assign t[263] = t[315] ^ x[35];
  assign t[264] = t[316] ^ x[39];
  assign t[265] = t[317] ^ x[38];
  assign t[266] = t[318] ^ x[42];
  assign t[267] = t[319] ^ x[41];
  assign t[268] = t[320] ^ x[45];
  assign t[269] = t[321] ^ x[44];
  assign t[26] = t[47] ? t[48] : t[166];
  assign t[270] = t[322] ^ x[48];
  assign t[271] = t[323] ^ x[47];
  assign t[272] = t[324] ^ x[51];
  assign t[273] = t[325] ^ x[50];
  assign t[274] = t[326] ^ x[56];
  assign t[275] = t[327] ^ x[55];
  assign t[276] = t[328] ^ x[59];
  assign t[277] = t[329] ^ x[58];
  assign t[278] = t[330] ^ x[64];
  assign t[279] = t[331] ^ x[63];
  assign t[27] = t[49] ^ t[50];
  assign t[280] = t[332] ^ x[67];
  assign t[281] = t[333] ^ x[66];
  assign t[282] = t[334] ^ x[70];
  assign t[283] = t[335] ^ x[69];
  assign t[284] = t[336] ^ x[81];
  assign t[285] = t[337] ^ x[80];
  assign t[286] = t[338] ^ x[90];
  assign t[287] = t[339] ^ x[89];
  assign t[288] = t[340] ^ x[95];
  assign t[289] = t[341] ^ x[94];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[342] ^ x[100];
  assign t[291] = t[343] ^ x[99];
  assign t[292] = t[344] ^ x[103];
  assign t[293] = t[345] ^ x[102];
  assign t[294] = (x[2]);
  assign t[295] = (x[2]);
  assign t[296] = (x[5]);
  assign t[297] = (x[5]);
  assign t[298] = (x[10]);
  assign t[299] = (x[10]);
  assign t[29] = ~(t[167] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[13]);
  assign t[301] = (x[13]);
  assign t[302] = (x[16]);
  assign t[303] = (x[16]);
  assign t[304] = (x[19]);
  assign t[305] = (x[19]);
  assign t[306] = (x[22]);
  assign t[307] = (x[22]);
  assign t[308] = (x[25]);
  assign t[309] = (x[25]);
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = (x[28]);
  assign t[311] = (x[28]);
  assign t[312] = (x[31]);
  assign t[313] = (x[31]);
  assign t[314] = (x[34]);
  assign t[315] = (x[34]);
  assign t[316] = (x[37]);
  assign t[317] = (x[37]);
  assign t[318] = (x[40]);
  assign t[319] = (x[40]);
  assign t[31] = ~(t[55]);
  assign t[320] = (x[43]);
  assign t[321] = (x[43]);
  assign t[322] = (x[46]);
  assign t[323] = (x[46]);
  assign t[324] = (x[49]);
  assign t[325] = (x[49]);
  assign t[326] = (x[54]);
  assign t[327] = (x[54]);
  assign t[328] = (x[57]);
  assign t[329] = (x[57]);
  assign t[32] = ~(t[168]);
  assign t[330] = (x[62]);
  assign t[331] = (x[62]);
  assign t[332] = (x[65]);
  assign t[333] = (x[65]);
  assign t[334] = (x[68]);
  assign t[335] = (x[68]);
  assign t[336] = (x[79]);
  assign t[337] = (x[79]);
  assign t[338] = (x[88]);
  assign t[339] = (x[88]);
  assign t[33] = ~(t[169]);
  assign t[340] = (x[93]);
  assign t[341] = (x[93]);
  assign t[342] = (x[98]);
  assign t[343] = (x[98]);
  assign t[344] = (x[101]);
  assign t[345] = (x[101]);
  assign t[34] = ~(t[170]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[36] = t[47] ? t[58] : t[171];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[61] ^ t[36];
  assign t[39] = t[62] & t[63];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[66] ^ t[67];
  assign t[42] = t[68] ^ t[66];
  assign t[43] = t[69] ^ t[70];
  assign t[44] = t[47] ? t[71] : t[172];
  assign t[45] = ~(t[72]);
  assign t[46] = t[47] ? t[73] : t[173];
  assign t[47] = ~(t[74]);
  assign t[48] = t[166] ^ t[75];
  assign t[49] = t[76] ^ t[25];
  assign t[4] = t[8] ? t[9] : t[164];
  assign t[50] = t[77] & t[78];
  assign t[51] = ~(t[79] & t[80]);
  assign t[52] = t[81] ^ t[174];
  assign t[53] = ~(t[167]);
  assign t[54] = t[82] & t[81];
  assign t[55] = ~(t[83]);
  assign t[56] = ~(t[175]);
  assign t[57] = ~(t[84] & t[176]);
  assign t[58] = t[171] ^ t[85];
  assign t[59] = t[86] ^ t[39];
  assign t[5] = ~(t[10]);
  assign t[60] = t[87] & t[88];
  assign t[61] = t[47] ? t[89] : t[177];
  assign t[62] = ~(t[90]);
  assign t[63] = t[47] ? t[91] : t[178];
  assign t[64] = t[92] ^ t[93];
  assign t[65] = t[94] & t[95];
  assign t[66] = t[96];
  assign t[67] = t[69] ^ t[97];
  assign t[68] = t[4];
  assign t[69] = t[98] ^ t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[100] & t[101];
  assign t[71] = t[172] ^ t[102];
  assign t[72] = t[47] ? t[103] : t[179];
  assign t[73] = t[173] ^ t[104];
  assign t[74] = ~(t[8]);
  assign t[75] = t[105] ? x[53] : x[52];
  assign t[76] = t[106] & t[107];
  assign t[77] = ~(t[108] ^ t[49]);
  assign t[78] = t[109] ^ t[46];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[110] | t[53]);
  assign t[81] = ~(t[180]);
  assign t[82] = ~(t[174]);
  assign t[83] = ~(t[16]);
  assign t[84] = ~(t[181]);
  assign t[85] = t[111] ? x[61] : x[60];
  assign t[86] = t[112] & t[113];
  assign t[87] = ~(t[114] ^ t[59]);
  assign t[88] = t[115] ^ t[63];
  assign t[89] = t[177] ^ t[116];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[47] ? t[117] : t[182];
  assign t[91] = t[178] ^ t[118];
  assign t[92] = t[8] ? t[119] : t[183];
  assign t[93] = t[170] ^ t[120];
  assign t[94] = ~(t[64] ^ t[121]);
  assign t[95] = t[122] ^ t[123];
  assign t[96] = t[8] ? t[124] : t[184];
  assign t[97] = t[125] & t[126];
  assign t[98] = t[127] & t[128];
  assign t[99] = t[129] & t[130];
  assign t[9] = t[164] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind28(x, y);
 input [111:0] x;
 output y;

 wire [334:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[129] ^ t[130];
  assign t[101] = t[70] ^ t[131];
  assign t[102] = t[59] ? t[132] : t[175];
  assign t[103] = t[81] ? x[78] : x[77];
  assign t[104] = ~(t[133]);
  assign t[105] = ~(t[36]);
  assign t[106] = t[36] ^ t[58];
  assign t[107] = t[58] ^ t[26];
  assign t[108] = ~(t[154]);
  assign t[109] = t[81] ? x[80] : x[79];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[171] ^ t[134];
  assign t[111] = ~(t[54]);
  assign t[112] = ~(t[135]);
  assign t[113] = ~(t[39]);
  assign t[114] = ~(t[40]);
  assign t[115] = t[172] ^ t[136];
  assign t[116] = t[111] ? x[82] : x[81];
  assign t[117] = t[173] ^ t[137];
  assign t[118] = ~(t[85]);
  assign t[119] = t[174] ^ t[138];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = ~(t[126]);
  assign t[121] = ~(t[139]);
  assign t[122] = ~(t[65]);
  assign t[123] = t[170] ^ t[140];
  assign t[124] = t[43] ^ t[139];
  assign t[125] = t[139] ^ t[66];
  assign t[126] = t[123] ^ t[65];
  assign t[127] = t[141] ? x[84] : x[83];
  assign t[128] = t[141] ? x[86] : x[85];
  assign t[129] = t[142] & t[143];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[144] & t[102];
  assign t[131] = t[59] ? t[145] : t[176];
  assign t[132] = t[175] ^ t[146];
  assign t[133] = t[38] ^ t[58];
  assign t[134] = t[31] ? x[91] : x[90];
  assign t[135] = t[64] ^ t[40];
  assign t[136] = t[111] ? x[93] : x[92];
  assign t[137] = t[111] ? x[95] : x[94];
  assign t[138] = t[31] ? x[97] : x[96];
  assign t[139] = t[8] ? t[147] : t[177];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[8] ? t[148] : t[178];
  assign t[141] = ~(t[54]);
  assign t[142] = ~(t[149]);
  assign t[143] = ~(t[69]);
  assign t[144] = ~(t[70]);
  assign t[145] = t[176] ^ t[150];
  assign t[146] = t[141] ? x[105] : x[104];
  assign t[147] = t[177] ^ t[151];
  assign t[148] = t[178] ^ t[152];
  assign t[149] = t[102] ^ t[70];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[141] ? x[107] : x[106];
  assign t[151] = t[111] ? x[109] : x[108];
  assign t[152] = t[81] ? x[111] : x[110];
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[154] | t[30];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = t[205] ^ x[4];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[206] ^ x[7];
  assign t[181] = t[207] ^ x[12];
  assign t[182] = t[208] ^ x[15];
  assign t[183] = t[209] ^ x[18];
  assign t[184] = t[210] ^ x[21];
  assign t[185] = t[211] ^ x[24];
  assign t[186] = t[212] ^ x[27];
  assign t[187] = t[213] ^ x[30];
  assign t[188] = t[214] ^ x[33];
  assign t[189] = t[215] ^ x[36];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[216] ^ x[39];
  assign t[191] = t[217] ^ x[42];
  assign t[192] = t[218] ^ x[45];
  assign t[193] = t[219] ^ x[48];
  assign t[194] = t[220] ^ x[51];
  assign t[195] = t[221] ^ x[54];
  assign t[196] = t[222] ^ x[57];
  assign t[197] = t[223] ^ x[60];
  assign t[198] = t[224] ^ x[67];
  assign t[199] = t[225] ^ x[70];
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[73];
  assign t[201] = t[227] ^ x[76];
  assign t[202] = t[228] ^ x[89];
  assign t[203] = t[229] ^ x[100];
  assign t[204] = t[230] ^ x[103];
  assign t[205] = (t[231] & ~t[232]);
  assign t[206] = (t[233] & ~t[234]);
  assign t[207] = (t[235] & ~t[236]);
  assign t[208] = (t[237] & ~t[238]);
  assign t[209] = (t[239] & ~t[240]);
  assign t[20] = t[36] ^ t[26];
  assign t[210] = (t[241] & ~t[242]);
  assign t[211] = (t[243] & ~t[244]);
  assign t[212] = (t[245] & ~t[246]);
  assign t[213] = (t[247] & ~t[248]);
  assign t[214] = (t[249] & ~t[250]);
  assign t[215] = (t[251] & ~t[252]);
  assign t[216] = (t[253] & ~t[254]);
  assign t[217] = (t[255] & ~t[256]);
  assign t[218] = (t[257] & ~t[258]);
  assign t[219] = (t[259] & ~t[260]);
  assign t[21] = t[37] & t[38];
  assign t[220] = (t[261] & ~t[262]);
  assign t[221] = (t[263] & ~t[264]);
  assign t[222] = (t[265] & ~t[266]);
  assign t[223] = (t[267] & ~t[268]);
  assign t[224] = (t[269] & ~t[270]);
  assign t[225] = (t[271] & ~t[272]);
  assign t[226] = (t[273] & ~t[274]);
  assign t[227] = (t[275] & ~t[276]);
  assign t[228] = (t[277] & ~t[278]);
  assign t[229] = (t[279] & ~t[280]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[281] & ~t[282]);
  assign t[231] = t[283] ^ x[4];
  assign t[232] = t[284] ^ x[3];
  assign t[233] = t[285] ^ x[7];
  assign t[234] = t[286] ^ x[6];
  assign t[235] = t[287] ^ x[12];
  assign t[236] = t[288] ^ x[11];
  assign t[237] = t[289] ^ x[15];
  assign t[238] = t[290] ^ x[14];
  assign t[239] = t[291] ^ x[18];
  assign t[23] = t[41] & t[42];
  assign t[240] = t[292] ^ x[17];
  assign t[241] = t[293] ^ x[21];
  assign t[242] = t[294] ^ x[20];
  assign t[243] = t[295] ^ x[24];
  assign t[244] = t[296] ^ x[23];
  assign t[245] = t[297] ^ x[27];
  assign t[246] = t[298] ^ x[26];
  assign t[247] = t[299] ^ x[30];
  assign t[248] = t[300] ^ x[29];
  assign t[249] = t[301] ^ x[33];
  assign t[24] = t[43] ^ t[44];
  assign t[250] = t[302] ^ x[32];
  assign t[251] = t[303] ^ x[36];
  assign t[252] = t[304] ^ x[35];
  assign t[253] = t[305] ^ x[39];
  assign t[254] = t[306] ^ x[38];
  assign t[255] = t[307] ^ x[42];
  assign t[256] = t[308] ^ x[41];
  assign t[257] = t[309] ^ x[45];
  assign t[258] = t[310] ^ x[44];
  assign t[259] = t[311] ^ x[48];
  assign t[25] = t[45] ^ t[46];
  assign t[260] = t[312] ^ x[47];
  assign t[261] = t[313] ^ x[51];
  assign t[262] = t[314] ^ x[50];
  assign t[263] = t[315] ^ x[54];
  assign t[264] = t[316] ^ x[53];
  assign t[265] = t[317] ^ x[57];
  assign t[266] = t[318] ^ x[56];
  assign t[267] = t[319] ^ x[60];
  assign t[268] = t[320] ^ x[59];
  assign t[269] = t[321] ^ x[67];
  assign t[26] = t[47];
  assign t[270] = t[322] ^ x[66];
  assign t[271] = t[323] ^ x[70];
  assign t[272] = t[324] ^ x[69];
  assign t[273] = t[325] ^ x[73];
  assign t[274] = t[326] ^ x[72];
  assign t[275] = t[327] ^ x[76];
  assign t[276] = t[328] ^ x[75];
  assign t[277] = t[329] ^ x[89];
  assign t[278] = t[330] ^ x[88];
  assign t[279] = t[331] ^ x[100];
  assign t[27] = t[48] ^ t[49];
  assign t[280] = t[332] ^ x[99];
  assign t[281] = t[333] ^ x[103];
  assign t[282] = t[334] ^ x[102];
  assign t[283] = (x[2]);
  assign t[284] = (x[2]);
  assign t[285] = (x[5]);
  assign t[286] = (x[5]);
  assign t[287] = (x[10]);
  assign t[288] = (x[10]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[30] & t[50]);
  assign t[290] = (x[13]);
  assign t[291] = (x[16]);
  assign t[292] = (x[16]);
  assign t[293] = (x[19]);
  assign t[294] = (x[19]);
  assign t[295] = (x[22]);
  assign t[296] = (x[22]);
  assign t[297] = (x[25]);
  assign t[298] = (x[25]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155] ^ t[51]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[28]);
  assign t[301] = (x[31]);
  assign t[302] = (x[31]);
  assign t[303] = (x[34]);
  assign t[304] = (x[34]);
  assign t[305] = (x[37]);
  assign t[306] = (x[37]);
  assign t[307] = (x[40]);
  assign t[308] = (x[40]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[52] & t[53]);
  assign t[310] = (x[43]);
  assign t[311] = (x[46]);
  assign t[312] = (x[46]);
  assign t[313] = (x[49]);
  assign t[314] = (x[49]);
  assign t[315] = (x[52]);
  assign t[316] = (x[52]);
  assign t[317] = (x[55]);
  assign t[318] = (x[55]);
  assign t[319] = (x[58]);
  assign t[31] = ~(t[54]);
  assign t[320] = (x[58]);
  assign t[321] = (x[65]);
  assign t[322] = (x[65]);
  assign t[323] = (x[68]);
  assign t[324] = (x[68]);
  assign t[325] = (x[71]);
  assign t[326] = (x[71]);
  assign t[327] = (x[74]);
  assign t[328] = (x[74]);
  assign t[329] = (x[87]);
  assign t[32] = ~(t[156]);
  assign t[330] = (x[87]);
  assign t[331] = (x[98]);
  assign t[332] = (x[98]);
  assign t[333] = (x[101]);
  assign t[334] = (x[101]);
  assign t[33] = ~(t[157]);
  assign t[34] = ~(t[158]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~t[57];
  assign t[37] = ~(t[58]);
  assign t[38] = t[4];
  assign t[39] = t[59] ? t[60] : t[159];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[59] ? t[61] : t[160];
  assign t[41] = ~(t[22] ^ t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[65] ^ t[66];
  assign t[44] = t[67] ^ t[68];
  assign t[45] = t[69] ^ t[70];
  assign t[46] = t[71] & t[72];
  assign t[47] = t[8] ? t[73] : t[161];
  assign t[48] = t[74] ^ t[21];
  assign t[49] = t[75] & t[76];
  assign t[4] = t[8] ? t[9] : t[153];
  assign t[50] = ~(t[77] & t[78]);
  assign t[51] = t[79] ^ t[162];
  assign t[52] = ~(t[155]);
  assign t[53] = t[80] & t[79];
  assign t[54] = ~(t[81]);
  assign t[55] = ~(t[163]);
  assign t[56] = ~(t[82] & t[164]);
  assign t[57] = t[8] ? t[83] : t[165];
  assign t[58] = t[84];
  assign t[59] = ~(t[85]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[159] ^ t[86];
  assign t[61] = t[160] ^ t[87];
  assign t[62] = t[88] ^ t[89];
  assign t[63] = t[40] ^ t[90];
  assign t[64] = t[59] ? t[91] : t[166];
  assign t[65] = t[158] ^ t[92];
  assign t[66] = t[163] ^ t[93];
  assign t[67] = t[94] ^ t[95];
  assign t[68] = t[96] & t[97];
  assign t[69] = t[59] ? t[98] : t[167];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[59] ? t[99] : t[168];
  assign t[71] = ~(t[45] ^ t[100]);
  assign t[72] = t[101] ^ t[102];
  assign t[73] = t[161] ^ t[103];
  assign t[74] = t[104] & t[105];
  assign t[75] = ~(t[106] ^ t[48]);
  assign t[76] = t[107] ^ t[38];
  assign t[77] = ~(t[80] | t[79]);
  assign t[78] = ~(t[108] | t[52]);
  assign t[79] = ~(t[169]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[162]);
  assign t[81] = ~(t[16]);
  assign t[82] = ~(t[170]);
  assign t[83] = t[165] ^ t[109];
  assign t[84] = t[8] ? t[110] : t[171];
  assign t[85] = ~(t[8]);
  assign t[86] = t[111] ? x[62] : x[61];
  assign t[87] = t[111] ? x[64] : x[63];
  assign t[88] = t[112] & t[113];
  assign t[89] = t[114] & t[64];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[59] ? t[115] : t[172];
  assign t[91] = t[166] ^ t[116];
  assign t[92] = t[8] ? t[117] : t[173];
  assign t[93] = t[118] ? t[119] : t[174];
  assign t[94] = t[120] & t[121];
  assign t[95] = t[122] & t[123];
  assign t[96] = ~(t[94] ^ t[124]);
  assign t[97] = t[125] ^ t[126];
  assign t[98] = t[167] ^ t[127];
  assign t[99] = t[168] ^ t[128];
  assign t[9] = t[153] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind29(x, y);
 input [111:0] x;
 output y;

 wire [334:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[129] ^ t[130];
  assign t[101] = t[70] ^ t[131];
  assign t[102] = t[59] ? t[132] : t[175];
  assign t[103] = t[81] ? x[78] : x[77];
  assign t[104] = ~(t[133]);
  assign t[105] = ~(t[36]);
  assign t[106] = t[36] ^ t[58];
  assign t[107] = t[58] ^ t[26];
  assign t[108] = ~(t[154]);
  assign t[109] = t[81] ? x[80] : x[79];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[171] ^ t[134];
  assign t[111] = ~(t[54]);
  assign t[112] = ~(t[135]);
  assign t[113] = ~(t[39]);
  assign t[114] = ~(t[40]);
  assign t[115] = t[172] ^ t[136];
  assign t[116] = t[111] ? x[82] : x[81];
  assign t[117] = t[173] ^ t[137];
  assign t[118] = ~(t[85]);
  assign t[119] = t[174] ^ t[138];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = ~(t[126]);
  assign t[121] = ~(t[139]);
  assign t[122] = ~(t[65]);
  assign t[123] = t[170] ^ t[140];
  assign t[124] = t[43] ^ t[139];
  assign t[125] = t[139] ^ t[66];
  assign t[126] = t[123] ^ t[65];
  assign t[127] = t[141] ? x[84] : x[83];
  assign t[128] = t[141] ? x[86] : x[85];
  assign t[129] = t[142] & t[143];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[144] & t[102];
  assign t[131] = t[59] ? t[145] : t[176];
  assign t[132] = t[175] ^ t[146];
  assign t[133] = t[38] ^ t[58];
  assign t[134] = t[31] ? x[91] : x[90];
  assign t[135] = t[64] ^ t[40];
  assign t[136] = t[111] ? x[93] : x[92];
  assign t[137] = t[111] ? x[95] : x[94];
  assign t[138] = t[31] ? x[97] : x[96];
  assign t[139] = t[8] ? t[147] : t[177];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[8] ? t[148] : t[178];
  assign t[141] = ~(t[54]);
  assign t[142] = ~(t[149]);
  assign t[143] = ~(t[69]);
  assign t[144] = ~(t[70]);
  assign t[145] = t[176] ^ t[150];
  assign t[146] = t[141] ? x[105] : x[104];
  assign t[147] = t[177] ^ t[151];
  assign t[148] = t[178] ^ t[152];
  assign t[149] = t[102] ^ t[70];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[141] ? x[107] : x[106];
  assign t[151] = t[111] ? x[109] : x[108];
  assign t[152] = t[81] ? x[111] : x[110];
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[154] | t[30];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = t[205] ^ x[4];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[206] ^ x[7];
  assign t[181] = t[207] ^ x[12];
  assign t[182] = t[208] ^ x[15];
  assign t[183] = t[209] ^ x[18];
  assign t[184] = t[210] ^ x[21];
  assign t[185] = t[211] ^ x[24];
  assign t[186] = t[212] ^ x[27];
  assign t[187] = t[213] ^ x[30];
  assign t[188] = t[214] ^ x[33];
  assign t[189] = t[215] ^ x[36];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[216] ^ x[39];
  assign t[191] = t[217] ^ x[42];
  assign t[192] = t[218] ^ x[45];
  assign t[193] = t[219] ^ x[48];
  assign t[194] = t[220] ^ x[51];
  assign t[195] = t[221] ^ x[54];
  assign t[196] = t[222] ^ x[57];
  assign t[197] = t[223] ^ x[60];
  assign t[198] = t[224] ^ x[67];
  assign t[199] = t[225] ^ x[70];
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[73];
  assign t[201] = t[227] ^ x[76];
  assign t[202] = t[228] ^ x[89];
  assign t[203] = t[229] ^ x[100];
  assign t[204] = t[230] ^ x[103];
  assign t[205] = (t[231] & ~t[232]);
  assign t[206] = (t[233] & ~t[234]);
  assign t[207] = (t[235] & ~t[236]);
  assign t[208] = (t[237] & ~t[238]);
  assign t[209] = (t[239] & ~t[240]);
  assign t[20] = t[36] ^ t[26];
  assign t[210] = (t[241] & ~t[242]);
  assign t[211] = (t[243] & ~t[244]);
  assign t[212] = (t[245] & ~t[246]);
  assign t[213] = (t[247] & ~t[248]);
  assign t[214] = (t[249] & ~t[250]);
  assign t[215] = (t[251] & ~t[252]);
  assign t[216] = (t[253] & ~t[254]);
  assign t[217] = (t[255] & ~t[256]);
  assign t[218] = (t[257] & ~t[258]);
  assign t[219] = (t[259] & ~t[260]);
  assign t[21] = t[37] & t[38];
  assign t[220] = (t[261] & ~t[262]);
  assign t[221] = (t[263] & ~t[264]);
  assign t[222] = (t[265] & ~t[266]);
  assign t[223] = (t[267] & ~t[268]);
  assign t[224] = (t[269] & ~t[270]);
  assign t[225] = (t[271] & ~t[272]);
  assign t[226] = (t[273] & ~t[274]);
  assign t[227] = (t[275] & ~t[276]);
  assign t[228] = (t[277] & ~t[278]);
  assign t[229] = (t[279] & ~t[280]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[281] & ~t[282]);
  assign t[231] = t[283] ^ x[4];
  assign t[232] = t[284] ^ x[3];
  assign t[233] = t[285] ^ x[7];
  assign t[234] = t[286] ^ x[6];
  assign t[235] = t[287] ^ x[12];
  assign t[236] = t[288] ^ x[11];
  assign t[237] = t[289] ^ x[15];
  assign t[238] = t[290] ^ x[14];
  assign t[239] = t[291] ^ x[18];
  assign t[23] = t[41] & t[42];
  assign t[240] = t[292] ^ x[17];
  assign t[241] = t[293] ^ x[21];
  assign t[242] = t[294] ^ x[20];
  assign t[243] = t[295] ^ x[24];
  assign t[244] = t[296] ^ x[23];
  assign t[245] = t[297] ^ x[27];
  assign t[246] = t[298] ^ x[26];
  assign t[247] = t[299] ^ x[30];
  assign t[248] = t[300] ^ x[29];
  assign t[249] = t[301] ^ x[33];
  assign t[24] = t[43] ^ t[44];
  assign t[250] = t[302] ^ x[32];
  assign t[251] = t[303] ^ x[36];
  assign t[252] = t[304] ^ x[35];
  assign t[253] = t[305] ^ x[39];
  assign t[254] = t[306] ^ x[38];
  assign t[255] = t[307] ^ x[42];
  assign t[256] = t[308] ^ x[41];
  assign t[257] = t[309] ^ x[45];
  assign t[258] = t[310] ^ x[44];
  assign t[259] = t[311] ^ x[48];
  assign t[25] = t[45] ^ t[46];
  assign t[260] = t[312] ^ x[47];
  assign t[261] = t[313] ^ x[51];
  assign t[262] = t[314] ^ x[50];
  assign t[263] = t[315] ^ x[54];
  assign t[264] = t[316] ^ x[53];
  assign t[265] = t[317] ^ x[57];
  assign t[266] = t[318] ^ x[56];
  assign t[267] = t[319] ^ x[60];
  assign t[268] = t[320] ^ x[59];
  assign t[269] = t[321] ^ x[67];
  assign t[26] = t[47];
  assign t[270] = t[322] ^ x[66];
  assign t[271] = t[323] ^ x[70];
  assign t[272] = t[324] ^ x[69];
  assign t[273] = t[325] ^ x[73];
  assign t[274] = t[326] ^ x[72];
  assign t[275] = t[327] ^ x[76];
  assign t[276] = t[328] ^ x[75];
  assign t[277] = t[329] ^ x[89];
  assign t[278] = t[330] ^ x[88];
  assign t[279] = t[331] ^ x[100];
  assign t[27] = t[48] ^ t[49];
  assign t[280] = t[332] ^ x[99];
  assign t[281] = t[333] ^ x[103];
  assign t[282] = t[334] ^ x[102];
  assign t[283] = (x[2]);
  assign t[284] = (x[2]);
  assign t[285] = (x[5]);
  assign t[286] = (x[5]);
  assign t[287] = (x[10]);
  assign t[288] = (x[10]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[30] & t[50]);
  assign t[290] = (x[13]);
  assign t[291] = (x[16]);
  assign t[292] = (x[16]);
  assign t[293] = (x[19]);
  assign t[294] = (x[19]);
  assign t[295] = (x[22]);
  assign t[296] = (x[22]);
  assign t[297] = (x[25]);
  assign t[298] = (x[25]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155] ^ t[51]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[28]);
  assign t[301] = (x[31]);
  assign t[302] = (x[31]);
  assign t[303] = (x[34]);
  assign t[304] = (x[34]);
  assign t[305] = (x[37]);
  assign t[306] = (x[37]);
  assign t[307] = (x[40]);
  assign t[308] = (x[40]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[52] & t[53]);
  assign t[310] = (x[43]);
  assign t[311] = (x[46]);
  assign t[312] = (x[46]);
  assign t[313] = (x[49]);
  assign t[314] = (x[49]);
  assign t[315] = (x[52]);
  assign t[316] = (x[52]);
  assign t[317] = (x[55]);
  assign t[318] = (x[55]);
  assign t[319] = (x[58]);
  assign t[31] = ~(t[54]);
  assign t[320] = (x[58]);
  assign t[321] = (x[65]);
  assign t[322] = (x[65]);
  assign t[323] = (x[68]);
  assign t[324] = (x[68]);
  assign t[325] = (x[71]);
  assign t[326] = (x[71]);
  assign t[327] = (x[74]);
  assign t[328] = (x[74]);
  assign t[329] = (x[87]);
  assign t[32] = ~(t[156]);
  assign t[330] = (x[87]);
  assign t[331] = (x[98]);
  assign t[332] = (x[98]);
  assign t[333] = (x[101]);
  assign t[334] = (x[101]);
  assign t[33] = ~(t[157]);
  assign t[34] = ~(t[158]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~t[57];
  assign t[37] = ~(t[58]);
  assign t[38] = t[4];
  assign t[39] = t[59] ? t[60] : t[159];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[59] ? t[61] : t[160];
  assign t[41] = ~(t[22] ^ t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[65] ^ t[66];
  assign t[44] = t[67] ^ t[68];
  assign t[45] = t[69] ^ t[70];
  assign t[46] = t[71] & t[72];
  assign t[47] = t[8] ? t[73] : t[161];
  assign t[48] = t[74] ^ t[21];
  assign t[49] = t[75] & t[76];
  assign t[4] = t[8] ? t[9] : t[153];
  assign t[50] = ~(t[77] & t[78]);
  assign t[51] = t[79] ^ t[162];
  assign t[52] = ~(t[155]);
  assign t[53] = t[80] & t[79];
  assign t[54] = ~(t[81]);
  assign t[55] = ~(t[163]);
  assign t[56] = ~(t[82] & t[164]);
  assign t[57] = t[8] ? t[83] : t[165];
  assign t[58] = t[84];
  assign t[59] = ~(t[85]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[159] ^ t[86];
  assign t[61] = t[160] ^ t[87];
  assign t[62] = t[88] ^ t[89];
  assign t[63] = t[40] ^ t[90];
  assign t[64] = t[59] ? t[91] : t[166];
  assign t[65] = t[158] ^ t[92];
  assign t[66] = t[163] ^ t[93];
  assign t[67] = t[94] ^ t[95];
  assign t[68] = t[96] & t[97];
  assign t[69] = t[59] ? t[98] : t[167];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[59] ? t[99] : t[168];
  assign t[71] = ~(t[45] ^ t[100]);
  assign t[72] = t[101] ^ t[102];
  assign t[73] = t[161] ^ t[103];
  assign t[74] = t[104] & t[105];
  assign t[75] = ~(t[106] ^ t[48]);
  assign t[76] = t[107] ^ t[38];
  assign t[77] = ~(t[80] | t[79]);
  assign t[78] = ~(t[108] | t[52]);
  assign t[79] = ~(t[169]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[162]);
  assign t[81] = ~(t[16]);
  assign t[82] = ~(t[170]);
  assign t[83] = t[165] ^ t[109];
  assign t[84] = t[8] ? t[110] : t[171];
  assign t[85] = ~(t[8]);
  assign t[86] = t[111] ? x[62] : x[61];
  assign t[87] = t[111] ? x[64] : x[63];
  assign t[88] = t[112] & t[113];
  assign t[89] = t[114] & t[64];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[59] ? t[115] : t[172];
  assign t[91] = t[166] ^ t[116];
  assign t[92] = t[8] ? t[117] : t[173];
  assign t[93] = t[118] ? t[119] : t[174];
  assign t[94] = t[120] & t[121];
  assign t[95] = t[122] & t[123];
  assign t[96] = ~(t[94] ^ t[124]);
  assign t[97] = t[125] ^ t[126];
  assign t[98] = t[167] ^ t[127];
  assign t[99] = t[168] ^ t[128];
  assign t[9] = t[153] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [111:0] x;
 output y;

 wire [333:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[126]);
  assign t[101] = t[44] ? t[127] : t[171];
  assign t[102] = t[167] ^ t[128];
  assign t[103] = ~(t[153]);
  assign t[104] = t[129] ? x[69] : x[68];
  assign t[105] = t[129] ? x[71] : x[70];
  assign t[106] = ~(t[112]);
  assign t[107] = ~(t[130]);
  assign t[108] = ~(t[57]);
  assign t[109] = t[44] ? t[131] : t[172];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[36] ^ t[130];
  assign t[111] = t[130] ^ t[58];
  assign t[112] = t[109] ^ t[57];
  assign t[113] = t[132] ? x[76] : x[75];
  assign t[114] = ~(t[133]);
  assign t[115] = ~(t[134]);
  assign t[116] = ~(t[135]);
  assign t[117] = t[169] ^ t[136];
  assign t[118] = t[134] ^ t[135];
  assign t[119] = t[135] ^ t[38];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[132] ? x[78] : x[77];
  assign t[121] = ~(t[137]);
  assign t[122] = ~(t[40]);
  assign t[123] = ~(t[41]);
  assign t[124] = t[8] ? t[138] : t[173];
  assign t[125] = t[170] ^ t[139];
  assign t[126] = ~(t[31]);
  assign t[127] = t[171] ^ t[140];
  assign t[128] = t[100] ? x[83] : x[82];
  assign t[129] = ~(t[126]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[44] ? t[141] : t[174];
  assign t[131] = t[172] ^ t[142];
  assign t[132] = ~(t[126]);
  assign t[133] = t[117] ^ t[135];
  assign t[134] = t[8] ? t[143] : t[175];
  assign t[135] = t[159] ^ t[144];
  assign t[136] = t[8] ? t[145] : t[176];
  assign t[137] = t[67] ^ t[41];
  assign t[138] = t[173] ^ t[146];
  assign t[139] = t[132] ? x[94] : x[93];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[100] ? x[96] : x[95];
  assign t[141] = t[174] ^ t[147];
  assign t[142] = t[129] ? x[98] : x[97];
  assign t[143] = t[175] ^ t[148];
  assign t[144] = t[8] ? t[149] : t[177];
  assign t[145] = t[176] ^ t[150];
  assign t[146] = t[31] ? x[103] : x[102];
  assign t[147] = t[129] ? x[105] : x[104];
  assign t[148] = t[100] ? x[107] : x[106];
  assign t[149] = t[177] ^ t[151];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[31] ? x[109] : x[108];
  assign t[151] = t[100] ? x[111] : x[110];
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[153] | t[30];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = t[204] ^ x[4];
  assign t[179] = t[205] ^ x[7];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[206] ^ x[12];
  assign t[181] = t[207] ^ x[15];
  assign t[182] = t[208] ^ x[18];
  assign t[183] = t[209] ^ x[21];
  assign t[184] = t[210] ^ x[24];
  assign t[185] = t[211] ^ x[27];
  assign t[186] = t[212] ^ x[30];
  assign t[187] = t[213] ^ x[33];
  assign t[188] = t[214] ^ x[36];
  assign t[189] = t[215] ^ x[39];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[216] ^ x[42];
  assign t[191] = t[217] ^ x[45];
  assign t[192] = t[218] ^ x[48];
  assign t[193] = t[219] ^ x[55];
  assign t[194] = t[220] ^ x[58];
  assign t[195] = t[221] ^ x[61];
  assign t[196] = t[222] ^ x[64];
  assign t[197] = t[223] ^ x[67];
  assign t[198] = t[224] ^ x[74];
  assign t[199] = t[225] ^ x[81];
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[86];
  assign t[201] = t[227] ^ x[89];
  assign t[202] = t[228] ^ x[92];
  assign t[203] = t[229] ^ x[101];
  assign t[204] = (t[230] & ~t[231]);
  assign t[205] = (t[232] & ~t[233]);
  assign t[206] = (t[234] & ~t[235]);
  assign t[207] = (t[236] & ~t[237]);
  assign t[208] = (t[238] & ~t[239]);
  assign t[209] = (t[240] & ~t[241]);
  assign t[20] = t[36] ^ t[37];
  assign t[210] = (t[242] & ~t[243]);
  assign t[211] = (t[244] & ~t[245]);
  assign t[212] = (t[246] & ~t[247]);
  assign t[213] = (t[248] & ~t[249]);
  assign t[214] = (t[250] & ~t[251]);
  assign t[215] = (t[252] & ~t[253]);
  assign t[216] = (t[254] & ~t[255]);
  assign t[217] = (t[256] & ~t[257]);
  assign t[218] = (t[258] & ~t[259]);
  assign t[219] = (t[260] & ~t[261]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = (t[262] & ~t[263]);
  assign t[221] = (t[264] & ~t[265]);
  assign t[222] = (t[266] & ~t[267]);
  assign t[223] = (t[268] & ~t[269]);
  assign t[224] = (t[270] & ~t[271]);
  assign t[225] = (t[272] & ~t[273]);
  assign t[226] = (t[274] & ~t[275]);
  assign t[227] = (t[276] & ~t[277]);
  assign t[228] = (t[278] & ~t[279]);
  assign t[229] = (t[280] & ~t[281]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[282] ^ x[4];
  assign t[231] = t[283] ^ x[3];
  assign t[232] = t[284] ^ x[7];
  assign t[233] = t[285] ^ x[6];
  assign t[234] = t[286] ^ x[12];
  assign t[235] = t[287] ^ x[11];
  assign t[236] = t[288] ^ x[15];
  assign t[237] = t[289] ^ x[14];
  assign t[238] = t[290] ^ x[18];
  assign t[239] = t[291] ^ x[17];
  assign t[23] = t[42] & t[43];
  assign t[240] = t[292] ^ x[21];
  assign t[241] = t[293] ^ x[20];
  assign t[242] = t[294] ^ x[24];
  assign t[243] = t[295] ^ x[23];
  assign t[244] = t[296] ^ x[27];
  assign t[245] = t[297] ^ x[26];
  assign t[246] = t[298] ^ x[30];
  assign t[247] = t[299] ^ x[29];
  assign t[248] = t[300] ^ x[33];
  assign t[249] = t[301] ^ x[32];
  assign t[24] = t[44] ? t[45] : t[154];
  assign t[250] = t[302] ^ x[36];
  assign t[251] = t[303] ^ x[35];
  assign t[252] = t[304] ^ x[39];
  assign t[253] = t[305] ^ x[38];
  assign t[254] = t[306] ^ x[42];
  assign t[255] = t[307] ^ x[41];
  assign t[256] = t[308] ^ x[45];
  assign t[257] = t[309] ^ x[44];
  assign t[258] = t[310] ^ x[48];
  assign t[259] = t[311] ^ x[47];
  assign t[25] = t[44] ? t[46] : t[155];
  assign t[260] = t[312] ^ x[55];
  assign t[261] = t[313] ^ x[54];
  assign t[262] = t[314] ^ x[58];
  assign t[263] = t[315] ^ x[57];
  assign t[264] = t[316] ^ x[61];
  assign t[265] = t[317] ^ x[60];
  assign t[266] = t[318] ^ x[64];
  assign t[267] = t[319] ^ x[63];
  assign t[268] = t[320] ^ x[67];
  assign t[269] = t[321] ^ x[66];
  assign t[26] = t[47] ^ t[48];
  assign t[270] = t[322] ^ x[74];
  assign t[271] = t[323] ^ x[73];
  assign t[272] = t[324] ^ x[81];
  assign t[273] = t[325] ^ x[80];
  assign t[274] = t[326] ^ x[86];
  assign t[275] = t[327] ^ x[85];
  assign t[276] = t[328] ^ x[89];
  assign t[277] = t[329] ^ x[88];
  assign t[278] = t[330] ^ x[92];
  assign t[279] = t[331] ^ x[91];
  assign t[27] = t[49] & t[50];
  assign t[280] = t[332] ^ x[101];
  assign t[281] = t[333] ^ x[100];
  assign t[282] = (x[2]);
  assign t[283] = (x[2]);
  assign t[284] = (x[5]);
  assign t[285] = (x[5]);
  assign t[286] = (x[10]);
  assign t[287] = (x[10]);
  assign t[288] = (x[13]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = (x[16]);
  assign t[291] = (x[16]);
  assign t[292] = (x[19]);
  assign t[293] = (x[19]);
  assign t[294] = (x[22]);
  assign t[295] = (x[22]);
  assign t[296] = (x[25]);
  assign t[297] = (x[25]);
  assign t[298] = (x[28]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[156] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[31]);
  assign t[301] = (x[31]);
  assign t[302] = (x[34]);
  assign t[303] = (x[34]);
  assign t[304] = (x[37]);
  assign t[305] = (x[37]);
  assign t[306] = (x[40]);
  assign t[307] = (x[40]);
  assign t[308] = (x[43]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = (x[46]);
  assign t[311] = (x[46]);
  assign t[312] = (x[53]);
  assign t[313] = (x[53]);
  assign t[314] = (x[56]);
  assign t[315] = (x[56]);
  assign t[316] = (x[59]);
  assign t[317] = (x[59]);
  assign t[318] = (x[62]);
  assign t[319] = (x[62]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[65]);
  assign t[321] = (x[65]);
  assign t[322] = (x[72]);
  assign t[323] = (x[72]);
  assign t[324] = (x[79]);
  assign t[325] = (x[79]);
  assign t[326] = (x[84]);
  assign t[327] = (x[84]);
  assign t[328] = (x[87]);
  assign t[329] = (x[87]);
  assign t[32] = ~(t[157]);
  assign t[330] = (x[90]);
  assign t[331] = (x[90]);
  assign t[332] = (x[99]);
  assign t[333] = (x[99]);
  assign t[33] = ~(t[158]);
  assign t[34] = ~(t[159]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[160] ^ t[61];
  assign t[39] = t[62] ^ t[63];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~t[4];
  assign t[41] = t[64];
  assign t[42] = ~(t[22] ^ t[65]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[68]);
  assign t[45] = t[154] ^ t[69];
  assign t[46] = t[155] ^ t[70];
  assign t[47] = t[71] & t[72];
  assign t[48] = t[73] & t[74];
  assign t[49] = ~(t[47] ^ t[75]);
  assign t[4] = t[8] ? t[9] : t[152];
  assign t[50] = t[76] ^ t[77];
  assign t[51] = ~(t[78] & t[79]);
  assign t[52] = t[80] ^ t[161];
  assign t[53] = ~(t[156]);
  assign t[54] = t[81] & t[80];
  assign t[55] = ~(t[160]);
  assign t[56] = ~(t[82] & t[162]);
  assign t[57] = t[44] ? t[83] : t[163];
  assign t[58] = t[44] ? t[84] : t[164];
  assign t[59] = t[85] ^ t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[87] & t[88];
  assign t[61] = t[89] ? t[90] : t[165];
  assign t[62] = t[91] ^ t[92];
  assign t[63] = t[93] & t[94];
  assign t[64] = t[8] ? t[95] : t[166];
  assign t[65] = t[96] ^ t[97];
  assign t[66] = t[41] ^ t[98];
  assign t[67] = t[99];
  assign t[68] = ~(t[8]);
  assign t[69] = t[100] ? x[50] : x[49];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[100] ? x[52] : x[51];
  assign t[71] = ~(t[77]);
  assign t[72] = ~(t[101]);
  assign t[73] = ~(t[24]);
  assign t[74] = t[44] ? t[102] : t[167];
  assign t[75] = t[13] ^ t[101];
  assign t[76] = t[101] ^ t[25];
  assign t[77] = t[74] ^ t[24];
  assign t[78] = ~(t[81] | t[80]);
  assign t[79] = ~(t[103] | t[53]);
  assign t[7] = t[13] ^ t[14];
  assign t[80] = ~(t[168]);
  assign t[81] = ~(t[161]);
  assign t[82] = ~(t[169]);
  assign t[83] = t[163] ^ t[104];
  assign t[84] = t[164] ^ t[105];
  assign t[85] = t[106] & t[107];
  assign t[86] = t[108] & t[109];
  assign t[87] = ~(t[85] ^ t[110]);
  assign t[88] = t[111] ^ t[112];
  assign t[89] = ~(t[68]);
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[165] ^ t[113];
  assign t[91] = t[114] & t[115];
  assign t[92] = t[116] & t[117];
  assign t[93] = ~(t[118] ^ t[62]);
  assign t[94] = t[119] ^ t[117];
  assign t[95] = t[166] ^ t[120];
  assign t[96] = t[121] & t[122];
  assign t[97] = t[123] & t[67];
  assign t[98] = t[124];
  assign t[99] = t[8] ? t[125] : t[170];
  assign t[9] = t[152] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind31(x, y);
 input [111:0] x;
 output y;

 wire [333:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[126]);
  assign t[101] = t[44] ? t[127] : t[171];
  assign t[102] = t[167] ^ t[128];
  assign t[103] = ~(t[153]);
  assign t[104] = t[129] ? x[69] : x[68];
  assign t[105] = t[129] ? x[71] : x[70];
  assign t[106] = ~(t[112]);
  assign t[107] = ~(t[130]);
  assign t[108] = ~(t[57]);
  assign t[109] = t[44] ? t[131] : t[172];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[36] ^ t[130];
  assign t[111] = t[130] ^ t[58];
  assign t[112] = t[109] ^ t[57];
  assign t[113] = t[132] ? x[76] : x[75];
  assign t[114] = ~(t[133]);
  assign t[115] = ~(t[134]);
  assign t[116] = ~(t[135]);
  assign t[117] = t[169] ^ t[136];
  assign t[118] = t[134] ^ t[135];
  assign t[119] = t[135] ^ t[38];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[132] ? x[78] : x[77];
  assign t[121] = ~(t[137]);
  assign t[122] = ~(t[40]);
  assign t[123] = ~(t[41]);
  assign t[124] = t[8] ? t[138] : t[173];
  assign t[125] = t[170] ^ t[139];
  assign t[126] = ~(t[31]);
  assign t[127] = t[171] ^ t[140];
  assign t[128] = t[100] ? x[83] : x[82];
  assign t[129] = ~(t[126]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[44] ? t[141] : t[174];
  assign t[131] = t[172] ^ t[142];
  assign t[132] = ~(t[126]);
  assign t[133] = t[117] ^ t[135];
  assign t[134] = t[8] ? t[143] : t[175];
  assign t[135] = t[159] ^ t[144];
  assign t[136] = t[8] ? t[145] : t[176];
  assign t[137] = t[67] ^ t[41];
  assign t[138] = t[173] ^ t[146];
  assign t[139] = t[132] ? x[94] : x[93];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[100] ? x[96] : x[95];
  assign t[141] = t[174] ^ t[147];
  assign t[142] = t[129] ? x[98] : x[97];
  assign t[143] = t[175] ^ t[148];
  assign t[144] = t[8] ? t[149] : t[177];
  assign t[145] = t[176] ^ t[150];
  assign t[146] = t[31] ? x[103] : x[102];
  assign t[147] = t[129] ? x[105] : x[104];
  assign t[148] = t[100] ? x[107] : x[106];
  assign t[149] = t[177] ^ t[151];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[31] ? x[109] : x[108];
  assign t[151] = t[100] ? x[111] : x[110];
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[153] | t[30];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = t[204] ^ x[4];
  assign t[179] = t[205] ^ x[7];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[206] ^ x[12];
  assign t[181] = t[207] ^ x[15];
  assign t[182] = t[208] ^ x[18];
  assign t[183] = t[209] ^ x[21];
  assign t[184] = t[210] ^ x[24];
  assign t[185] = t[211] ^ x[27];
  assign t[186] = t[212] ^ x[30];
  assign t[187] = t[213] ^ x[33];
  assign t[188] = t[214] ^ x[36];
  assign t[189] = t[215] ^ x[39];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[216] ^ x[42];
  assign t[191] = t[217] ^ x[45];
  assign t[192] = t[218] ^ x[48];
  assign t[193] = t[219] ^ x[55];
  assign t[194] = t[220] ^ x[58];
  assign t[195] = t[221] ^ x[61];
  assign t[196] = t[222] ^ x[64];
  assign t[197] = t[223] ^ x[67];
  assign t[198] = t[224] ^ x[74];
  assign t[199] = t[225] ^ x[81];
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[86];
  assign t[201] = t[227] ^ x[89];
  assign t[202] = t[228] ^ x[92];
  assign t[203] = t[229] ^ x[101];
  assign t[204] = (t[230] & ~t[231]);
  assign t[205] = (t[232] & ~t[233]);
  assign t[206] = (t[234] & ~t[235]);
  assign t[207] = (t[236] & ~t[237]);
  assign t[208] = (t[238] & ~t[239]);
  assign t[209] = (t[240] & ~t[241]);
  assign t[20] = t[36] ^ t[37];
  assign t[210] = (t[242] & ~t[243]);
  assign t[211] = (t[244] & ~t[245]);
  assign t[212] = (t[246] & ~t[247]);
  assign t[213] = (t[248] & ~t[249]);
  assign t[214] = (t[250] & ~t[251]);
  assign t[215] = (t[252] & ~t[253]);
  assign t[216] = (t[254] & ~t[255]);
  assign t[217] = (t[256] & ~t[257]);
  assign t[218] = (t[258] & ~t[259]);
  assign t[219] = (t[260] & ~t[261]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = (t[262] & ~t[263]);
  assign t[221] = (t[264] & ~t[265]);
  assign t[222] = (t[266] & ~t[267]);
  assign t[223] = (t[268] & ~t[269]);
  assign t[224] = (t[270] & ~t[271]);
  assign t[225] = (t[272] & ~t[273]);
  assign t[226] = (t[274] & ~t[275]);
  assign t[227] = (t[276] & ~t[277]);
  assign t[228] = (t[278] & ~t[279]);
  assign t[229] = (t[280] & ~t[281]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[282] ^ x[4];
  assign t[231] = t[283] ^ x[3];
  assign t[232] = t[284] ^ x[7];
  assign t[233] = t[285] ^ x[6];
  assign t[234] = t[286] ^ x[12];
  assign t[235] = t[287] ^ x[11];
  assign t[236] = t[288] ^ x[15];
  assign t[237] = t[289] ^ x[14];
  assign t[238] = t[290] ^ x[18];
  assign t[239] = t[291] ^ x[17];
  assign t[23] = t[42] & t[43];
  assign t[240] = t[292] ^ x[21];
  assign t[241] = t[293] ^ x[20];
  assign t[242] = t[294] ^ x[24];
  assign t[243] = t[295] ^ x[23];
  assign t[244] = t[296] ^ x[27];
  assign t[245] = t[297] ^ x[26];
  assign t[246] = t[298] ^ x[30];
  assign t[247] = t[299] ^ x[29];
  assign t[248] = t[300] ^ x[33];
  assign t[249] = t[301] ^ x[32];
  assign t[24] = t[44] ? t[45] : t[154];
  assign t[250] = t[302] ^ x[36];
  assign t[251] = t[303] ^ x[35];
  assign t[252] = t[304] ^ x[39];
  assign t[253] = t[305] ^ x[38];
  assign t[254] = t[306] ^ x[42];
  assign t[255] = t[307] ^ x[41];
  assign t[256] = t[308] ^ x[45];
  assign t[257] = t[309] ^ x[44];
  assign t[258] = t[310] ^ x[48];
  assign t[259] = t[311] ^ x[47];
  assign t[25] = t[44] ? t[46] : t[155];
  assign t[260] = t[312] ^ x[55];
  assign t[261] = t[313] ^ x[54];
  assign t[262] = t[314] ^ x[58];
  assign t[263] = t[315] ^ x[57];
  assign t[264] = t[316] ^ x[61];
  assign t[265] = t[317] ^ x[60];
  assign t[266] = t[318] ^ x[64];
  assign t[267] = t[319] ^ x[63];
  assign t[268] = t[320] ^ x[67];
  assign t[269] = t[321] ^ x[66];
  assign t[26] = t[47] ^ t[48];
  assign t[270] = t[322] ^ x[74];
  assign t[271] = t[323] ^ x[73];
  assign t[272] = t[324] ^ x[81];
  assign t[273] = t[325] ^ x[80];
  assign t[274] = t[326] ^ x[86];
  assign t[275] = t[327] ^ x[85];
  assign t[276] = t[328] ^ x[89];
  assign t[277] = t[329] ^ x[88];
  assign t[278] = t[330] ^ x[92];
  assign t[279] = t[331] ^ x[91];
  assign t[27] = t[49] & t[50];
  assign t[280] = t[332] ^ x[101];
  assign t[281] = t[333] ^ x[100];
  assign t[282] = (x[2]);
  assign t[283] = (x[2]);
  assign t[284] = (x[5]);
  assign t[285] = (x[5]);
  assign t[286] = (x[10]);
  assign t[287] = (x[10]);
  assign t[288] = (x[13]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = (x[16]);
  assign t[291] = (x[16]);
  assign t[292] = (x[19]);
  assign t[293] = (x[19]);
  assign t[294] = (x[22]);
  assign t[295] = (x[22]);
  assign t[296] = (x[25]);
  assign t[297] = (x[25]);
  assign t[298] = (x[28]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[156] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[31]);
  assign t[301] = (x[31]);
  assign t[302] = (x[34]);
  assign t[303] = (x[34]);
  assign t[304] = (x[37]);
  assign t[305] = (x[37]);
  assign t[306] = (x[40]);
  assign t[307] = (x[40]);
  assign t[308] = (x[43]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = (x[46]);
  assign t[311] = (x[46]);
  assign t[312] = (x[53]);
  assign t[313] = (x[53]);
  assign t[314] = (x[56]);
  assign t[315] = (x[56]);
  assign t[316] = (x[59]);
  assign t[317] = (x[59]);
  assign t[318] = (x[62]);
  assign t[319] = (x[62]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[65]);
  assign t[321] = (x[65]);
  assign t[322] = (x[72]);
  assign t[323] = (x[72]);
  assign t[324] = (x[79]);
  assign t[325] = (x[79]);
  assign t[326] = (x[84]);
  assign t[327] = (x[84]);
  assign t[328] = (x[87]);
  assign t[329] = (x[87]);
  assign t[32] = ~(t[157]);
  assign t[330] = (x[90]);
  assign t[331] = (x[90]);
  assign t[332] = (x[99]);
  assign t[333] = (x[99]);
  assign t[33] = ~(t[158]);
  assign t[34] = ~(t[159]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[160] ^ t[61];
  assign t[39] = t[62] ^ t[63];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~t[4];
  assign t[41] = t[64];
  assign t[42] = ~(t[22] ^ t[65]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[68]);
  assign t[45] = t[154] ^ t[69];
  assign t[46] = t[155] ^ t[70];
  assign t[47] = t[71] & t[72];
  assign t[48] = t[73] & t[74];
  assign t[49] = ~(t[47] ^ t[75]);
  assign t[4] = t[8] ? t[9] : t[152];
  assign t[50] = t[76] ^ t[77];
  assign t[51] = ~(t[78] & t[79]);
  assign t[52] = t[80] ^ t[161];
  assign t[53] = ~(t[156]);
  assign t[54] = t[81] & t[80];
  assign t[55] = ~(t[160]);
  assign t[56] = ~(t[82] & t[162]);
  assign t[57] = t[44] ? t[83] : t[163];
  assign t[58] = t[44] ? t[84] : t[164];
  assign t[59] = t[85] ^ t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[87] & t[88];
  assign t[61] = t[89] ? t[90] : t[165];
  assign t[62] = t[91] ^ t[92];
  assign t[63] = t[93] & t[94];
  assign t[64] = t[8] ? t[95] : t[166];
  assign t[65] = t[96] ^ t[97];
  assign t[66] = t[41] ^ t[98];
  assign t[67] = t[99];
  assign t[68] = ~(t[8]);
  assign t[69] = t[100] ? x[50] : x[49];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[100] ? x[52] : x[51];
  assign t[71] = ~(t[77]);
  assign t[72] = ~(t[101]);
  assign t[73] = ~(t[24]);
  assign t[74] = t[44] ? t[102] : t[167];
  assign t[75] = t[13] ^ t[101];
  assign t[76] = t[101] ^ t[25];
  assign t[77] = t[74] ^ t[24];
  assign t[78] = ~(t[81] | t[80]);
  assign t[79] = ~(t[103] | t[53]);
  assign t[7] = t[13] ^ t[14];
  assign t[80] = ~(t[168]);
  assign t[81] = ~(t[161]);
  assign t[82] = ~(t[169]);
  assign t[83] = t[163] ^ t[104];
  assign t[84] = t[164] ^ t[105];
  assign t[85] = t[106] & t[107];
  assign t[86] = t[108] & t[109];
  assign t[87] = ~(t[85] ^ t[110]);
  assign t[88] = t[111] ^ t[112];
  assign t[89] = ~(t[68]);
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[165] ^ t[113];
  assign t[91] = t[114] & t[115];
  assign t[92] = t[116] & t[117];
  assign t[93] = ~(t[118] ^ t[62]);
  assign t[94] = t[119] ^ t[117];
  assign t[95] = t[166] ^ t[120];
  assign t[96] = t[121] & t[122];
  assign t[97] = t[123] & t[67];
  assign t[98] = t[124];
  assign t[99] = t[8] ? t[125] : t[170];
  assign t[9] = t[152] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind32(x, y);
 input [111:0] x;
 output y;

 wire [323:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[44] ? t[119] : t[158];
  assign t[101] = t[117] ^ t[118];
  assign t[102] = t[118] ^ t[25];
  assign t[103] = ~(t[120] & t[121]);
  assign t[104] = t[122] ^ t[159];
  assign t[105] = ~(t[156]);
  assign t[106] = t[123] & t[122];
  assign t[107] = t[28] ? x[69] : x[68];
  assign t[108] = t[8] ? t[124] : t[160];
  assign t[109] = t[8] ? t[125] : t[161];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[50]);
  assign t[111] = t[110] ? x[77] : x[76];
  assign t[112] = t[93] ^ t[114];
  assign t[113] = t[126];
  assign t[114] = ~t[127];
  assign t[115] = t[27] ? t[128] : t[162];
  assign t[116] = t[100] ^ t[118];
  assign t[117] = t[44] ? t[129] : t[163];
  assign t[118] = t[44] ? t[130] : t[164];
  assign t[119] = t[158] ^ t[131];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[123] | t[122]);
  assign t[121] = ~(t[132] | t[105]);
  assign t[122] = ~(t[165]);
  assign t[123] = ~(t[159]);
  assign t[124] = t[160] ^ t[133];
  assign t[125] = t[161] ^ t[134];
  assign t[126] = t[44] ? t[135] : t[166];
  assign t[127] = t[44] ? t[136] : t[167];
  assign t[128] = t[162] ^ t[137];
  assign t[129] = t[163] ^ t[138];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[164] ^ t[139];
  assign t[131] = t[96] ? x[97] : x[96];
  assign t[132] = ~(t[152]);
  assign t[133] = t[28] ? x[99] : x[98];
  assign t[134] = t[28] ? x[101] : x[100];
  assign t[135] = t[166] ^ t[140];
  assign t[136] = t[167] ^ t[141];
  assign t[137] = t[96] ? x[103] : x[102];
  assign t[138] = t[96] ? x[105] : x[104];
  assign t[139] = t[96] ? x[107] : x[106];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[96] ? x[109] : x[108];
  assign t[141] = t[96] ? x[111] : x[110];
  assign t[142] = (t[168]);
  assign t[143] = (t[169]);
  assign t[144] = (t[170]);
  assign t[145] = (t[171]);
  assign t[146] = (t[172]);
  assign t[147] = (t[173]);
  assign t[148] = (t[174]);
  assign t[149] = (t[175]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = (t[176]);
  assign t[151] = (t[177]);
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = t[194] ^ x[4];
  assign t[169] = t[195] ^ x[9];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[196] ^ x[12];
  assign t[171] = t[197] ^ x[15];
  assign t[172] = t[198] ^ x[18];
  assign t[173] = t[199] ^ x[21];
  assign t[174] = t[200] ^ x[24];
  assign t[175] = t[201] ^ x[27];
  assign t[176] = t[202] ^ x[30];
  assign t[177] = t[203] ^ x[33];
  assign t[178] = t[204] ^ x[36];
  assign t[179] = t[205] ^ x[39];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[42];
  assign t[181] = t[207] ^ x[45];
  assign t[182] = t[208] ^ x[50];
  assign t[183] = t[209] ^ x[53];
  assign t[184] = t[210] ^ x[64];
  assign t[185] = t[211] ^ x[67];
  assign t[186] = t[212] ^ x[72];
  assign t[187] = t[213] ^ x[75];
  assign t[188] = t[214] ^ x[80];
  assign t[189] = t[215] ^ x[83];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[86];
  assign t[191] = t[217] ^ x[89];
  assign t[192] = t[218] ^ x[92];
  assign t[193] = t[219] ^ x[95];
  assign t[194] = (t[220] & ~t[221]);
  assign t[195] = (t[222] & ~t[223]);
  assign t[196] = (t[224] & ~t[225]);
  assign t[197] = (t[226] & ~t[227]);
  assign t[198] = (t[228] & ~t[229]);
  assign t[199] = (t[230] & ~t[231]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[232] & ~t[233]);
  assign t[201] = (t[234] & ~t[235]);
  assign t[202] = (t[236] & ~t[237]);
  assign t[203] = (t[238] & ~t[239]);
  assign t[204] = (t[240] & ~t[241]);
  assign t[205] = (t[242] & ~t[243]);
  assign t[206] = (t[244] & ~t[245]);
  assign t[207] = (t[246] & ~t[247]);
  assign t[208] = (t[248] & ~t[249]);
  assign t[209] = (t[250] & ~t[251]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[252] & ~t[253]);
  assign t[211] = (t[254] & ~t[255]);
  assign t[212] = (t[256] & ~t[257]);
  assign t[213] = (t[258] & ~t[259]);
  assign t[214] = (t[260] & ~t[261]);
  assign t[215] = (t[262] & ~t[263]);
  assign t[216] = (t[264] & ~t[265]);
  assign t[217] = (t[266] & ~t[267]);
  assign t[218] = (t[268] & ~t[269]);
  assign t[219] = (t[270] & ~t[271]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[272] ^ x[4];
  assign t[221] = t[273] ^ x[3];
  assign t[222] = t[274] ^ x[9];
  assign t[223] = t[275] ^ x[8];
  assign t[224] = t[276] ^ x[12];
  assign t[225] = t[277] ^ x[11];
  assign t[226] = t[278] ^ x[15];
  assign t[227] = t[279] ^ x[14];
  assign t[228] = t[280] ^ x[18];
  assign t[229] = t[281] ^ x[17];
  assign t[22] = t[39] & t[40];
  assign t[230] = t[282] ^ x[21];
  assign t[231] = t[283] ^ x[20];
  assign t[232] = t[284] ^ x[24];
  assign t[233] = t[285] ^ x[23];
  assign t[234] = t[286] ^ x[27];
  assign t[235] = t[287] ^ x[26];
  assign t[236] = t[288] ^ x[30];
  assign t[237] = t[289] ^ x[29];
  assign t[238] = t[290] ^ x[33];
  assign t[239] = t[291] ^ x[32];
  assign t[23] = ~t[41];
  assign t[240] = t[292] ^ x[36];
  assign t[241] = t[293] ^ x[35];
  assign t[242] = t[294] ^ x[39];
  assign t[243] = t[295] ^ x[38];
  assign t[244] = t[296] ^ x[42];
  assign t[245] = t[297] ^ x[41];
  assign t[246] = t[298] ^ x[45];
  assign t[247] = t[299] ^ x[44];
  assign t[248] = t[300] ^ x[50];
  assign t[249] = t[301] ^ x[49];
  assign t[24] = t[42] ^ t[43];
  assign t[250] = t[302] ^ x[53];
  assign t[251] = t[303] ^ x[52];
  assign t[252] = t[304] ^ x[64];
  assign t[253] = t[305] ^ x[63];
  assign t[254] = t[306] ^ x[67];
  assign t[255] = t[307] ^ x[66];
  assign t[256] = t[308] ^ x[72];
  assign t[257] = t[309] ^ x[71];
  assign t[258] = t[310] ^ x[75];
  assign t[259] = t[311] ^ x[74];
  assign t[25] = t[44] ? t[45] : t[143];
  assign t[260] = t[312] ^ x[80];
  assign t[261] = t[313] ^ x[79];
  assign t[262] = t[314] ^ x[83];
  assign t[263] = t[315] ^ x[82];
  assign t[264] = t[316] ^ x[86];
  assign t[265] = t[317] ^ x[85];
  assign t[266] = t[318] ^ x[89];
  assign t[267] = t[319] ^ x[88];
  assign t[268] = t[320] ^ x[92];
  assign t[269] = t[321] ^ x[91];
  assign t[26] = t[46] ^ t[47];
  assign t[270] = t[322] ^ x[95];
  assign t[271] = t[323] ^ x[94];
  assign t[272] = (x[2]);
  assign t[273] = (x[2]);
  assign t[274] = (x[7]);
  assign t[275] = (x[7]);
  assign t[276] = (x[10]);
  assign t[277] = (x[10]);
  assign t[278] = (x[13]);
  assign t[279] = (x[13]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = (x[16]);
  assign t[281] = (x[16]);
  assign t[282] = (x[19]);
  assign t[283] = (x[19]);
  assign t[284] = (x[22]);
  assign t[285] = (x[22]);
  assign t[286] = (x[25]);
  assign t[287] = (x[25]);
  assign t[288] = (x[28]);
  assign t[289] = (x[28]);
  assign t[28] = ~(t[50]);
  assign t[290] = (x[31]);
  assign t[291] = (x[31]);
  assign t[292] = (x[34]);
  assign t[293] = (x[34]);
  assign t[294] = (x[37]);
  assign t[295] = (x[37]);
  assign t[296] = (x[40]);
  assign t[297] = (x[40]);
  assign t[298] = (x[43]);
  assign t[299] = (x[43]);
  assign t[29] = ~(t[144]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[48]);
  assign t[301] = (x[48]);
  assign t[302] = (x[51]);
  assign t[303] = (x[51]);
  assign t[304] = (x[62]);
  assign t[305] = (x[62]);
  assign t[306] = (x[65]);
  assign t[307] = (x[65]);
  assign t[308] = (x[70]);
  assign t[309] = (x[70]);
  assign t[30] = ~(t[145]);
  assign t[310] = (x[73]);
  assign t[311] = (x[73]);
  assign t[312] = (x[78]);
  assign t[313] = (x[78]);
  assign t[314] = (x[81]);
  assign t[315] = (x[81]);
  assign t[316] = (x[84]);
  assign t[317] = (x[84]);
  assign t[318] = (x[87]);
  assign t[319] = (x[87]);
  assign t[31] = ~(t[146]);
  assign t[320] = (x[90]);
  assign t[321] = (x[90]);
  assign t[322] = (x[93]);
  assign t[323] = (x[93]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[33] = t[144] ^ t[53];
  assign t[34] = t[147] ^ t[4];
  assign t[35] = t[54] ^ t[55];
  assign t[36] = t[56] & t[57];
  assign t[37] = t[27] ? t[58] : t[148];
  assign t[38] = t[27] ? t[59] : t[149];
  assign t[39] = ~(t[60]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[27] ? t[61] : t[150];
  assign t[41] = t[44] ? t[62] : t[151];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[65] & t[66];
  assign t[44] = ~(t[15]);
  assign t[45] = t[143] ^ t[67];
  assign t[46] = t[68] ^ t[69];
  assign t[47] = t[70] & t[71];
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = t[152] | t[74];
  assign t[4] = t[8] ? t[9] : t[142];
  assign t[50] = ~(t[75]);
  assign t[51] = ~(t[153]);
  assign t[52] = ~(t[76] & t[147]);
  assign t[53] = t[8] ? t[77] : t[154];
  assign t[54] = t[78] & t[79];
  assign t[55] = t[80] & t[81];
  assign t[56] = ~(t[54] ^ t[82]);
  assign t[57] = t[83] ^ t[84];
  assign t[58] = t[148] ^ t[85];
  assign t[59] = t[149] ^ t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[27] ? t[87] : t[155];
  assign t[61] = t[150] ^ t[88];
  assign t[62] = t[151] ^ t[89];
  assign t[63] = t[90] & t[91];
  assign t[64] = t[92] & t[93];
  assign t[65] = ~(t[94] ^ t[42]);
  assign t[66] = t[95] ^ t[93];
  assign t[67] = t[96] ? x[47] : x[46];
  assign t[68] = t[97] & t[98];
  assign t[69] = t[99] & t[100];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[101] ^ t[46]);
  assign t[71] = t[102] ^ t[100];
  assign t[72] = ~(t[74] & t[103]);
  assign t[73] = ~(t[156] ^ t[104]);
  assign t[74] = ~(t[105] & t[106]);
  assign t[75] = ~(t[49]);
  assign t[76] = ~(t[157]);
  assign t[77] = t[154] ^ t[107];
  assign t[78] = ~(t[84]);
  assign t[79] = ~(t[108]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[33]);
  assign t[81] = t[145] ^ t[109];
  assign t[82] = t[19] ^ t[108];
  assign t[83] = t[108] ^ t[34];
  assign t[84] = t[81] ^ t[33];
  assign t[85] = t[110] ? x[55] : x[54];
  assign t[86] = t[75] ? x[57] : x[56];
  assign t[87] = t[155] ^ t[111];
  assign t[88] = t[75] ? x[59] : x[58];
  assign t[89] = t[96] ? x[61] : x[60];
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[112]);
  assign t[91] = ~(t[113]);
  assign t[92] = ~(t[114]);
  assign t[93] = t[115];
  assign t[94] = t[113] ^ t[114];
  assign t[95] = t[114] ^ t[23];
  assign t[96] = ~(t[50]);
  assign t[97] = ~(t[116]);
  assign t[98] = ~(t[117]);
  assign t[99] = ~(t[118]);
  assign t[9] = t[142] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind33(x, y);
 input [111:0] x;
 output y;

 wire [323:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[44] ? t[119] : t[158];
  assign t[101] = t[117] ^ t[118];
  assign t[102] = t[118] ^ t[25];
  assign t[103] = ~(t[120] & t[121]);
  assign t[104] = t[122] ^ t[159];
  assign t[105] = ~(t[156]);
  assign t[106] = t[123] & t[122];
  assign t[107] = t[28] ? x[69] : x[68];
  assign t[108] = t[8] ? t[124] : t[160];
  assign t[109] = t[8] ? t[125] : t[161];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[50]);
  assign t[111] = t[110] ? x[77] : x[76];
  assign t[112] = t[93] ^ t[114];
  assign t[113] = t[126];
  assign t[114] = ~t[127];
  assign t[115] = t[27] ? t[128] : t[162];
  assign t[116] = t[100] ^ t[118];
  assign t[117] = t[44] ? t[129] : t[163];
  assign t[118] = t[44] ? t[130] : t[164];
  assign t[119] = t[158] ^ t[131];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[123] | t[122]);
  assign t[121] = ~(t[132] | t[105]);
  assign t[122] = ~(t[165]);
  assign t[123] = ~(t[159]);
  assign t[124] = t[160] ^ t[133];
  assign t[125] = t[161] ^ t[134];
  assign t[126] = t[44] ? t[135] : t[166];
  assign t[127] = t[44] ? t[136] : t[167];
  assign t[128] = t[162] ^ t[137];
  assign t[129] = t[163] ^ t[138];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[164] ^ t[139];
  assign t[131] = t[96] ? x[97] : x[96];
  assign t[132] = ~(t[152]);
  assign t[133] = t[28] ? x[99] : x[98];
  assign t[134] = t[28] ? x[101] : x[100];
  assign t[135] = t[166] ^ t[140];
  assign t[136] = t[167] ^ t[141];
  assign t[137] = t[96] ? x[103] : x[102];
  assign t[138] = t[96] ? x[105] : x[104];
  assign t[139] = t[96] ? x[107] : x[106];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[96] ? x[109] : x[108];
  assign t[141] = t[96] ? x[111] : x[110];
  assign t[142] = (t[168]);
  assign t[143] = (t[169]);
  assign t[144] = (t[170]);
  assign t[145] = (t[171]);
  assign t[146] = (t[172]);
  assign t[147] = (t[173]);
  assign t[148] = (t[174]);
  assign t[149] = (t[175]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = (t[176]);
  assign t[151] = (t[177]);
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = t[194] ^ x[4];
  assign t[169] = t[195] ^ x[9];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[196] ^ x[12];
  assign t[171] = t[197] ^ x[15];
  assign t[172] = t[198] ^ x[18];
  assign t[173] = t[199] ^ x[21];
  assign t[174] = t[200] ^ x[24];
  assign t[175] = t[201] ^ x[27];
  assign t[176] = t[202] ^ x[30];
  assign t[177] = t[203] ^ x[33];
  assign t[178] = t[204] ^ x[36];
  assign t[179] = t[205] ^ x[39];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[42];
  assign t[181] = t[207] ^ x[45];
  assign t[182] = t[208] ^ x[50];
  assign t[183] = t[209] ^ x[53];
  assign t[184] = t[210] ^ x[64];
  assign t[185] = t[211] ^ x[67];
  assign t[186] = t[212] ^ x[72];
  assign t[187] = t[213] ^ x[75];
  assign t[188] = t[214] ^ x[80];
  assign t[189] = t[215] ^ x[83];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[86];
  assign t[191] = t[217] ^ x[89];
  assign t[192] = t[218] ^ x[92];
  assign t[193] = t[219] ^ x[95];
  assign t[194] = (t[220] & ~t[221]);
  assign t[195] = (t[222] & ~t[223]);
  assign t[196] = (t[224] & ~t[225]);
  assign t[197] = (t[226] & ~t[227]);
  assign t[198] = (t[228] & ~t[229]);
  assign t[199] = (t[230] & ~t[231]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[232] & ~t[233]);
  assign t[201] = (t[234] & ~t[235]);
  assign t[202] = (t[236] & ~t[237]);
  assign t[203] = (t[238] & ~t[239]);
  assign t[204] = (t[240] & ~t[241]);
  assign t[205] = (t[242] & ~t[243]);
  assign t[206] = (t[244] & ~t[245]);
  assign t[207] = (t[246] & ~t[247]);
  assign t[208] = (t[248] & ~t[249]);
  assign t[209] = (t[250] & ~t[251]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[252] & ~t[253]);
  assign t[211] = (t[254] & ~t[255]);
  assign t[212] = (t[256] & ~t[257]);
  assign t[213] = (t[258] & ~t[259]);
  assign t[214] = (t[260] & ~t[261]);
  assign t[215] = (t[262] & ~t[263]);
  assign t[216] = (t[264] & ~t[265]);
  assign t[217] = (t[266] & ~t[267]);
  assign t[218] = (t[268] & ~t[269]);
  assign t[219] = (t[270] & ~t[271]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[272] ^ x[4];
  assign t[221] = t[273] ^ x[3];
  assign t[222] = t[274] ^ x[9];
  assign t[223] = t[275] ^ x[8];
  assign t[224] = t[276] ^ x[12];
  assign t[225] = t[277] ^ x[11];
  assign t[226] = t[278] ^ x[15];
  assign t[227] = t[279] ^ x[14];
  assign t[228] = t[280] ^ x[18];
  assign t[229] = t[281] ^ x[17];
  assign t[22] = t[39] & t[40];
  assign t[230] = t[282] ^ x[21];
  assign t[231] = t[283] ^ x[20];
  assign t[232] = t[284] ^ x[24];
  assign t[233] = t[285] ^ x[23];
  assign t[234] = t[286] ^ x[27];
  assign t[235] = t[287] ^ x[26];
  assign t[236] = t[288] ^ x[30];
  assign t[237] = t[289] ^ x[29];
  assign t[238] = t[290] ^ x[33];
  assign t[239] = t[291] ^ x[32];
  assign t[23] = ~t[41];
  assign t[240] = t[292] ^ x[36];
  assign t[241] = t[293] ^ x[35];
  assign t[242] = t[294] ^ x[39];
  assign t[243] = t[295] ^ x[38];
  assign t[244] = t[296] ^ x[42];
  assign t[245] = t[297] ^ x[41];
  assign t[246] = t[298] ^ x[45];
  assign t[247] = t[299] ^ x[44];
  assign t[248] = t[300] ^ x[50];
  assign t[249] = t[301] ^ x[49];
  assign t[24] = t[42] ^ t[43];
  assign t[250] = t[302] ^ x[53];
  assign t[251] = t[303] ^ x[52];
  assign t[252] = t[304] ^ x[64];
  assign t[253] = t[305] ^ x[63];
  assign t[254] = t[306] ^ x[67];
  assign t[255] = t[307] ^ x[66];
  assign t[256] = t[308] ^ x[72];
  assign t[257] = t[309] ^ x[71];
  assign t[258] = t[310] ^ x[75];
  assign t[259] = t[311] ^ x[74];
  assign t[25] = t[44] ? t[45] : t[143];
  assign t[260] = t[312] ^ x[80];
  assign t[261] = t[313] ^ x[79];
  assign t[262] = t[314] ^ x[83];
  assign t[263] = t[315] ^ x[82];
  assign t[264] = t[316] ^ x[86];
  assign t[265] = t[317] ^ x[85];
  assign t[266] = t[318] ^ x[89];
  assign t[267] = t[319] ^ x[88];
  assign t[268] = t[320] ^ x[92];
  assign t[269] = t[321] ^ x[91];
  assign t[26] = t[46] ^ t[47];
  assign t[270] = t[322] ^ x[95];
  assign t[271] = t[323] ^ x[94];
  assign t[272] = (x[2]);
  assign t[273] = (x[2]);
  assign t[274] = (x[7]);
  assign t[275] = (x[7]);
  assign t[276] = (x[10]);
  assign t[277] = (x[10]);
  assign t[278] = (x[13]);
  assign t[279] = (x[13]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = (x[16]);
  assign t[281] = (x[16]);
  assign t[282] = (x[19]);
  assign t[283] = (x[19]);
  assign t[284] = (x[22]);
  assign t[285] = (x[22]);
  assign t[286] = (x[25]);
  assign t[287] = (x[25]);
  assign t[288] = (x[28]);
  assign t[289] = (x[28]);
  assign t[28] = ~(t[50]);
  assign t[290] = (x[31]);
  assign t[291] = (x[31]);
  assign t[292] = (x[34]);
  assign t[293] = (x[34]);
  assign t[294] = (x[37]);
  assign t[295] = (x[37]);
  assign t[296] = (x[40]);
  assign t[297] = (x[40]);
  assign t[298] = (x[43]);
  assign t[299] = (x[43]);
  assign t[29] = ~(t[144]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[48]);
  assign t[301] = (x[48]);
  assign t[302] = (x[51]);
  assign t[303] = (x[51]);
  assign t[304] = (x[62]);
  assign t[305] = (x[62]);
  assign t[306] = (x[65]);
  assign t[307] = (x[65]);
  assign t[308] = (x[70]);
  assign t[309] = (x[70]);
  assign t[30] = ~(t[145]);
  assign t[310] = (x[73]);
  assign t[311] = (x[73]);
  assign t[312] = (x[78]);
  assign t[313] = (x[78]);
  assign t[314] = (x[81]);
  assign t[315] = (x[81]);
  assign t[316] = (x[84]);
  assign t[317] = (x[84]);
  assign t[318] = (x[87]);
  assign t[319] = (x[87]);
  assign t[31] = ~(t[146]);
  assign t[320] = (x[90]);
  assign t[321] = (x[90]);
  assign t[322] = (x[93]);
  assign t[323] = (x[93]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[33] = t[144] ^ t[53];
  assign t[34] = t[147] ^ t[4];
  assign t[35] = t[54] ^ t[55];
  assign t[36] = t[56] & t[57];
  assign t[37] = t[27] ? t[58] : t[148];
  assign t[38] = t[27] ? t[59] : t[149];
  assign t[39] = ~(t[60]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[27] ? t[61] : t[150];
  assign t[41] = t[44] ? t[62] : t[151];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[65] & t[66];
  assign t[44] = ~(t[15]);
  assign t[45] = t[143] ^ t[67];
  assign t[46] = t[68] ^ t[69];
  assign t[47] = t[70] & t[71];
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = t[152] | t[74];
  assign t[4] = t[8] ? t[9] : t[142];
  assign t[50] = ~(t[75]);
  assign t[51] = ~(t[153]);
  assign t[52] = ~(t[76] & t[147]);
  assign t[53] = t[8] ? t[77] : t[154];
  assign t[54] = t[78] & t[79];
  assign t[55] = t[80] & t[81];
  assign t[56] = ~(t[54] ^ t[82]);
  assign t[57] = t[83] ^ t[84];
  assign t[58] = t[148] ^ t[85];
  assign t[59] = t[149] ^ t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[27] ? t[87] : t[155];
  assign t[61] = t[150] ^ t[88];
  assign t[62] = t[151] ^ t[89];
  assign t[63] = t[90] & t[91];
  assign t[64] = t[92] & t[93];
  assign t[65] = ~(t[94] ^ t[42]);
  assign t[66] = t[95] ^ t[93];
  assign t[67] = t[96] ? x[47] : x[46];
  assign t[68] = t[97] & t[98];
  assign t[69] = t[99] & t[100];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[101] ^ t[46]);
  assign t[71] = t[102] ^ t[100];
  assign t[72] = ~(t[74] & t[103]);
  assign t[73] = ~(t[156] ^ t[104]);
  assign t[74] = ~(t[105] & t[106]);
  assign t[75] = ~(t[49]);
  assign t[76] = ~(t[157]);
  assign t[77] = t[154] ^ t[107];
  assign t[78] = ~(t[84]);
  assign t[79] = ~(t[108]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[33]);
  assign t[81] = t[145] ^ t[109];
  assign t[82] = t[19] ^ t[108];
  assign t[83] = t[108] ^ t[34];
  assign t[84] = t[81] ^ t[33];
  assign t[85] = t[110] ? x[55] : x[54];
  assign t[86] = t[75] ? x[57] : x[56];
  assign t[87] = t[155] ^ t[111];
  assign t[88] = t[75] ? x[59] : x[58];
  assign t[89] = t[96] ? x[61] : x[60];
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[112]);
  assign t[91] = ~(t[113]);
  assign t[92] = ~(t[114]);
  assign t[93] = t[115];
  assign t[94] = t[113] ^ t[114];
  assign t[95] = t[114] ^ t[23];
  assign t[96] = ~(t[50]);
  assign t[97] = ~(t[116]);
  assign t[98] = ~(t[117]);
  assign t[99] = ~(t[118]);
  assign t[9] = t[142] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind34(x, y);
 input [111:0] x;
 output y;

 wire [345:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[41]);
  assign t[101] = t[41] ^ t[67];
  assign t[102] = t[67] ^ t[25];
  assign t[103] = ~(t[132] & t[133]);
  assign t[104] = t[134] ^ t[183];
  assign t[105] = ~(t[176]);
  assign t[106] = t[135] & t[134];
  assign t[107] = t[98] ? x[71] : x[70];
  assign t[108] = ~(t[136]);
  assign t[109] = ~(t[56]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[56] ^ t[83];
  assign t[111] = t[83] ^ t[33];
  assign t[112] = t[178] ^ t[137];
  assign t[113] = t[44] ? t[138] : t[184];
  assign t[114] = t[179] ^ t[139];
  assign t[115] = t[180] ^ t[140];
  assign t[116] = t[181] ^ t[141];
  assign t[117] = t[142] ^ t[143];
  assign t[118] = t[86] ^ t[144];
  assign t[119] = t[27] ? t[145] : t[185];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[182] ^ t[146];
  assign t[121] = ~(t[147] ^ t[64]);
  assign t[122] = t[39] ^ t[126];
  assign t[123] = ~(t[129]);
  assign t[124] = ~(t[148]);
  assign t[125] = ~(t[63]);
  assign t[126] = t[167] ^ t[149];
  assign t[127] = t[39] ^ t[148];
  assign t[128] = t[148] ^ t[61];
  assign t[129] = t[126] ^ t[63];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[98] ? x[79] : x[78];
  assign t[131] = t[43] ^ t[67];
  assign t[132] = ~(t[135] | t[134]);
  assign t[133] = ~(t[150] | t[105]);
  assign t[134] = ~(t[186]);
  assign t[135] = ~(t[183]);
  assign t[136] = t[58] ^ t[83];
  assign t[137] = t[98] ? x[84] : x[83];
  assign t[138] = t[184] ^ t[151];
  assign t[139] = t[98] ? x[86] : x[85];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[152] ? x[88] : x[87];
  assign t[141] = t[152] ? x[90] : x[89];
  assign t[142] = t[153] & t[154];
  assign t[143] = t[155] & t[119];
  assign t[144] = t[27] ? t[156] : t[187];
  assign t[145] = t[185] ^ t[157];
  assign t[146] = t[28] ? x[95] : x[94];
  assign t[147] = t[148] ^ t[63];
  assign t[148] = t[8] ? t[158] : t[188];
  assign t[149] = t[8] ? t[159] : t[189];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = ~(t[171]);
  assign t[151] = t[98] ? x[103] : x[102];
  assign t[152] = ~(t[50]);
  assign t[153] = ~(t[160]);
  assign t[154] = ~(t[85]);
  assign t[155] = ~(t[86]);
  assign t[156] = t[187] ^ t[161];
  assign t[157] = t[76] ? x[105] : x[104];
  assign t[158] = t[188] ^ t[162];
  assign t[159] = t[189] ^ t[163];
  assign t[15] = ~(t[27]);
  assign t[160] = t[119] ^ t[86];
  assign t[161] = t[76] ? x[107] : x[106];
  assign t[162] = t[28] ? x[109] : x[108];
  assign t[163] = t[28] ? x[111] : x[110];
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = (t[205]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[206]);
  assign t[181] = (t[207]);
  assign t[182] = (t[208]);
  assign t[183] = (t[209]);
  assign t[184] = (t[210]);
  assign t[185] = (t[211]);
  assign t[186] = (t[212]);
  assign t[187] = (t[213]);
  assign t[188] = (t[214]);
  assign t[189] = (t[215]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[4];
  assign t[191] = t[217] ^ x[9];
  assign t[192] = t[218] ^ x[12];
  assign t[193] = t[219] ^ x[15];
  assign t[194] = t[220] ^ x[18];
  assign t[195] = t[221] ^ x[21];
  assign t[196] = t[222] ^ x[24];
  assign t[197] = t[223] ^ x[27];
  assign t[198] = t[224] ^ x[30];
  assign t[199] = t[225] ^ x[33];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[36];
  assign t[201] = t[227] ^ x[39];
  assign t[202] = t[228] ^ x[44];
  assign t[203] = t[229] ^ x[47];
  assign t[204] = t[230] ^ x[50];
  assign t[205] = t[231] ^ x[53];
  assign t[206] = t[232] ^ x[56];
  assign t[207] = t[233] ^ x[59];
  assign t[208] = t[234] ^ x[62];
  assign t[209] = t[235] ^ x[69];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[236] ^ x[74];
  assign t[211] = t[237] ^ x[77];
  assign t[212] = t[238] ^ x[82];
  assign t[213] = t[239] ^ x[93];
  assign t[214] = t[240] ^ x[98];
  assign t[215] = t[241] ^ x[101];
  assign t[216] = (t[242] & ~t[243]);
  assign t[217] = (t[244] & ~t[245]);
  assign t[218] = (t[246] & ~t[247]);
  assign t[219] = (t[248] & ~t[249]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[250] & ~t[251]);
  assign t[221] = (t[252] & ~t[253]);
  assign t[222] = (t[254] & ~t[255]);
  assign t[223] = (t[256] & ~t[257]);
  assign t[224] = (t[258] & ~t[259]);
  assign t[225] = (t[260] & ~t[261]);
  assign t[226] = (t[262] & ~t[263]);
  assign t[227] = (t[264] & ~t[265]);
  assign t[228] = (t[266] & ~t[267]);
  assign t[229] = (t[268] & ~t[269]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[270] & ~t[271]);
  assign t[231] = (t[272] & ~t[273]);
  assign t[232] = (t[274] & ~t[275]);
  assign t[233] = (t[276] & ~t[277]);
  assign t[234] = (t[278] & ~t[279]);
  assign t[235] = (t[280] & ~t[281]);
  assign t[236] = (t[282] & ~t[283]);
  assign t[237] = (t[284] & ~t[285]);
  assign t[238] = (t[286] & ~t[287]);
  assign t[239] = (t[288] & ~t[289]);
  assign t[23] = t[41] ^ t[25];
  assign t[240] = (t[290] & ~t[291]);
  assign t[241] = (t[292] & ~t[293]);
  assign t[242] = t[294] ^ x[4];
  assign t[243] = t[295] ^ x[3];
  assign t[244] = t[296] ^ x[9];
  assign t[245] = t[297] ^ x[8];
  assign t[246] = t[298] ^ x[12];
  assign t[247] = t[299] ^ x[11];
  assign t[248] = t[300] ^ x[15];
  assign t[249] = t[301] ^ x[14];
  assign t[24] = t[42] & t[43];
  assign t[250] = t[302] ^ x[18];
  assign t[251] = t[303] ^ x[17];
  assign t[252] = t[304] ^ x[21];
  assign t[253] = t[305] ^ x[20];
  assign t[254] = t[306] ^ x[24];
  assign t[255] = t[307] ^ x[23];
  assign t[256] = t[308] ^ x[27];
  assign t[257] = t[309] ^ x[26];
  assign t[258] = t[310] ^ x[30];
  assign t[259] = t[311] ^ x[29];
  assign t[25] = t[44] ? t[45] : t[165];
  assign t[260] = t[312] ^ x[33];
  assign t[261] = t[313] ^ x[32];
  assign t[262] = t[314] ^ x[36];
  assign t[263] = t[315] ^ x[35];
  assign t[264] = t[316] ^ x[39];
  assign t[265] = t[317] ^ x[38];
  assign t[266] = t[318] ^ x[44];
  assign t[267] = t[319] ^ x[43];
  assign t[268] = t[320] ^ x[47];
  assign t[269] = t[321] ^ x[46];
  assign t[26] = t[46] ^ t[47];
  assign t[270] = t[322] ^ x[50];
  assign t[271] = t[323] ^ x[49];
  assign t[272] = t[324] ^ x[53];
  assign t[273] = t[325] ^ x[52];
  assign t[274] = t[326] ^ x[56];
  assign t[275] = t[327] ^ x[55];
  assign t[276] = t[328] ^ x[59];
  assign t[277] = t[329] ^ x[58];
  assign t[278] = t[330] ^ x[62];
  assign t[279] = t[331] ^ x[61];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[332] ^ x[69];
  assign t[281] = t[333] ^ x[68];
  assign t[282] = t[334] ^ x[74];
  assign t[283] = t[335] ^ x[73];
  assign t[284] = t[336] ^ x[77];
  assign t[285] = t[337] ^ x[76];
  assign t[286] = t[338] ^ x[82];
  assign t[287] = t[339] ^ x[81];
  assign t[288] = t[340] ^ x[93];
  assign t[289] = t[341] ^ x[92];
  assign t[28] = ~(t[50]);
  assign t[290] = t[342] ^ x[98];
  assign t[291] = t[343] ^ x[97];
  assign t[292] = t[344] ^ x[101];
  assign t[293] = t[345] ^ x[100];
  assign t[294] = (x[2]);
  assign t[295] = (x[2]);
  assign t[296] = (x[7]);
  assign t[297] = (x[7]);
  assign t[298] = (x[10]);
  assign t[299] = (x[10]);
  assign t[29] = ~(t[166]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[13]);
  assign t[301] = (x[13]);
  assign t[302] = (x[16]);
  assign t[303] = (x[16]);
  assign t[304] = (x[19]);
  assign t[305] = (x[19]);
  assign t[306] = (x[22]);
  assign t[307] = (x[22]);
  assign t[308] = (x[25]);
  assign t[309] = (x[25]);
  assign t[30] = ~(t[167]);
  assign t[310] = (x[28]);
  assign t[311] = (x[28]);
  assign t[312] = (x[31]);
  assign t[313] = (x[31]);
  assign t[314] = (x[34]);
  assign t[315] = (x[34]);
  assign t[316] = (x[37]);
  assign t[317] = (x[37]);
  assign t[318] = (x[42]);
  assign t[319] = (x[42]);
  assign t[31] = ~(t[168]);
  assign t[320] = (x[45]);
  assign t[321] = (x[45]);
  assign t[322] = (x[48]);
  assign t[323] = (x[48]);
  assign t[324] = (x[51]);
  assign t[325] = (x[51]);
  assign t[326] = (x[54]);
  assign t[327] = (x[54]);
  assign t[328] = (x[57]);
  assign t[329] = (x[57]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[60]);
  assign t[331] = (x[60]);
  assign t[332] = (x[67]);
  assign t[333] = (x[67]);
  assign t[334] = (x[72]);
  assign t[335] = (x[72]);
  assign t[336] = (x[75]);
  assign t[337] = (x[75]);
  assign t[338] = (x[80]);
  assign t[339] = (x[80]);
  assign t[33] = ~t[53];
  assign t[340] = (x[91]);
  assign t[341] = (x[91]);
  assign t[342] = (x[96]);
  assign t[343] = (x[96]);
  assign t[344] = (x[99]);
  assign t[345] = (x[99]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] ^ t[33];
  assign t[36] = t[57] & t[58];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[44] ? t[66] : t[169];
  assign t[42] = ~(t[67]);
  assign t[43] = t[44] ? t[68] : t[170];
  assign t[44] = ~(t[15]);
  assign t[45] = t[165] ^ t[69];
  assign t[46] = t[70] ^ t[24];
  assign t[47] = t[71] & t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[171] | t[75];
  assign t[4] = t[8] ? t[9] : t[164];
  assign t[50] = ~(t[76]);
  assign t[51] = ~(t[172]);
  assign t[52] = ~(t[77] & t[173]);
  assign t[53] = t[44] ? t[78] : t[174];
  assign t[54] = t[79] ^ t[36];
  assign t[55] = t[80] & t[81];
  assign t[56] = t[82];
  assign t[57] = ~(t[83]);
  assign t[58] = t[84];
  assign t[59] = t[85] ^ t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[87] & t[88];
  assign t[61] = t[173] ^ t[89];
  assign t[62] = t[64] ^ t[90];
  assign t[63] = t[166] ^ t[4];
  assign t[64] = t[91] ^ t[92];
  assign t[65] = t[93] & t[94];
  assign t[66] = t[169] ^ t[95];
  assign t[67] = t[44] ? t[96] : t[175];
  assign t[68] = t[170] ^ t[97];
  assign t[69] = t[98] ? x[41] : x[40];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[99] & t[100];
  assign t[71] = ~(t[101] ^ t[46]);
  assign t[72] = t[102] ^ t[43];
  assign t[73] = ~(t[75] & t[103]);
  assign t[74] = ~(t[176] ^ t[104]);
  assign t[75] = ~(t[105] & t[106]);
  assign t[76] = ~(t[49]);
  assign t[77] = ~(t[177]);
  assign t[78] = t[174] ^ t[107];
  assign t[79] = t[108] & t[109];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[110] ^ t[54]);
  assign t[81] = t[111] ^ t[58];
  assign t[82] = t[44] ? t[112] : t[178];
  assign t[83] = ~t[113];
  assign t[84] = t[27] ? t[114] : t[179];
  assign t[85] = t[27] ? t[115] : t[180];
  assign t[86] = t[27] ? t[116] : t[181];
  assign t[87] = ~(t[59] ^ t[117]);
  assign t[88] = t[118] ^ t[119];
  assign t[89] = t[8] ? t[120] : t[182];
  assign t[8] = ~(t[15]);
  assign t[90] = t[121] & t[122];
  assign t[91] = t[123] & t[124];
  assign t[92] = t[125] & t[126];
  assign t[93] = ~(t[91] ^ t[127]);
  assign t[94] = t[128] ^ t[129];
  assign t[95] = t[98] ? x[64] : x[63];
  assign t[96] = t[175] ^ t[130];
  assign t[97] = t[98] ? x[66] : x[65];
  assign t[98] = ~(t[50]);
  assign t[99] = ~(t[131]);
  assign t[9] = t[164] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [111:0] x;
 output y;

 wire [345:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[41]);
  assign t[101] = t[41] ^ t[67];
  assign t[102] = t[67] ^ t[25];
  assign t[103] = ~(t[132] & t[133]);
  assign t[104] = t[134] ^ t[183];
  assign t[105] = ~(t[176]);
  assign t[106] = t[135] & t[134];
  assign t[107] = t[98] ? x[71] : x[70];
  assign t[108] = ~(t[136]);
  assign t[109] = ~(t[56]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[56] ^ t[83];
  assign t[111] = t[83] ^ t[33];
  assign t[112] = t[178] ^ t[137];
  assign t[113] = t[44] ? t[138] : t[184];
  assign t[114] = t[179] ^ t[139];
  assign t[115] = t[180] ^ t[140];
  assign t[116] = t[181] ^ t[141];
  assign t[117] = t[142] ^ t[143];
  assign t[118] = t[86] ^ t[144];
  assign t[119] = t[27] ? t[145] : t[185];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[182] ^ t[146];
  assign t[121] = ~(t[147] ^ t[64]);
  assign t[122] = t[39] ^ t[126];
  assign t[123] = ~(t[129]);
  assign t[124] = ~(t[148]);
  assign t[125] = ~(t[63]);
  assign t[126] = t[167] ^ t[149];
  assign t[127] = t[39] ^ t[148];
  assign t[128] = t[148] ^ t[61];
  assign t[129] = t[126] ^ t[63];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[98] ? x[79] : x[78];
  assign t[131] = t[43] ^ t[67];
  assign t[132] = ~(t[135] | t[134]);
  assign t[133] = ~(t[150] | t[105]);
  assign t[134] = ~(t[186]);
  assign t[135] = ~(t[183]);
  assign t[136] = t[58] ^ t[83];
  assign t[137] = t[98] ? x[84] : x[83];
  assign t[138] = t[184] ^ t[151];
  assign t[139] = t[98] ? x[86] : x[85];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[152] ? x[88] : x[87];
  assign t[141] = t[152] ? x[90] : x[89];
  assign t[142] = t[153] & t[154];
  assign t[143] = t[155] & t[119];
  assign t[144] = t[27] ? t[156] : t[187];
  assign t[145] = t[185] ^ t[157];
  assign t[146] = t[28] ? x[95] : x[94];
  assign t[147] = t[148] ^ t[63];
  assign t[148] = t[8] ? t[158] : t[188];
  assign t[149] = t[8] ? t[159] : t[189];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = ~(t[171]);
  assign t[151] = t[98] ? x[103] : x[102];
  assign t[152] = ~(t[50]);
  assign t[153] = ~(t[160]);
  assign t[154] = ~(t[85]);
  assign t[155] = ~(t[86]);
  assign t[156] = t[187] ^ t[161];
  assign t[157] = t[76] ? x[105] : x[104];
  assign t[158] = t[188] ^ t[162];
  assign t[159] = t[189] ^ t[163];
  assign t[15] = ~(t[27]);
  assign t[160] = t[119] ^ t[86];
  assign t[161] = t[76] ? x[107] : x[106];
  assign t[162] = t[28] ? x[109] : x[108];
  assign t[163] = t[28] ? x[111] : x[110];
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = (t[205]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[206]);
  assign t[181] = (t[207]);
  assign t[182] = (t[208]);
  assign t[183] = (t[209]);
  assign t[184] = (t[210]);
  assign t[185] = (t[211]);
  assign t[186] = (t[212]);
  assign t[187] = (t[213]);
  assign t[188] = (t[214]);
  assign t[189] = (t[215]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[4];
  assign t[191] = t[217] ^ x[9];
  assign t[192] = t[218] ^ x[12];
  assign t[193] = t[219] ^ x[15];
  assign t[194] = t[220] ^ x[18];
  assign t[195] = t[221] ^ x[21];
  assign t[196] = t[222] ^ x[24];
  assign t[197] = t[223] ^ x[27];
  assign t[198] = t[224] ^ x[30];
  assign t[199] = t[225] ^ x[33];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[36];
  assign t[201] = t[227] ^ x[39];
  assign t[202] = t[228] ^ x[44];
  assign t[203] = t[229] ^ x[47];
  assign t[204] = t[230] ^ x[50];
  assign t[205] = t[231] ^ x[53];
  assign t[206] = t[232] ^ x[56];
  assign t[207] = t[233] ^ x[59];
  assign t[208] = t[234] ^ x[62];
  assign t[209] = t[235] ^ x[69];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[236] ^ x[74];
  assign t[211] = t[237] ^ x[77];
  assign t[212] = t[238] ^ x[82];
  assign t[213] = t[239] ^ x[93];
  assign t[214] = t[240] ^ x[98];
  assign t[215] = t[241] ^ x[101];
  assign t[216] = (t[242] & ~t[243]);
  assign t[217] = (t[244] & ~t[245]);
  assign t[218] = (t[246] & ~t[247]);
  assign t[219] = (t[248] & ~t[249]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[250] & ~t[251]);
  assign t[221] = (t[252] & ~t[253]);
  assign t[222] = (t[254] & ~t[255]);
  assign t[223] = (t[256] & ~t[257]);
  assign t[224] = (t[258] & ~t[259]);
  assign t[225] = (t[260] & ~t[261]);
  assign t[226] = (t[262] & ~t[263]);
  assign t[227] = (t[264] & ~t[265]);
  assign t[228] = (t[266] & ~t[267]);
  assign t[229] = (t[268] & ~t[269]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[270] & ~t[271]);
  assign t[231] = (t[272] & ~t[273]);
  assign t[232] = (t[274] & ~t[275]);
  assign t[233] = (t[276] & ~t[277]);
  assign t[234] = (t[278] & ~t[279]);
  assign t[235] = (t[280] & ~t[281]);
  assign t[236] = (t[282] & ~t[283]);
  assign t[237] = (t[284] & ~t[285]);
  assign t[238] = (t[286] & ~t[287]);
  assign t[239] = (t[288] & ~t[289]);
  assign t[23] = t[41] ^ t[25];
  assign t[240] = (t[290] & ~t[291]);
  assign t[241] = (t[292] & ~t[293]);
  assign t[242] = t[294] ^ x[4];
  assign t[243] = t[295] ^ x[3];
  assign t[244] = t[296] ^ x[9];
  assign t[245] = t[297] ^ x[8];
  assign t[246] = t[298] ^ x[12];
  assign t[247] = t[299] ^ x[11];
  assign t[248] = t[300] ^ x[15];
  assign t[249] = t[301] ^ x[14];
  assign t[24] = t[42] & t[43];
  assign t[250] = t[302] ^ x[18];
  assign t[251] = t[303] ^ x[17];
  assign t[252] = t[304] ^ x[21];
  assign t[253] = t[305] ^ x[20];
  assign t[254] = t[306] ^ x[24];
  assign t[255] = t[307] ^ x[23];
  assign t[256] = t[308] ^ x[27];
  assign t[257] = t[309] ^ x[26];
  assign t[258] = t[310] ^ x[30];
  assign t[259] = t[311] ^ x[29];
  assign t[25] = t[44] ? t[45] : t[165];
  assign t[260] = t[312] ^ x[33];
  assign t[261] = t[313] ^ x[32];
  assign t[262] = t[314] ^ x[36];
  assign t[263] = t[315] ^ x[35];
  assign t[264] = t[316] ^ x[39];
  assign t[265] = t[317] ^ x[38];
  assign t[266] = t[318] ^ x[44];
  assign t[267] = t[319] ^ x[43];
  assign t[268] = t[320] ^ x[47];
  assign t[269] = t[321] ^ x[46];
  assign t[26] = t[46] ^ t[47];
  assign t[270] = t[322] ^ x[50];
  assign t[271] = t[323] ^ x[49];
  assign t[272] = t[324] ^ x[53];
  assign t[273] = t[325] ^ x[52];
  assign t[274] = t[326] ^ x[56];
  assign t[275] = t[327] ^ x[55];
  assign t[276] = t[328] ^ x[59];
  assign t[277] = t[329] ^ x[58];
  assign t[278] = t[330] ^ x[62];
  assign t[279] = t[331] ^ x[61];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[332] ^ x[69];
  assign t[281] = t[333] ^ x[68];
  assign t[282] = t[334] ^ x[74];
  assign t[283] = t[335] ^ x[73];
  assign t[284] = t[336] ^ x[77];
  assign t[285] = t[337] ^ x[76];
  assign t[286] = t[338] ^ x[82];
  assign t[287] = t[339] ^ x[81];
  assign t[288] = t[340] ^ x[93];
  assign t[289] = t[341] ^ x[92];
  assign t[28] = ~(t[50]);
  assign t[290] = t[342] ^ x[98];
  assign t[291] = t[343] ^ x[97];
  assign t[292] = t[344] ^ x[101];
  assign t[293] = t[345] ^ x[100];
  assign t[294] = (x[2]);
  assign t[295] = (x[2]);
  assign t[296] = (x[7]);
  assign t[297] = (x[7]);
  assign t[298] = (x[10]);
  assign t[299] = (x[10]);
  assign t[29] = ~(t[166]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[13]);
  assign t[301] = (x[13]);
  assign t[302] = (x[16]);
  assign t[303] = (x[16]);
  assign t[304] = (x[19]);
  assign t[305] = (x[19]);
  assign t[306] = (x[22]);
  assign t[307] = (x[22]);
  assign t[308] = (x[25]);
  assign t[309] = (x[25]);
  assign t[30] = ~(t[167]);
  assign t[310] = (x[28]);
  assign t[311] = (x[28]);
  assign t[312] = (x[31]);
  assign t[313] = (x[31]);
  assign t[314] = (x[34]);
  assign t[315] = (x[34]);
  assign t[316] = (x[37]);
  assign t[317] = (x[37]);
  assign t[318] = (x[42]);
  assign t[319] = (x[42]);
  assign t[31] = ~(t[168]);
  assign t[320] = (x[45]);
  assign t[321] = (x[45]);
  assign t[322] = (x[48]);
  assign t[323] = (x[48]);
  assign t[324] = (x[51]);
  assign t[325] = (x[51]);
  assign t[326] = (x[54]);
  assign t[327] = (x[54]);
  assign t[328] = (x[57]);
  assign t[329] = (x[57]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[60]);
  assign t[331] = (x[60]);
  assign t[332] = (x[67]);
  assign t[333] = (x[67]);
  assign t[334] = (x[72]);
  assign t[335] = (x[72]);
  assign t[336] = (x[75]);
  assign t[337] = (x[75]);
  assign t[338] = (x[80]);
  assign t[339] = (x[80]);
  assign t[33] = ~t[53];
  assign t[340] = (x[91]);
  assign t[341] = (x[91]);
  assign t[342] = (x[96]);
  assign t[343] = (x[96]);
  assign t[344] = (x[99]);
  assign t[345] = (x[99]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] ^ t[33];
  assign t[36] = t[57] & t[58];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[44] ? t[66] : t[169];
  assign t[42] = ~(t[67]);
  assign t[43] = t[44] ? t[68] : t[170];
  assign t[44] = ~(t[15]);
  assign t[45] = t[165] ^ t[69];
  assign t[46] = t[70] ^ t[24];
  assign t[47] = t[71] & t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[171] | t[75];
  assign t[4] = t[8] ? t[9] : t[164];
  assign t[50] = ~(t[76]);
  assign t[51] = ~(t[172]);
  assign t[52] = ~(t[77] & t[173]);
  assign t[53] = t[44] ? t[78] : t[174];
  assign t[54] = t[79] ^ t[36];
  assign t[55] = t[80] & t[81];
  assign t[56] = t[82];
  assign t[57] = ~(t[83]);
  assign t[58] = t[84];
  assign t[59] = t[85] ^ t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[87] & t[88];
  assign t[61] = t[173] ^ t[89];
  assign t[62] = t[64] ^ t[90];
  assign t[63] = t[166] ^ t[4];
  assign t[64] = t[91] ^ t[92];
  assign t[65] = t[93] & t[94];
  assign t[66] = t[169] ^ t[95];
  assign t[67] = t[44] ? t[96] : t[175];
  assign t[68] = t[170] ^ t[97];
  assign t[69] = t[98] ? x[41] : x[40];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[99] & t[100];
  assign t[71] = ~(t[101] ^ t[46]);
  assign t[72] = t[102] ^ t[43];
  assign t[73] = ~(t[75] & t[103]);
  assign t[74] = ~(t[176] ^ t[104]);
  assign t[75] = ~(t[105] & t[106]);
  assign t[76] = ~(t[49]);
  assign t[77] = ~(t[177]);
  assign t[78] = t[174] ^ t[107];
  assign t[79] = t[108] & t[109];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[110] ^ t[54]);
  assign t[81] = t[111] ^ t[58];
  assign t[82] = t[44] ? t[112] : t[178];
  assign t[83] = ~t[113];
  assign t[84] = t[27] ? t[114] : t[179];
  assign t[85] = t[27] ? t[115] : t[180];
  assign t[86] = t[27] ? t[116] : t[181];
  assign t[87] = ~(t[59] ^ t[117]);
  assign t[88] = t[118] ^ t[119];
  assign t[89] = t[8] ? t[120] : t[182];
  assign t[8] = ~(t[15]);
  assign t[90] = t[121] & t[122];
  assign t[91] = t[123] & t[124];
  assign t[92] = t[125] & t[126];
  assign t[93] = ~(t[91] ^ t[127]);
  assign t[94] = t[128] ^ t[129];
  assign t[95] = t[98] ? x[64] : x[63];
  assign t[96] = t[175] ^ t[130];
  assign t[97] = t[98] ? x[66] : x[65];
  assign t[98] = ~(t[50]);
  assign t[99] = ~(t[131]);
  assign t[9] = t[164] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind36(x, y);
 input [111:0] x;
 output y;

 wire [334:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[53] ^ t[25];
  assign t[101] = ~(t[129] & t[130]);
  assign t[102] = t[131] ^ t[173];
  assign t[103] = ~(t[168]);
  assign t[104] = t[132] & t[131];
  assign t[105] = t[170] ^ t[133];
  assign t[106] = t[134] ? x[72] : x[71];
  assign t[107] = t[134] ? x[74] : x[73];
  assign t[108] = ~(t[135]);
  assign t[109] = ~(t[36]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[37]);
  assign t[111] = t[78] ? t[136] : t[174];
  assign t[112] = t[171] ^ t[137];
  assign t[113] = t[138] ? x[79] : x[78];
  assign t[114] = t[74] ? x[81] : x[80];
  assign t[115] = ~(t[121]);
  assign t[116] = ~(t[139]);
  assign t[117] = ~(t[59]);
  assign t[118] = t[27] ? t[140] : t[175];
  assign t[119] = t[40] ^ t[139];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[139] ^ t[60];
  assign t[121] = t[118] ^ t[59];
  assign t[122] = t[134] ? x[86] : x[85];
  assign t[123] = t[134] ? x[88] : x[87];
  assign t[124] = t[141] & t[142];
  assign t[125] = t[143] & t[95];
  assign t[126] = t[78] ? t[144] : t[176];
  assign t[127] = t[172] ^ t[145];
  assign t[128] = t[35] ^ t[53];
  assign t[129] = ~(t[132] | t[131]);
  assign t[12] = t[21] ^ t[22];
  assign t[130] = ~(t[146] | t[103]);
  assign t[131] = ~(t[177]);
  assign t[132] = ~(t[173]);
  assign t[133] = t[28] ? x[96] : x[95];
  assign t[134] = ~(t[49]);
  assign t[135] = t[58] ^ t[37];
  assign t[136] = t[174] ^ t[147];
  assign t[137] = t[134] ? x[98] : x[97];
  assign t[138] = ~(t[49]);
  assign t[139] = t[27] ? t[148] : t[178];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[175] ^ t[149];
  assign t[141] = ~(t[150]);
  assign t[142] = ~(t[63]);
  assign t[143] = ~(t[64]);
  assign t[144] = t[176] ^ t[151];
  assign t[145] = t[134] ? x[103] : x[102];
  assign t[146] = ~(t[160]);
  assign t[147] = t[134] ? x[105] : x[104];
  assign t[148] = t[178] ^ t[152];
  assign t[149] = t[74] ? x[107] : x[106];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[95] ^ t[64];
  assign t[151] = t[134] ? x[109] : x[108];
  assign t[152] = t[138] ? x[111] : x[110];
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = t[205] ^ x[4];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[9];
  assign t[181] = t[207] ^ x[12];
  assign t[182] = t[208] ^ x[15];
  assign t[183] = t[209] ^ x[18];
  assign t[184] = t[210] ^ x[21];
  assign t[185] = t[211] ^ x[24];
  assign t[186] = t[212] ^ x[27];
  assign t[187] = t[213] ^ x[30];
  assign t[188] = t[214] ^ x[33];
  assign t[189] = t[215] ^ x[36];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[39];
  assign t[191] = t[217] ^ x[42];
  assign t[192] = t[218] ^ x[45];
  assign t[193] = t[219] ^ x[48];
  assign t[194] = t[220] ^ x[51];
  assign t[195] = t[221] ^ x[54];
  assign t[196] = t[222] ^ x[59];
  assign t[197] = t[223] ^ x[62];
  assign t[198] = t[224] ^ x[65];
  assign t[199] = t[225] ^ x[70];
  assign t[19] = t[33] ^ t[25];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[77];
  assign t[201] = t[227] ^ x[84];
  assign t[202] = t[228] ^ x[91];
  assign t[203] = t[229] ^ x[94];
  assign t[204] = t[230] ^ x[101];
  assign t[205] = (t[231] & ~t[232]);
  assign t[206] = (t[233] & ~t[234]);
  assign t[207] = (t[235] & ~t[236]);
  assign t[208] = (t[237] & ~t[238]);
  assign t[209] = (t[239] & ~t[240]);
  assign t[20] = t[34] & t[35];
  assign t[210] = (t[241] & ~t[242]);
  assign t[211] = (t[243] & ~t[244]);
  assign t[212] = (t[245] & ~t[246]);
  assign t[213] = (t[247] & ~t[248]);
  assign t[214] = (t[249] & ~t[250]);
  assign t[215] = (t[251] & ~t[252]);
  assign t[216] = (t[253] & ~t[254]);
  assign t[217] = (t[255] & ~t[256]);
  assign t[218] = (t[257] & ~t[258]);
  assign t[219] = (t[259] & ~t[260]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = (t[261] & ~t[262]);
  assign t[221] = (t[263] & ~t[264]);
  assign t[222] = (t[265] & ~t[266]);
  assign t[223] = (t[267] & ~t[268]);
  assign t[224] = (t[269] & ~t[270]);
  assign t[225] = (t[271] & ~t[272]);
  assign t[226] = (t[273] & ~t[274]);
  assign t[227] = (t[275] & ~t[276]);
  assign t[228] = (t[277] & ~t[278]);
  assign t[229] = (t[279] & ~t[280]);
  assign t[22] = t[38] & t[39];
  assign t[230] = (t[281] & ~t[282]);
  assign t[231] = t[283] ^ x[4];
  assign t[232] = t[284] ^ x[3];
  assign t[233] = t[285] ^ x[9];
  assign t[234] = t[286] ^ x[8];
  assign t[235] = t[287] ^ x[12];
  assign t[236] = t[288] ^ x[11];
  assign t[237] = t[289] ^ x[15];
  assign t[238] = t[290] ^ x[14];
  assign t[239] = t[291] ^ x[18];
  assign t[23] = t[40] ^ t[41];
  assign t[240] = t[292] ^ x[17];
  assign t[241] = t[293] ^ x[21];
  assign t[242] = t[294] ^ x[20];
  assign t[243] = t[295] ^ x[24];
  assign t[244] = t[296] ^ x[23];
  assign t[245] = t[297] ^ x[27];
  assign t[246] = t[298] ^ x[26];
  assign t[247] = t[299] ^ x[30];
  assign t[248] = t[300] ^ x[29];
  assign t[249] = t[301] ^ x[33];
  assign t[24] = t[42] ^ t[43];
  assign t[250] = t[302] ^ x[32];
  assign t[251] = t[303] ^ x[36];
  assign t[252] = t[304] ^ x[35];
  assign t[253] = t[305] ^ x[39];
  assign t[254] = t[306] ^ x[38];
  assign t[255] = t[307] ^ x[42];
  assign t[256] = t[308] ^ x[41];
  assign t[257] = t[309] ^ x[45];
  assign t[258] = t[310] ^ x[44];
  assign t[259] = t[311] ^ x[48];
  assign t[25] = t[154] ^ t[44];
  assign t[260] = t[312] ^ x[47];
  assign t[261] = t[313] ^ x[51];
  assign t[262] = t[314] ^ x[50];
  assign t[263] = t[315] ^ x[54];
  assign t[264] = t[316] ^ x[53];
  assign t[265] = t[317] ^ x[59];
  assign t[266] = t[318] ^ x[58];
  assign t[267] = t[319] ^ x[62];
  assign t[268] = t[320] ^ x[61];
  assign t[269] = t[321] ^ x[65];
  assign t[26] = t[45] ^ t[46];
  assign t[270] = t[322] ^ x[64];
  assign t[271] = t[323] ^ x[70];
  assign t[272] = t[324] ^ x[69];
  assign t[273] = t[325] ^ x[77];
  assign t[274] = t[326] ^ x[76];
  assign t[275] = t[327] ^ x[84];
  assign t[276] = t[328] ^ x[83];
  assign t[277] = t[329] ^ x[91];
  assign t[278] = t[330] ^ x[90];
  assign t[279] = t[331] ^ x[94];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[332] ^ x[93];
  assign t[281] = t[333] ^ x[101];
  assign t[282] = t[334] ^ x[100];
  assign t[283] = (x[2]);
  assign t[284] = (x[2]);
  assign t[285] = (x[7]);
  assign t[286] = (x[7]);
  assign t[287] = (x[10]);
  assign t[288] = (x[10]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[49]);
  assign t[290] = (x[13]);
  assign t[291] = (x[16]);
  assign t[292] = (x[16]);
  assign t[293] = (x[19]);
  assign t[294] = (x[19]);
  assign t[295] = (x[22]);
  assign t[296] = (x[22]);
  assign t[297] = (x[25]);
  assign t[298] = (x[25]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[28]);
  assign t[301] = (x[31]);
  assign t[302] = (x[31]);
  assign t[303] = (x[34]);
  assign t[304] = (x[34]);
  assign t[305] = (x[37]);
  assign t[306] = (x[37]);
  assign t[307] = (x[40]);
  assign t[308] = (x[40]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[156]);
  assign t[310] = (x[43]);
  assign t[311] = (x[46]);
  assign t[312] = (x[46]);
  assign t[313] = (x[49]);
  assign t[314] = (x[49]);
  assign t[315] = (x[52]);
  assign t[316] = (x[52]);
  assign t[317] = (x[57]);
  assign t[318] = (x[57]);
  assign t[319] = (x[60]);
  assign t[31] = ~(t[157]);
  assign t[320] = (x[60]);
  assign t[321] = (x[63]);
  assign t[322] = (x[63]);
  assign t[323] = (x[68]);
  assign t[324] = (x[68]);
  assign t[325] = (x[75]);
  assign t[326] = (x[75]);
  assign t[327] = (x[82]);
  assign t[328] = (x[82]);
  assign t[329] = (x[89]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[89]);
  assign t[331] = (x[92]);
  assign t[332] = (x[92]);
  assign t[333] = (x[99]);
  assign t[334] = (x[99]);
  assign t[33] = t[8] ? t[52] : t[158];
  assign t[34] = ~(t[53]);
  assign t[35] = t[156] ^ t[4];
  assign t[36] = t[54];
  assign t[37] = ~t[55];
  assign t[38] = ~(t[21] ^ t[56]);
  assign t[39] = t[57] ^ t[58];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[59] ^ t[60];
  assign t[41] = t[61] ^ t[62];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[65] & t[66];
  assign t[44] = t[8] ? t[67] : t[159];
  assign t[45] = t[68] ^ t[20];
  assign t[46] = t[69] & t[70];
  assign t[47] = ~(t[71] & t[72]);
  assign t[48] = t[160] | t[73];
  assign t[49] = ~(t[74]);
  assign t[4] = t[8] ? t[9] : t[153];
  assign t[50] = ~(t[161]);
  assign t[51] = ~(t[75] & t[154]);
  assign t[52] = t[158] ^ t[76];
  assign t[53] = t[155] ^ t[77];
  assign t[54] = t[78] ? t[79] : t[162];
  assign t[55] = t[78] ? t[80] : t[163];
  assign t[56] = t[81] ^ t[82];
  assign t[57] = t[37] ^ t[83];
  assign t[58] = t[84];
  assign t[59] = t[27] ? t[85] : t[164];
  assign t[5] = ~(t[10]);
  assign t[60] = t[27] ? t[86] : t[165];
  assign t[61] = t[87] ^ t[88];
  assign t[62] = t[89] & t[90];
  assign t[63] = t[78] ? t[91] : t[166];
  assign t[64] = t[78] ? t[92] : t[167];
  assign t[65] = ~(t[42] ^ t[93]);
  assign t[66] = t[94] ^ t[95];
  assign t[67] = t[159] ^ t[96];
  assign t[68] = t[97] & t[98];
  assign t[69] = ~(t[99] ^ t[45]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[100] ^ t[35];
  assign t[71] = ~(t[73] & t[101]);
  assign t[72] = ~(t[168] ^ t[102]);
  assign t[73] = ~(t[103] & t[104]);
  assign t[74] = ~(t[48]);
  assign t[75] = ~(t[169]);
  assign t[76] = t[28] ? x[56] : x[55];
  assign t[77] = t[8] ? t[105] : t[170];
  assign t[78] = ~(t[15]);
  assign t[79] = t[162] ^ t[106];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[163] ^ t[107];
  assign t[81] = t[108] & t[109];
  assign t[82] = t[110] & t[58];
  assign t[83] = ~t[111];
  assign t[84] = t[27] ? t[112] : t[171];
  assign t[85] = t[164] ^ t[113];
  assign t[86] = t[165] ^ t[114];
  assign t[87] = t[115] & t[116];
  assign t[88] = t[117] & t[118];
  assign t[89] = ~(t[87] ^ t[119]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[120] ^ t[121];
  assign t[91] = t[166] ^ t[122];
  assign t[92] = t[167] ^ t[123];
  assign t[93] = t[124] ^ t[125];
  assign t[94] = t[64] ^ t[126];
  assign t[95] = t[78] ? t[127] : t[172];
  assign t[96] = t[28] ? x[67] : x[66];
  assign t[97] = ~(t[128]);
  assign t[98] = ~(t[33]);
  assign t[99] = t[33] ^ t[53];
  assign t[9] = t[153] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind37(x, y);
 input [111:0] x;
 output y;

 wire [334:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[53] ^ t[25];
  assign t[101] = ~(t[129] & t[130]);
  assign t[102] = t[131] ^ t[173];
  assign t[103] = ~(t[168]);
  assign t[104] = t[132] & t[131];
  assign t[105] = t[170] ^ t[133];
  assign t[106] = t[134] ? x[72] : x[71];
  assign t[107] = t[134] ? x[74] : x[73];
  assign t[108] = ~(t[135]);
  assign t[109] = ~(t[36]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[37]);
  assign t[111] = t[78] ? t[136] : t[174];
  assign t[112] = t[171] ^ t[137];
  assign t[113] = t[138] ? x[79] : x[78];
  assign t[114] = t[74] ? x[81] : x[80];
  assign t[115] = ~(t[121]);
  assign t[116] = ~(t[139]);
  assign t[117] = ~(t[59]);
  assign t[118] = t[27] ? t[140] : t[175];
  assign t[119] = t[40] ^ t[139];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[139] ^ t[60];
  assign t[121] = t[118] ^ t[59];
  assign t[122] = t[134] ? x[86] : x[85];
  assign t[123] = t[134] ? x[88] : x[87];
  assign t[124] = t[141] & t[142];
  assign t[125] = t[143] & t[95];
  assign t[126] = t[78] ? t[144] : t[176];
  assign t[127] = t[172] ^ t[145];
  assign t[128] = t[35] ^ t[53];
  assign t[129] = ~(t[132] | t[131]);
  assign t[12] = t[21] ^ t[22];
  assign t[130] = ~(t[146] | t[103]);
  assign t[131] = ~(t[177]);
  assign t[132] = ~(t[173]);
  assign t[133] = t[28] ? x[96] : x[95];
  assign t[134] = ~(t[49]);
  assign t[135] = t[58] ^ t[37];
  assign t[136] = t[174] ^ t[147];
  assign t[137] = t[134] ? x[98] : x[97];
  assign t[138] = ~(t[49]);
  assign t[139] = t[27] ? t[148] : t[178];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[175] ^ t[149];
  assign t[141] = ~(t[150]);
  assign t[142] = ~(t[63]);
  assign t[143] = ~(t[64]);
  assign t[144] = t[176] ^ t[151];
  assign t[145] = t[134] ? x[103] : x[102];
  assign t[146] = ~(t[160]);
  assign t[147] = t[134] ? x[105] : x[104];
  assign t[148] = t[178] ^ t[152];
  assign t[149] = t[74] ? x[107] : x[106];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[95] ^ t[64];
  assign t[151] = t[134] ? x[109] : x[108];
  assign t[152] = t[138] ? x[111] : x[110];
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = t[205] ^ x[4];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[9];
  assign t[181] = t[207] ^ x[12];
  assign t[182] = t[208] ^ x[15];
  assign t[183] = t[209] ^ x[18];
  assign t[184] = t[210] ^ x[21];
  assign t[185] = t[211] ^ x[24];
  assign t[186] = t[212] ^ x[27];
  assign t[187] = t[213] ^ x[30];
  assign t[188] = t[214] ^ x[33];
  assign t[189] = t[215] ^ x[36];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[39];
  assign t[191] = t[217] ^ x[42];
  assign t[192] = t[218] ^ x[45];
  assign t[193] = t[219] ^ x[48];
  assign t[194] = t[220] ^ x[51];
  assign t[195] = t[221] ^ x[54];
  assign t[196] = t[222] ^ x[59];
  assign t[197] = t[223] ^ x[62];
  assign t[198] = t[224] ^ x[65];
  assign t[199] = t[225] ^ x[70];
  assign t[19] = t[33] ^ t[25];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[77];
  assign t[201] = t[227] ^ x[84];
  assign t[202] = t[228] ^ x[91];
  assign t[203] = t[229] ^ x[94];
  assign t[204] = t[230] ^ x[101];
  assign t[205] = (t[231] & ~t[232]);
  assign t[206] = (t[233] & ~t[234]);
  assign t[207] = (t[235] & ~t[236]);
  assign t[208] = (t[237] & ~t[238]);
  assign t[209] = (t[239] & ~t[240]);
  assign t[20] = t[34] & t[35];
  assign t[210] = (t[241] & ~t[242]);
  assign t[211] = (t[243] & ~t[244]);
  assign t[212] = (t[245] & ~t[246]);
  assign t[213] = (t[247] & ~t[248]);
  assign t[214] = (t[249] & ~t[250]);
  assign t[215] = (t[251] & ~t[252]);
  assign t[216] = (t[253] & ~t[254]);
  assign t[217] = (t[255] & ~t[256]);
  assign t[218] = (t[257] & ~t[258]);
  assign t[219] = (t[259] & ~t[260]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = (t[261] & ~t[262]);
  assign t[221] = (t[263] & ~t[264]);
  assign t[222] = (t[265] & ~t[266]);
  assign t[223] = (t[267] & ~t[268]);
  assign t[224] = (t[269] & ~t[270]);
  assign t[225] = (t[271] & ~t[272]);
  assign t[226] = (t[273] & ~t[274]);
  assign t[227] = (t[275] & ~t[276]);
  assign t[228] = (t[277] & ~t[278]);
  assign t[229] = (t[279] & ~t[280]);
  assign t[22] = t[38] & t[39];
  assign t[230] = (t[281] & ~t[282]);
  assign t[231] = t[283] ^ x[4];
  assign t[232] = t[284] ^ x[3];
  assign t[233] = t[285] ^ x[9];
  assign t[234] = t[286] ^ x[8];
  assign t[235] = t[287] ^ x[12];
  assign t[236] = t[288] ^ x[11];
  assign t[237] = t[289] ^ x[15];
  assign t[238] = t[290] ^ x[14];
  assign t[239] = t[291] ^ x[18];
  assign t[23] = t[40] ^ t[41];
  assign t[240] = t[292] ^ x[17];
  assign t[241] = t[293] ^ x[21];
  assign t[242] = t[294] ^ x[20];
  assign t[243] = t[295] ^ x[24];
  assign t[244] = t[296] ^ x[23];
  assign t[245] = t[297] ^ x[27];
  assign t[246] = t[298] ^ x[26];
  assign t[247] = t[299] ^ x[30];
  assign t[248] = t[300] ^ x[29];
  assign t[249] = t[301] ^ x[33];
  assign t[24] = t[42] ^ t[43];
  assign t[250] = t[302] ^ x[32];
  assign t[251] = t[303] ^ x[36];
  assign t[252] = t[304] ^ x[35];
  assign t[253] = t[305] ^ x[39];
  assign t[254] = t[306] ^ x[38];
  assign t[255] = t[307] ^ x[42];
  assign t[256] = t[308] ^ x[41];
  assign t[257] = t[309] ^ x[45];
  assign t[258] = t[310] ^ x[44];
  assign t[259] = t[311] ^ x[48];
  assign t[25] = t[154] ^ t[44];
  assign t[260] = t[312] ^ x[47];
  assign t[261] = t[313] ^ x[51];
  assign t[262] = t[314] ^ x[50];
  assign t[263] = t[315] ^ x[54];
  assign t[264] = t[316] ^ x[53];
  assign t[265] = t[317] ^ x[59];
  assign t[266] = t[318] ^ x[58];
  assign t[267] = t[319] ^ x[62];
  assign t[268] = t[320] ^ x[61];
  assign t[269] = t[321] ^ x[65];
  assign t[26] = t[45] ^ t[46];
  assign t[270] = t[322] ^ x[64];
  assign t[271] = t[323] ^ x[70];
  assign t[272] = t[324] ^ x[69];
  assign t[273] = t[325] ^ x[77];
  assign t[274] = t[326] ^ x[76];
  assign t[275] = t[327] ^ x[84];
  assign t[276] = t[328] ^ x[83];
  assign t[277] = t[329] ^ x[91];
  assign t[278] = t[330] ^ x[90];
  assign t[279] = t[331] ^ x[94];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[332] ^ x[93];
  assign t[281] = t[333] ^ x[101];
  assign t[282] = t[334] ^ x[100];
  assign t[283] = (x[2]);
  assign t[284] = (x[2]);
  assign t[285] = (x[7]);
  assign t[286] = (x[7]);
  assign t[287] = (x[10]);
  assign t[288] = (x[10]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[49]);
  assign t[290] = (x[13]);
  assign t[291] = (x[16]);
  assign t[292] = (x[16]);
  assign t[293] = (x[19]);
  assign t[294] = (x[19]);
  assign t[295] = (x[22]);
  assign t[296] = (x[22]);
  assign t[297] = (x[25]);
  assign t[298] = (x[25]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[28]);
  assign t[301] = (x[31]);
  assign t[302] = (x[31]);
  assign t[303] = (x[34]);
  assign t[304] = (x[34]);
  assign t[305] = (x[37]);
  assign t[306] = (x[37]);
  assign t[307] = (x[40]);
  assign t[308] = (x[40]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[156]);
  assign t[310] = (x[43]);
  assign t[311] = (x[46]);
  assign t[312] = (x[46]);
  assign t[313] = (x[49]);
  assign t[314] = (x[49]);
  assign t[315] = (x[52]);
  assign t[316] = (x[52]);
  assign t[317] = (x[57]);
  assign t[318] = (x[57]);
  assign t[319] = (x[60]);
  assign t[31] = ~(t[157]);
  assign t[320] = (x[60]);
  assign t[321] = (x[63]);
  assign t[322] = (x[63]);
  assign t[323] = (x[68]);
  assign t[324] = (x[68]);
  assign t[325] = (x[75]);
  assign t[326] = (x[75]);
  assign t[327] = (x[82]);
  assign t[328] = (x[82]);
  assign t[329] = (x[89]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[89]);
  assign t[331] = (x[92]);
  assign t[332] = (x[92]);
  assign t[333] = (x[99]);
  assign t[334] = (x[99]);
  assign t[33] = t[8] ? t[52] : t[158];
  assign t[34] = ~(t[53]);
  assign t[35] = t[156] ^ t[4];
  assign t[36] = t[54];
  assign t[37] = ~t[55];
  assign t[38] = ~(t[21] ^ t[56]);
  assign t[39] = t[57] ^ t[58];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[59] ^ t[60];
  assign t[41] = t[61] ^ t[62];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[65] & t[66];
  assign t[44] = t[8] ? t[67] : t[159];
  assign t[45] = t[68] ^ t[20];
  assign t[46] = t[69] & t[70];
  assign t[47] = ~(t[71] & t[72]);
  assign t[48] = t[160] | t[73];
  assign t[49] = ~(t[74]);
  assign t[4] = t[8] ? t[9] : t[153];
  assign t[50] = ~(t[161]);
  assign t[51] = ~(t[75] & t[154]);
  assign t[52] = t[158] ^ t[76];
  assign t[53] = t[155] ^ t[77];
  assign t[54] = t[78] ? t[79] : t[162];
  assign t[55] = t[78] ? t[80] : t[163];
  assign t[56] = t[81] ^ t[82];
  assign t[57] = t[37] ^ t[83];
  assign t[58] = t[84];
  assign t[59] = t[27] ? t[85] : t[164];
  assign t[5] = ~(t[10]);
  assign t[60] = t[27] ? t[86] : t[165];
  assign t[61] = t[87] ^ t[88];
  assign t[62] = t[89] & t[90];
  assign t[63] = t[78] ? t[91] : t[166];
  assign t[64] = t[78] ? t[92] : t[167];
  assign t[65] = ~(t[42] ^ t[93]);
  assign t[66] = t[94] ^ t[95];
  assign t[67] = t[159] ^ t[96];
  assign t[68] = t[97] & t[98];
  assign t[69] = ~(t[99] ^ t[45]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[100] ^ t[35];
  assign t[71] = ~(t[73] & t[101]);
  assign t[72] = ~(t[168] ^ t[102]);
  assign t[73] = ~(t[103] & t[104]);
  assign t[74] = ~(t[48]);
  assign t[75] = ~(t[169]);
  assign t[76] = t[28] ? x[56] : x[55];
  assign t[77] = t[8] ? t[105] : t[170];
  assign t[78] = ~(t[15]);
  assign t[79] = t[162] ^ t[106];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[163] ^ t[107];
  assign t[81] = t[108] & t[109];
  assign t[82] = t[110] & t[58];
  assign t[83] = ~t[111];
  assign t[84] = t[27] ? t[112] : t[171];
  assign t[85] = t[164] ^ t[113];
  assign t[86] = t[165] ^ t[114];
  assign t[87] = t[115] & t[116];
  assign t[88] = t[117] & t[118];
  assign t[89] = ~(t[87] ^ t[119]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[120] ^ t[121];
  assign t[91] = t[166] ^ t[122];
  assign t[92] = t[167] ^ t[123];
  assign t[93] = t[124] ^ t[125];
  assign t[94] = t[64] ^ t[126];
  assign t[95] = t[78] ? t[127] : t[172];
  assign t[96] = t[28] ? x[67] : x[66];
  assign t[97] = ~(t[128]);
  assign t[98] = ~(t[33]);
  assign t[99] = t[33] ^ t[53];
  assign t[9] = t[153] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind38(x, y);
 input [111:0] x;
 output y;

 wire [333:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[128] & t[127];
  assign t[101] = t[122] ? x[65] : x[64];
  assign t[102] = t[122] ? x[67] : x[66];
  assign t[103] = ~(t[109]);
  assign t[104] = ~(t[129]);
  assign t[105] = ~(t[51]);
  assign t[106] = t[62] ? t[130] : t[170];
  assign t[107] = t[33] ^ t[129];
  assign t[108] = t[129] ^ t[52];
  assign t[109] = t[106] ^ t[51];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[131]);
  assign t[111] = ~(t[132]);
  assign t[112] = ~(t[133]);
  assign t[113] = t[27] ? t[134] : t[171];
  assign t[114] = t[132] ^ t[133];
  assign t[115] = t[133] ^ t[35];
  assign t[116] = t[28] ? x[75] : x[74];
  assign t[117] = ~(t[135]);
  assign t[118] = ~(t[4]);
  assign t[119] = ~(t[37]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[8] ? t[136] : t[172];
  assign t[121] = t[167] ^ t[137];
  assign t[122] = ~(t[48]);
  assign t[123] = t[62] ? t[138] : t[173];
  assign t[124] = t[168] ^ t[139];
  assign t[125] = ~(t[128] | t[127]);
  assign t[126] = ~(t[140] | t[99]);
  assign t[127] = ~(t[174]);
  assign t[128] = ~(t[169]);
  assign t[129] = t[62] ? t[141] : t[175];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[170] ^ t[142];
  assign t[131] = t[113] ^ t[133];
  assign t[132] = t[27] ? t[143] : t[176];
  assign t[133] = t[27] ? t[144] : t[177];
  assign t[134] = t[171] ^ t[145];
  assign t[135] = t[61] ^ t[37];
  assign t[136] = t[172] ^ t[146];
  assign t[137] = t[28] ? x[95] : x[94];
  assign t[138] = t[173] ^ t[147];
  assign t[139] = t[122] ? x[97] : x[96];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[159]);
  assign t[141] = t[175] ^ t[148];
  assign t[142] = t[122] ? x[99] : x[98];
  assign t[143] = t[176] ^ t[149];
  assign t[144] = t[177] ^ t[150];
  assign t[145] = t[75] ? x[101] : x[100];
  assign t[146] = t[28] ? x[103] : x[102];
  assign t[147] = t[122] ? x[105] : x[104];
  assign t[148] = t[122] ? x[107] : x[106];
  assign t[149] = t[151] ? x[109] : x[108];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[151] ? x[111] : x[110];
  assign t[151] = ~(t[48]);
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = t[204] ^ x[4];
  assign t[179] = t[205] ^ x[9];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[12];
  assign t[181] = t[207] ^ x[15];
  assign t[182] = t[208] ^ x[18];
  assign t[183] = t[209] ^ x[21];
  assign t[184] = t[210] ^ x[24];
  assign t[185] = t[211] ^ x[27];
  assign t[186] = t[212] ^ x[30];
  assign t[187] = t[213] ^ x[33];
  assign t[188] = t[214] ^ x[36];
  assign t[189] = t[215] ^ x[39];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[42];
  assign t[191] = t[217] ^ x[45];
  assign t[192] = t[218] ^ x[48];
  assign t[193] = t[219] ^ x[53];
  assign t[194] = t[220] ^ x[60];
  assign t[195] = t[221] ^ x[63];
  assign t[196] = t[222] ^ x[70];
  assign t[197] = t[223] ^ x[73];
  assign t[198] = t[224] ^ x[78];
  assign t[199] = t[225] ^ x[81];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[84];
  assign t[201] = t[227] ^ x[87];
  assign t[202] = t[228] ^ x[90];
  assign t[203] = t[229] ^ x[93];
  assign t[204] = (t[230] & ~t[231]);
  assign t[205] = (t[232] & ~t[233]);
  assign t[206] = (t[234] & ~t[235]);
  assign t[207] = (t[236] & ~t[237]);
  assign t[208] = (t[238] & ~t[239]);
  assign t[209] = (t[240] & ~t[241]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[242] & ~t[243]);
  assign t[211] = (t[244] & ~t[245]);
  assign t[212] = (t[246] & ~t[247]);
  assign t[213] = (t[248] & ~t[249]);
  assign t[214] = (t[250] & ~t[251]);
  assign t[215] = (t[252] & ~t[253]);
  assign t[216] = (t[254] & ~t[255]);
  assign t[217] = (t[256] & ~t[257]);
  assign t[218] = (t[258] & ~t[259]);
  assign t[219] = (t[260] & ~t[261]);
  assign t[21] = t[4] ^ t[37];
  assign t[220] = (t[262] & ~t[263]);
  assign t[221] = (t[264] & ~t[265]);
  assign t[222] = (t[266] & ~t[267]);
  assign t[223] = (t[268] & ~t[269]);
  assign t[224] = (t[270] & ~t[271]);
  assign t[225] = (t[272] & ~t[273]);
  assign t[226] = (t[274] & ~t[275]);
  assign t[227] = (t[276] & ~t[277]);
  assign t[228] = (t[278] & ~t[279]);
  assign t[229] = (t[280] & ~t[281]);
  assign t[22] = t[38] & t[39];
  assign t[230] = t[282] ^ x[4];
  assign t[231] = t[283] ^ x[3];
  assign t[232] = t[284] ^ x[9];
  assign t[233] = t[285] ^ x[8];
  assign t[234] = t[286] ^ x[12];
  assign t[235] = t[287] ^ x[11];
  assign t[236] = t[288] ^ x[15];
  assign t[237] = t[289] ^ x[14];
  assign t[238] = t[290] ^ x[18];
  assign t[239] = t[291] ^ x[17];
  assign t[23] = ~t[40];
  assign t[240] = t[292] ^ x[21];
  assign t[241] = t[293] ^ x[20];
  assign t[242] = t[294] ^ x[24];
  assign t[243] = t[295] ^ x[23];
  assign t[244] = t[296] ^ x[27];
  assign t[245] = t[297] ^ x[26];
  assign t[246] = t[298] ^ x[30];
  assign t[247] = t[299] ^ x[29];
  assign t[248] = t[300] ^ x[33];
  assign t[249] = t[301] ^ x[32];
  assign t[24] = ~t[41];
  assign t[250] = t[302] ^ x[36];
  assign t[251] = t[303] ^ x[35];
  assign t[252] = t[304] ^ x[39];
  assign t[253] = t[305] ^ x[38];
  assign t[254] = t[306] ^ x[42];
  assign t[255] = t[307] ^ x[41];
  assign t[256] = t[308] ^ x[45];
  assign t[257] = t[309] ^ x[44];
  assign t[258] = t[310] ^ x[48];
  assign t[259] = t[311] ^ x[47];
  assign t[25] = t[42] ^ t[43];
  assign t[260] = t[312] ^ x[53];
  assign t[261] = t[313] ^ x[52];
  assign t[262] = t[314] ^ x[60];
  assign t[263] = t[315] ^ x[59];
  assign t[264] = t[316] ^ x[63];
  assign t[265] = t[317] ^ x[62];
  assign t[266] = t[318] ^ x[70];
  assign t[267] = t[319] ^ x[69];
  assign t[268] = t[320] ^ x[73];
  assign t[269] = t[321] ^ x[72];
  assign t[26] = t[44] & t[45];
  assign t[270] = t[322] ^ x[78];
  assign t[271] = t[323] ^ x[77];
  assign t[272] = t[324] ^ x[81];
  assign t[273] = t[325] ^ x[80];
  assign t[274] = t[326] ^ x[84];
  assign t[275] = t[327] ^ x[83];
  assign t[276] = t[328] ^ x[87];
  assign t[277] = t[329] ^ x[86];
  assign t[278] = t[330] ^ x[90];
  assign t[279] = t[331] ^ x[89];
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = t[332] ^ x[93];
  assign t[281] = t[333] ^ x[92];
  assign t[282] = (x[2]);
  assign t[283] = (x[2]);
  assign t[284] = (x[7]);
  assign t[285] = (x[7]);
  assign t[286] = (x[10]);
  assign t[287] = (x[10]);
  assign t[288] = (x[13]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[48]);
  assign t[290] = (x[16]);
  assign t[291] = (x[16]);
  assign t[292] = (x[19]);
  assign t[293] = (x[19]);
  assign t[294] = (x[22]);
  assign t[295] = (x[22]);
  assign t[296] = (x[25]);
  assign t[297] = (x[25]);
  assign t[298] = (x[28]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[153]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[31]);
  assign t[301] = (x[31]);
  assign t[302] = (x[34]);
  assign t[303] = (x[34]);
  assign t[304] = (x[37]);
  assign t[305] = (x[37]);
  assign t[306] = (x[40]);
  assign t[307] = (x[40]);
  assign t[308] = (x[43]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[154]);
  assign t[310] = (x[46]);
  assign t[311] = (x[46]);
  assign t[312] = (x[51]);
  assign t[313] = (x[51]);
  assign t[314] = (x[58]);
  assign t[315] = (x[58]);
  assign t[316] = (x[61]);
  assign t[317] = (x[61]);
  assign t[318] = (x[68]);
  assign t[319] = (x[68]);
  assign t[31] = ~(t[155]);
  assign t[320] = (x[71]);
  assign t[321] = (x[71]);
  assign t[322] = (x[76]);
  assign t[323] = (x[76]);
  assign t[324] = (x[79]);
  assign t[325] = (x[79]);
  assign t[326] = (x[82]);
  assign t[327] = (x[82]);
  assign t[328] = (x[85]);
  assign t[329] = (x[85]);
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = (x[88]);
  assign t[331] = (x[88]);
  assign t[332] = (x[91]);
  assign t[333] = (x[91]);
  assign t[33] = t[51] ^ t[52];
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[27] ? t[55] : t[156];
  assign t[36] = t[56] ^ t[57];
  assign t[37] = t[153] ^ t[58];
  assign t[38] = ~(t[21] ^ t[59]);
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[62] ? t[63] : t[157];
  assign t[41] = t[62] ? t[64] : t[158];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[67] & t[68];
  assign t[44] = ~(t[42] ^ t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[159] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[160]);
  assign t[4] = t[8] ? t[9] : t[152];
  assign t[50] = ~(t[76] & t[161]);
  assign t[51] = t[62] ? t[77] : t[162];
  assign t[52] = t[62] ? t[78] : t[163];
  assign t[53] = t[79] ^ t[80];
  assign t[54] = t[81] & t[82];
  assign t[55] = t[156] ^ t[83];
  assign t[56] = t[84] ^ t[85];
  assign t[57] = t[86] & t[87];
  assign t[58] = t[8] ? t[88] : t[164];
  assign t[59] = t[89] ^ t[90];
  assign t[5] = ~(t[10]);
  assign t[60] = t[37] ^ t[91];
  assign t[61] = t[154] ^ t[92];
  assign t[62] = ~(t[15]);
  assign t[63] = t[157] ^ t[93];
  assign t[64] = t[158] ^ t[94];
  assign t[65] = ~(t[71]);
  assign t[66] = ~(t[95]);
  assign t[67] = ~(t[23]);
  assign t[68] = t[96];
  assign t[69] = t[13] ^ t[95];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[95] ^ t[24];
  assign t[71] = t[68] ^ t[23];
  assign t[72] = ~(t[74] & t[97]);
  assign t[73] = ~(t[165] ^ t[98]);
  assign t[74] = ~(t[99] & t[100]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[166]);
  assign t[77] = t[162] ^ t[101];
  assign t[78] = t[163] ^ t[102];
  assign t[79] = t[103] & t[104];
  assign t[7] = t[13] ^ t[14];
  assign t[80] = t[105] & t[106];
  assign t[81] = ~(t[79] ^ t[107]);
  assign t[82] = t[108] ^ t[109];
  assign t[83] = t[75] ? x[50] : x[49];
  assign t[84] = t[110] & t[111];
  assign t[85] = t[112] & t[113];
  assign t[86] = ~(t[114] ^ t[56]);
  assign t[87] = t[115] ^ t[113];
  assign t[88] = t[164] ^ t[116];
  assign t[89] = t[117] & t[118];
  assign t[8] = ~(t[15]);
  assign t[90] = t[119] & t[61];
  assign t[91] = t[161] ^ t[120];
  assign t[92] = t[8] ? t[121] : t[167];
  assign t[93] = t[122] ? x[55] : x[54];
  assign t[94] = t[122] ? x[57] : x[56];
  assign t[95] = t[123];
  assign t[96] = t[27] ? t[124] : t[168];
  assign t[97] = ~(t[125] & t[126]);
  assign t[98] = t[127] ^ t[169];
  assign t[99] = ~(t[165]);
  assign t[9] = t[152] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind39(x, y);
 input [111:0] x;
 output y;

 wire [333:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[128] & t[127];
  assign t[101] = t[122] ? x[65] : x[64];
  assign t[102] = t[122] ? x[67] : x[66];
  assign t[103] = ~(t[109]);
  assign t[104] = ~(t[129]);
  assign t[105] = ~(t[51]);
  assign t[106] = t[62] ? t[130] : t[170];
  assign t[107] = t[33] ^ t[129];
  assign t[108] = t[129] ^ t[52];
  assign t[109] = t[106] ^ t[51];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[131]);
  assign t[111] = ~(t[132]);
  assign t[112] = ~(t[133]);
  assign t[113] = t[27] ? t[134] : t[171];
  assign t[114] = t[132] ^ t[133];
  assign t[115] = t[133] ^ t[35];
  assign t[116] = t[28] ? x[75] : x[74];
  assign t[117] = ~(t[135]);
  assign t[118] = ~(t[4]);
  assign t[119] = ~(t[37]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[8] ? t[136] : t[172];
  assign t[121] = t[167] ^ t[137];
  assign t[122] = ~(t[48]);
  assign t[123] = t[62] ? t[138] : t[173];
  assign t[124] = t[168] ^ t[139];
  assign t[125] = ~(t[128] | t[127]);
  assign t[126] = ~(t[140] | t[99]);
  assign t[127] = ~(t[174]);
  assign t[128] = ~(t[169]);
  assign t[129] = t[62] ? t[141] : t[175];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[170] ^ t[142];
  assign t[131] = t[113] ^ t[133];
  assign t[132] = t[27] ? t[143] : t[176];
  assign t[133] = t[27] ? t[144] : t[177];
  assign t[134] = t[171] ^ t[145];
  assign t[135] = t[61] ^ t[37];
  assign t[136] = t[172] ^ t[146];
  assign t[137] = t[28] ? x[95] : x[94];
  assign t[138] = t[173] ^ t[147];
  assign t[139] = t[122] ? x[97] : x[96];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[159]);
  assign t[141] = t[175] ^ t[148];
  assign t[142] = t[122] ? x[99] : x[98];
  assign t[143] = t[176] ^ t[149];
  assign t[144] = t[177] ^ t[150];
  assign t[145] = t[75] ? x[101] : x[100];
  assign t[146] = t[28] ? x[103] : x[102];
  assign t[147] = t[122] ? x[105] : x[104];
  assign t[148] = t[122] ? x[107] : x[106];
  assign t[149] = t[151] ? x[109] : x[108];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[151] ? x[111] : x[110];
  assign t[151] = ~(t[48]);
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = t[204] ^ x[4];
  assign t[179] = t[205] ^ x[9];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[12];
  assign t[181] = t[207] ^ x[15];
  assign t[182] = t[208] ^ x[18];
  assign t[183] = t[209] ^ x[21];
  assign t[184] = t[210] ^ x[24];
  assign t[185] = t[211] ^ x[27];
  assign t[186] = t[212] ^ x[30];
  assign t[187] = t[213] ^ x[33];
  assign t[188] = t[214] ^ x[36];
  assign t[189] = t[215] ^ x[39];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[42];
  assign t[191] = t[217] ^ x[45];
  assign t[192] = t[218] ^ x[48];
  assign t[193] = t[219] ^ x[53];
  assign t[194] = t[220] ^ x[60];
  assign t[195] = t[221] ^ x[63];
  assign t[196] = t[222] ^ x[70];
  assign t[197] = t[223] ^ x[73];
  assign t[198] = t[224] ^ x[78];
  assign t[199] = t[225] ^ x[81];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[84];
  assign t[201] = t[227] ^ x[87];
  assign t[202] = t[228] ^ x[90];
  assign t[203] = t[229] ^ x[93];
  assign t[204] = (t[230] & ~t[231]);
  assign t[205] = (t[232] & ~t[233]);
  assign t[206] = (t[234] & ~t[235]);
  assign t[207] = (t[236] & ~t[237]);
  assign t[208] = (t[238] & ~t[239]);
  assign t[209] = (t[240] & ~t[241]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[242] & ~t[243]);
  assign t[211] = (t[244] & ~t[245]);
  assign t[212] = (t[246] & ~t[247]);
  assign t[213] = (t[248] & ~t[249]);
  assign t[214] = (t[250] & ~t[251]);
  assign t[215] = (t[252] & ~t[253]);
  assign t[216] = (t[254] & ~t[255]);
  assign t[217] = (t[256] & ~t[257]);
  assign t[218] = (t[258] & ~t[259]);
  assign t[219] = (t[260] & ~t[261]);
  assign t[21] = t[4] ^ t[37];
  assign t[220] = (t[262] & ~t[263]);
  assign t[221] = (t[264] & ~t[265]);
  assign t[222] = (t[266] & ~t[267]);
  assign t[223] = (t[268] & ~t[269]);
  assign t[224] = (t[270] & ~t[271]);
  assign t[225] = (t[272] & ~t[273]);
  assign t[226] = (t[274] & ~t[275]);
  assign t[227] = (t[276] & ~t[277]);
  assign t[228] = (t[278] & ~t[279]);
  assign t[229] = (t[280] & ~t[281]);
  assign t[22] = t[38] & t[39];
  assign t[230] = t[282] ^ x[4];
  assign t[231] = t[283] ^ x[3];
  assign t[232] = t[284] ^ x[9];
  assign t[233] = t[285] ^ x[8];
  assign t[234] = t[286] ^ x[12];
  assign t[235] = t[287] ^ x[11];
  assign t[236] = t[288] ^ x[15];
  assign t[237] = t[289] ^ x[14];
  assign t[238] = t[290] ^ x[18];
  assign t[239] = t[291] ^ x[17];
  assign t[23] = ~t[40];
  assign t[240] = t[292] ^ x[21];
  assign t[241] = t[293] ^ x[20];
  assign t[242] = t[294] ^ x[24];
  assign t[243] = t[295] ^ x[23];
  assign t[244] = t[296] ^ x[27];
  assign t[245] = t[297] ^ x[26];
  assign t[246] = t[298] ^ x[30];
  assign t[247] = t[299] ^ x[29];
  assign t[248] = t[300] ^ x[33];
  assign t[249] = t[301] ^ x[32];
  assign t[24] = ~t[41];
  assign t[250] = t[302] ^ x[36];
  assign t[251] = t[303] ^ x[35];
  assign t[252] = t[304] ^ x[39];
  assign t[253] = t[305] ^ x[38];
  assign t[254] = t[306] ^ x[42];
  assign t[255] = t[307] ^ x[41];
  assign t[256] = t[308] ^ x[45];
  assign t[257] = t[309] ^ x[44];
  assign t[258] = t[310] ^ x[48];
  assign t[259] = t[311] ^ x[47];
  assign t[25] = t[42] ^ t[43];
  assign t[260] = t[312] ^ x[53];
  assign t[261] = t[313] ^ x[52];
  assign t[262] = t[314] ^ x[60];
  assign t[263] = t[315] ^ x[59];
  assign t[264] = t[316] ^ x[63];
  assign t[265] = t[317] ^ x[62];
  assign t[266] = t[318] ^ x[70];
  assign t[267] = t[319] ^ x[69];
  assign t[268] = t[320] ^ x[73];
  assign t[269] = t[321] ^ x[72];
  assign t[26] = t[44] & t[45];
  assign t[270] = t[322] ^ x[78];
  assign t[271] = t[323] ^ x[77];
  assign t[272] = t[324] ^ x[81];
  assign t[273] = t[325] ^ x[80];
  assign t[274] = t[326] ^ x[84];
  assign t[275] = t[327] ^ x[83];
  assign t[276] = t[328] ^ x[87];
  assign t[277] = t[329] ^ x[86];
  assign t[278] = t[330] ^ x[90];
  assign t[279] = t[331] ^ x[89];
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = t[332] ^ x[93];
  assign t[281] = t[333] ^ x[92];
  assign t[282] = (x[2]);
  assign t[283] = (x[2]);
  assign t[284] = (x[7]);
  assign t[285] = (x[7]);
  assign t[286] = (x[10]);
  assign t[287] = (x[10]);
  assign t[288] = (x[13]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[48]);
  assign t[290] = (x[16]);
  assign t[291] = (x[16]);
  assign t[292] = (x[19]);
  assign t[293] = (x[19]);
  assign t[294] = (x[22]);
  assign t[295] = (x[22]);
  assign t[296] = (x[25]);
  assign t[297] = (x[25]);
  assign t[298] = (x[28]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[153]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[31]);
  assign t[301] = (x[31]);
  assign t[302] = (x[34]);
  assign t[303] = (x[34]);
  assign t[304] = (x[37]);
  assign t[305] = (x[37]);
  assign t[306] = (x[40]);
  assign t[307] = (x[40]);
  assign t[308] = (x[43]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[154]);
  assign t[310] = (x[46]);
  assign t[311] = (x[46]);
  assign t[312] = (x[51]);
  assign t[313] = (x[51]);
  assign t[314] = (x[58]);
  assign t[315] = (x[58]);
  assign t[316] = (x[61]);
  assign t[317] = (x[61]);
  assign t[318] = (x[68]);
  assign t[319] = (x[68]);
  assign t[31] = ~(t[155]);
  assign t[320] = (x[71]);
  assign t[321] = (x[71]);
  assign t[322] = (x[76]);
  assign t[323] = (x[76]);
  assign t[324] = (x[79]);
  assign t[325] = (x[79]);
  assign t[326] = (x[82]);
  assign t[327] = (x[82]);
  assign t[328] = (x[85]);
  assign t[329] = (x[85]);
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = (x[88]);
  assign t[331] = (x[88]);
  assign t[332] = (x[91]);
  assign t[333] = (x[91]);
  assign t[33] = t[51] ^ t[52];
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[27] ? t[55] : t[156];
  assign t[36] = t[56] ^ t[57];
  assign t[37] = t[153] ^ t[58];
  assign t[38] = ~(t[21] ^ t[59]);
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[62] ? t[63] : t[157];
  assign t[41] = t[62] ? t[64] : t[158];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[67] & t[68];
  assign t[44] = ~(t[42] ^ t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[159] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[160]);
  assign t[4] = t[8] ? t[9] : t[152];
  assign t[50] = ~(t[76] & t[161]);
  assign t[51] = t[62] ? t[77] : t[162];
  assign t[52] = t[62] ? t[78] : t[163];
  assign t[53] = t[79] ^ t[80];
  assign t[54] = t[81] & t[82];
  assign t[55] = t[156] ^ t[83];
  assign t[56] = t[84] ^ t[85];
  assign t[57] = t[86] & t[87];
  assign t[58] = t[8] ? t[88] : t[164];
  assign t[59] = t[89] ^ t[90];
  assign t[5] = ~(t[10]);
  assign t[60] = t[37] ^ t[91];
  assign t[61] = t[154] ^ t[92];
  assign t[62] = ~(t[15]);
  assign t[63] = t[157] ^ t[93];
  assign t[64] = t[158] ^ t[94];
  assign t[65] = ~(t[71]);
  assign t[66] = ~(t[95]);
  assign t[67] = ~(t[23]);
  assign t[68] = t[96];
  assign t[69] = t[13] ^ t[95];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[95] ^ t[24];
  assign t[71] = t[68] ^ t[23];
  assign t[72] = ~(t[74] & t[97]);
  assign t[73] = ~(t[165] ^ t[98]);
  assign t[74] = ~(t[99] & t[100]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[166]);
  assign t[77] = t[162] ^ t[101];
  assign t[78] = t[163] ^ t[102];
  assign t[79] = t[103] & t[104];
  assign t[7] = t[13] ^ t[14];
  assign t[80] = t[105] & t[106];
  assign t[81] = ~(t[79] ^ t[107]);
  assign t[82] = t[108] ^ t[109];
  assign t[83] = t[75] ? x[50] : x[49];
  assign t[84] = t[110] & t[111];
  assign t[85] = t[112] & t[113];
  assign t[86] = ~(t[114] ^ t[56]);
  assign t[87] = t[115] ^ t[113];
  assign t[88] = t[164] ^ t[116];
  assign t[89] = t[117] & t[118];
  assign t[8] = ~(t[15]);
  assign t[90] = t[119] & t[61];
  assign t[91] = t[161] ^ t[120];
  assign t[92] = t[8] ? t[121] : t[167];
  assign t[93] = t[122] ? x[55] : x[54];
  assign t[94] = t[122] ? x[57] : x[56];
  assign t[95] = t[123];
  assign t[96] = t[27] ? t[124] : t[168];
  assign t[97] = ~(t[125] & t[126]);
  assign t[98] = t[127] ^ t[169];
  assign t[99] = ~(t[165]);
  assign t[9] = t[152] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [111:0] x;
 output y;

 wire [323:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[116] ^ t[117];
  assign t[101] = t[117] ^ t[25];
  assign t[102] = ~(t[119] & t[120]);
  assign t[103] = t[121] ^ t[159];
  assign t[104] = ~(t[156]);
  assign t[105] = t[122] & t[121];
  assign t[106] = t[8] ? t[123] : t[160];
  assign t[107] = t[158] ^ t[124];
  assign t[108] = ~(t[48]);
  assign t[109] = t[108] ? x[74] : x[73];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[48]);
  assign t[111] = t[92] ^ t[113];
  assign t[112] = t[56] ? t[125] : t[161];
  assign t[113] = t[146] ^ t[126];
  assign t[114] = t[56] ? t[127] : t[162];
  assign t[115] = t[99] ^ t[117];
  assign t[116] = t[128];
  assign t[117] = ~t[129];
  assign t[118] = t[56] ? t[130] : t[163];
  assign t[119] = ~(t[122] | t[121]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[131] | t[104]);
  assign t[121] = ~(t[164]);
  assign t[122] = ~(t[159]);
  assign t[123] = t[160] ^ t[132];
  assign t[124] = t[28] ? x[88] : x[87];
  assign t[125] = t[161] ^ t[133];
  assign t[126] = t[56] ? t[134] : t[165];
  assign t[127] = t[162] ^ t[135];
  assign t[128] = t[56] ? t[136] : t[166];
  assign t[129] = t[56] ? t[137] : t[167];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[163] ^ t[138];
  assign t[131] = ~(t[153]);
  assign t[132] = t[28] ? x[99] : x[98];
  assign t[133] = t[110] ? x[101] : x[100];
  assign t[134] = t[165] ^ t[139];
  assign t[135] = t[110] ? x[103] : x[102];
  assign t[136] = t[166] ^ t[140];
  assign t[137] = t[167] ^ t[141];
  assign t[138] = t[74] ? x[105] : x[104];
  assign t[139] = t[110] ? x[107] : x[106];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[74] ? x[109] : x[108];
  assign t[141] = t[110] ? x[111] : x[110];
  assign t[142] = (t[168]);
  assign t[143] = (t[169]);
  assign t[144] = (t[170]);
  assign t[145] = (t[171]);
  assign t[146] = (t[172]);
  assign t[147] = (t[173]);
  assign t[148] = (t[174]);
  assign t[149] = (t[175]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = (t[176]);
  assign t[151] = (t[177]);
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = t[194] ^ x[4];
  assign t[169] = t[195] ^ x[9];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[196] ^ x[12];
  assign t[171] = t[197] ^ x[15];
  assign t[172] = t[198] ^ x[18];
  assign t[173] = t[199] ^ x[21];
  assign t[174] = t[200] ^ x[24];
  assign t[175] = t[201] ^ x[27];
  assign t[176] = t[202] ^ x[30];
  assign t[177] = t[203] ^ x[33];
  assign t[178] = t[204] ^ x[36];
  assign t[179] = t[205] ^ x[39];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[42];
  assign t[181] = t[207] ^ x[45];
  assign t[182] = t[208] ^ x[48];
  assign t[183] = t[209] ^ x[51];
  assign t[184] = t[210] ^ x[56];
  assign t[185] = t[211] ^ x[69];
  assign t[186] = t[212] ^ x[72];
  assign t[187] = t[213] ^ x[77];
  assign t[188] = t[214] ^ x[80];
  assign t[189] = t[215] ^ x[83];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[86];
  assign t[191] = t[217] ^ x[91];
  assign t[192] = t[218] ^ x[94];
  assign t[193] = t[219] ^ x[97];
  assign t[194] = (t[220] & ~t[221]);
  assign t[195] = (t[222] & ~t[223]);
  assign t[196] = (t[224] & ~t[225]);
  assign t[197] = (t[226] & ~t[227]);
  assign t[198] = (t[228] & ~t[229]);
  assign t[199] = (t[230] & ~t[231]);
  assign t[19] = t[33] ^ t[4];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[232] & ~t[233]);
  assign t[201] = (t[234] & ~t[235]);
  assign t[202] = (t[236] & ~t[237]);
  assign t[203] = (t[238] & ~t[239]);
  assign t[204] = (t[240] & ~t[241]);
  assign t[205] = (t[242] & ~t[243]);
  assign t[206] = (t[244] & ~t[245]);
  assign t[207] = (t[246] & ~t[247]);
  assign t[208] = (t[248] & ~t[249]);
  assign t[209] = (t[250] & ~t[251]);
  assign t[20] = t[34] ^ t[35];
  assign t[210] = (t[252] & ~t[253]);
  assign t[211] = (t[254] & ~t[255]);
  assign t[212] = (t[256] & ~t[257]);
  assign t[213] = (t[258] & ~t[259]);
  assign t[214] = (t[260] & ~t[261]);
  assign t[215] = (t[262] & ~t[263]);
  assign t[216] = (t[264] & ~t[265]);
  assign t[217] = (t[266] & ~t[267]);
  assign t[218] = (t[268] & ~t[269]);
  assign t[219] = (t[270] & ~t[271]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = t[272] ^ x[4];
  assign t[221] = t[273] ^ x[3];
  assign t[222] = t[274] ^ x[9];
  assign t[223] = t[275] ^ x[8];
  assign t[224] = t[276] ^ x[12];
  assign t[225] = t[277] ^ x[11];
  assign t[226] = t[278] ^ x[15];
  assign t[227] = t[279] ^ x[14];
  assign t[228] = t[280] ^ x[18];
  assign t[229] = t[281] ^ x[17];
  assign t[22] = t[38] & t[39];
  assign t[230] = t[282] ^ x[21];
  assign t[231] = t[283] ^ x[20];
  assign t[232] = t[284] ^ x[24];
  assign t[233] = t[285] ^ x[23];
  assign t[234] = t[286] ^ x[27];
  assign t[235] = t[287] ^ x[26];
  assign t[236] = t[288] ^ x[30];
  assign t[237] = t[289] ^ x[29];
  assign t[238] = t[290] ^ x[33];
  assign t[239] = t[291] ^ x[32];
  assign t[23] = t[143] ^ t[40];
  assign t[240] = t[292] ^ x[36];
  assign t[241] = t[293] ^ x[35];
  assign t[242] = t[294] ^ x[39];
  assign t[243] = t[295] ^ x[38];
  assign t[244] = t[296] ^ x[42];
  assign t[245] = t[297] ^ x[41];
  assign t[246] = t[298] ^ x[45];
  assign t[247] = t[299] ^ x[44];
  assign t[248] = t[300] ^ x[48];
  assign t[249] = t[301] ^ x[47];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[302] ^ x[51];
  assign t[251] = t[303] ^ x[50];
  assign t[252] = t[304] ^ x[56];
  assign t[253] = t[305] ^ x[55];
  assign t[254] = t[306] ^ x[69];
  assign t[255] = t[307] ^ x[68];
  assign t[256] = t[308] ^ x[72];
  assign t[257] = t[309] ^ x[71];
  assign t[258] = t[310] ^ x[77];
  assign t[259] = t[311] ^ x[76];
  assign t[25] = t[43];
  assign t[260] = t[312] ^ x[80];
  assign t[261] = t[313] ^ x[79];
  assign t[262] = t[314] ^ x[83];
  assign t[263] = t[315] ^ x[82];
  assign t[264] = t[316] ^ x[86];
  assign t[265] = t[317] ^ x[85];
  assign t[266] = t[318] ^ x[91];
  assign t[267] = t[319] ^ x[90];
  assign t[268] = t[320] ^ x[94];
  assign t[269] = t[321] ^ x[93];
  assign t[26] = t[44] ^ t[45];
  assign t[270] = t[322] ^ x[97];
  assign t[271] = t[323] ^ x[96];
  assign t[272] = (x[2]);
  assign t[273] = (x[2]);
  assign t[274] = (x[7]);
  assign t[275] = (x[7]);
  assign t[276] = (x[10]);
  assign t[277] = (x[10]);
  assign t[278] = (x[13]);
  assign t[279] = (x[13]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (x[16]);
  assign t[281] = (x[16]);
  assign t[282] = (x[19]);
  assign t[283] = (x[19]);
  assign t[284] = (x[22]);
  assign t[285] = (x[22]);
  assign t[286] = (x[25]);
  assign t[287] = (x[25]);
  assign t[288] = (x[28]);
  assign t[289] = (x[28]);
  assign t[28] = ~(t[48]);
  assign t[290] = (x[31]);
  assign t[291] = (x[31]);
  assign t[292] = (x[34]);
  assign t[293] = (x[34]);
  assign t[294] = (x[37]);
  assign t[295] = (x[37]);
  assign t[296] = (x[40]);
  assign t[297] = (x[40]);
  assign t[298] = (x[43]);
  assign t[299] = (x[43]);
  assign t[29] = ~(t[144]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[46]);
  assign t[301] = (x[46]);
  assign t[302] = (x[49]);
  assign t[303] = (x[49]);
  assign t[304] = (x[54]);
  assign t[305] = (x[54]);
  assign t[306] = (x[67]);
  assign t[307] = (x[67]);
  assign t[308] = (x[70]);
  assign t[309] = (x[70]);
  assign t[30] = ~(t[145]);
  assign t[310] = (x[75]);
  assign t[311] = (x[75]);
  assign t[312] = (x[78]);
  assign t[313] = (x[78]);
  assign t[314] = (x[81]);
  assign t[315] = (x[81]);
  assign t[316] = (x[84]);
  assign t[317] = (x[84]);
  assign t[318] = (x[89]);
  assign t[319] = (x[89]);
  assign t[31] = ~(t[146]);
  assign t[320] = (x[92]);
  assign t[321] = (x[92]);
  assign t[322] = (x[95]);
  assign t[323] = (x[95]);
  assign t[32] = ~(t[49] | t[50]);
  assign t[33] = t[8] ? t[51] : t[147];
  assign t[34] = t[52] ^ t[53];
  assign t[35] = t[54] & t[55];
  assign t[36] = t[56] ? t[57] : t[148];
  assign t[37] = t[56] ? t[58] : t[149];
  assign t[38] = ~(t[59]);
  assign t[39] = t[56] ? t[60] : t[150];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[56] ? t[61] : t[151];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] & t[65];
  assign t[43] = t[56] ? t[66] : t[152];
  assign t[44] = t[67] ^ t[68];
  assign t[45] = t[69] & t[70];
  assign t[46] = ~(t[71] & t[72]);
  assign t[47] = t[153] | t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = ~(t[143]);
  assign t[4] = t[8] ? t[9] : t[142];
  assign t[50] = ~(t[75] & t[154]);
  assign t[51] = t[147] ^ t[76];
  assign t[52] = t[77] & t[78];
  assign t[53] = t[79] & t[80];
  assign t[54] = ~(t[52] ^ t[81]);
  assign t[55] = t[82] ^ t[83];
  assign t[56] = ~(t[15]);
  assign t[57] = t[148] ^ t[84];
  assign t[58] = t[149] ^ t[85];
  assign t[59] = t[56] ? t[86] : t[155];
  assign t[5] = ~(t[10]);
  assign t[60] = t[150] ^ t[87];
  assign t[61] = t[151] ^ t[88];
  assign t[62] = t[89] & t[90];
  assign t[63] = t[91] & t[92];
  assign t[64] = ~(t[93] ^ t[41]);
  assign t[65] = t[94] ^ t[92];
  assign t[66] = t[152] ^ t[95];
  assign t[67] = t[96] & t[97];
  assign t[68] = t[98] & t[99];
  assign t[69] = ~(t[100] ^ t[44]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[101] ^ t[99];
  assign t[71] = ~(t[73] & t[102]);
  assign t[72] = ~(t[156] ^ t[103]);
  assign t[73] = ~(t[104] & t[105]);
  assign t[74] = ~(t[47]);
  assign t[75] = ~(t[157]);
  assign t[76] = t[28] ? x[53] : x[52];
  assign t[77] = ~(t[83]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[33]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[107] : t[158];
  assign t[81] = t[19] ^ t[106];
  assign t[82] = t[106] ^ t[4];
  assign t[83] = t[80] ^ t[33];
  assign t[84] = t[108] ? x[58] : x[57];
  assign t[85] = t[74] ? x[60] : x[59];
  assign t[86] = t[155] ^ t[109];
  assign t[87] = t[108] ? x[62] : x[61];
  assign t[88] = t[110] ? x[64] : x[63];
  assign t[89] = ~(t[111]);
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[112]);
  assign t[91] = ~(t[113]);
  assign t[92] = t[157] ^ t[114];
  assign t[93] = t[112] ^ t[113];
  assign t[94] = t[113] ^ t[23];
  assign t[95] = t[74] ? x[66] : x[65];
  assign t[96] = ~(t[115]);
  assign t[97] = ~(t[116]);
  assign t[98] = ~(t[117]);
  assign t[99] = t[118];
  assign t[9] = t[142] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind41(x, y);
 input [111:0] x;
 output y;

 wire [323:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[116] ^ t[117];
  assign t[101] = t[117] ^ t[25];
  assign t[102] = ~(t[119] & t[120]);
  assign t[103] = t[121] ^ t[159];
  assign t[104] = ~(t[156]);
  assign t[105] = t[122] & t[121];
  assign t[106] = t[8] ? t[123] : t[160];
  assign t[107] = t[158] ^ t[124];
  assign t[108] = ~(t[48]);
  assign t[109] = t[108] ? x[74] : x[73];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[48]);
  assign t[111] = t[92] ^ t[113];
  assign t[112] = t[56] ? t[125] : t[161];
  assign t[113] = t[146] ^ t[126];
  assign t[114] = t[56] ? t[127] : t[162];
  assign t[115] = t[99] ^ t[117];
  assign t[116] = t[128];
  assign t[117] = ~t[129];
  assign t[118] = t[56] ? t[130] : t[163];
  assign t[119] = ~(t[122] | t[121]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[131] | t[104]);
  assign t[121] = ~(t[164]);
  assign t[122] = ~(t[159]);
  assign t[123] = t[160] ^ t[132];
  assign t[124] = t[28] ? x[88] : x[87];
  assign t[125] = t[161] ^ t[133];
  assign t[126] = t[56] ? t[134] : t[165];
  assign t[127] = t[162] ^ t[135];
  assign t[128] = t[56] ? t[136] : t[166];
  assign t[129] = t[56] ? t[137] : t[167];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[163] ^ t[138];
  assign t[131] = ~(t[153]);
  assign t[132] = t[28] ? x[99] : x[98];
  assign t[133] = t[110] ? x[101] : x[100];
  assign t[134] = t[165] ^ t[139];
  assign t[135] = t[110] ? x[103] : x[102];
  assign t[136] = t[166] ^ t[140];
  assign t[137] = t[167] ^ t[141];
  assign t[138] = t[74] ? x[105] : x[104];
  assign t[139] = t[110] ? x[107] : x[106];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[74] ? x[109] : x[108];
  assign t[141] = t[110] ? x[111] : x[110];
  assign t[142] = (t[168]);
  assign t[143] = (t[169]);
  assign t[144] = (t[170]);
  assign t[145] = (t[171]);
  assign t[146] = (t[172]);
  assign t[147] = (t[173]);
  assign t[148] = (t[174]);
  assign t[149] = (t[175]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = (t[176]);
  assign t[151] = (t[177]);
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = t[194] ^ x[4];
  assign t[169] = t[195] ^ x[9];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[196] ^ x[12];
  assign t[171] = t[197] ^ x[15];
  assign t[172] = t[198] ^ x[18];
  assign t[173] = t[199] ^ x[21];
  assign t[174] = t[200] ^ x[24];
  assign t[175] = t[201] ^ x[27];
  assign t[176] = t[202] ^ x[30];
  assign t[177] = t[203] ^ x[33];
  assign t[178] = t[204] ^ x[36];
  assign t[179] = t[205] ^ x[39];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[42];
  assign t[181] = t[207] ^ x[45];
  assign t[182] = t[208] ^ x[48];
  assign t[183] = t[209] ^ x[51];
  assign t[184] = t[210] ^ x[56];
  assign t[185] = t[211] ^ x[69];
  assign t[186] = t[212] ^ x[72];
  assign t[187] = t[213] ^ x[77];
  assign t[188] = t[214] ^ x[80];
  assign t[189] = t[215] ^ x[83];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[86];
  assign t[191] = t[217] ^ x[91];
  assign t[192] = t[218] ^ x[94];
  assign t[193] = t[219] ^ x[97];
  assign t[194] = (t[220] & ~t[221]);
  assign t[195] = (t[222] & ~t[223]);
  assign t[196] = (t[224] & ~t[225]);
  assign t[197] = (t[226] & ~t[227]);
  assign t[198] = (t[228] & ~t[229]);
  assign t[199] = (t[230] & ~t[231]);
  assign t[19] = t[33] ^ t[4];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[232] & ~t[233]);
  assign t[201] = (t[234] & ~t[235]);
  assign t[202] = (t[236] & ~t[237]);
  assign t[203] = (t[238] & ~t[239]);
  assign t[204] = (t[240] & ~t[241]);
  assign t[205] = (t[242] & ~t[243]);
  assign t[206] = (t[244] & ~t[245]);
  assign t[207] = (t[246] & ~t[247]);
  assign t[208] = (t[248] & ~t[249]);
  assign t[209] = (t[250] & ~t[251]);
  assign t[20] = t[34] ^ t[35];
  assign t[210] = (t[252] & ~t[253]);
  assign t[211] = (t[254] & ~t[255]);
  assign t[212] = (t[256] & ~t[257]);
  assign t[213] = (t[258] & ~t[259]);
  assign t[214] = (t[260] & ~t[261]);
  assign t[215] = (t[262] & ~t[263]);
  assign t[216] = (t[264] & ~t[265]);
  assign t[217] = (t[266] & ~t[267]);
  assign t[218] = (t[268] & ~t[269]);
  assign t[219] = (t[270] & ~t[271]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = t[272] ^ x[4];
  assign t[221] = t[273] ^ x[3];
  assign t[222] = t[274] ^ x[9];
  assign t[223] = t[275] ^ x[8];
  assign t[224] = t[276] ^ x[12];
  assign t[225] = t[277] ^ x[11];
  assign t[226] = t[278] ^ x[15];
  assign t[227] = t[279] ^ x[14];
  assign t[228] = t[280] ^ x[18];
  assign t[229] = t[281] ^ x[17];
  assign t[22] = t[38] & t[39];
  assign t[230] = t[282] ^ x[21];
  assign t[231] = t[283] ^ x[20];
  assign t[232] = t[284] ^ x[24];
  assign t[233] = t[285] ^ x[23];
  assign t[234] = t[286] ^ x[27];
  assign t[235] = t[287] ^ x[26];
  assign t[236] = t[288] ^ x[30];
  assign t[237] = t[289] ^ x[29];
  assign t[238] = t[290] ^ x[33];
  assign t[239] = t[291] ^ x[32];
  assign t[23] = t[143] ^ t[40];
  assign t[240] = t[292] ^ x[36];
  assign t[241] = t[293] ^ x[35];
  assign t[242] = t[294] ^ x[39];
  assign t[243] = t[295] ^ x[38];
  assign t[244] = t[296] ^ x[42];
  assign t[245] = t[297] ^ x[41];
  assign t[246] = t[298] ^ x[45];
  assign t[247] = t[299] ^ x[44];
  assign t[248] = t[300] ^ x[48];
  assign t[249] = t[301] ^ x[47];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[302] ^ x[51];
  assign t[251] = t[303] ^ x[50];
  assign t[252] = t[304] ^ x[56];
  assign t[253] = t[305] ^ x[55];
  assign t[254] = t[306] ^ x[69];
  assign t[255] = t[307] ^ x[68];
  assign t[256] = t[308] ^ x[72];
  assign t[257] = t[309] ^ x[71];
  assign t[258] = t[310] ^ x[77];
  assign t[259] = t[311] ^ x[76];
  assign t[25] = t[43];
  assign t[260] = t[312] ^ x[80];
  assign t[261] = t[313] ^ x[79];
  assign t[262] = t[314] ^ x[83];
  assign t[263] = t[315] ^ x[82];
  assign t[264] = t[316] ^ x[86];
  assign t[265] = t[317] ^ x[85];
  assign t[266] = t[318] ^ x[91];
  assign t[267] = t[319] ^ x[90];
  assign t[268] = t[320] ^ x[94];
  assign t[269] = t[321] ^ x[93];
  assign t[26] = t[44] ^ t[45];
  assign t[270] = t[322] ^ x[97];
  assign t[271] = t[323] ^ x[96];
  assign t[272] = (x[2]);
  assign t[273] = (x[2]);
  assign t[274] = (x[7]);
  assign t[275] = (x[7]);
  assign t[276] = (x[10]);
  assign t[277] = (x[10]);
  assign t[278] = (x[13]);
  assign t[279] = (x[13]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (x[16]);
  assign t[281] = (x[16]);
  assign t[282] = (x[19]);
  assign t[283] = (x[19]);
  assign t[284] = (x[22]);
  assign t[285] = (x[22]);
  assign t[286] = (x[25]);
  assign t[287] = (x[25]);
  assign t[288] = (x[28]);
  assign t[289] = (x[28]);
  assign t[28] = ~(t[48]);
  assign t[290] = (x[31]);
  assign t[291] = (x[31]);
  assign t[292] = (x[34]);
  assign t[293] = (x[34]);
  assign t[294] = (x[37]);
  assign t[295] = (x[37]);
  assign t[296] = (x[40]);
  assign t[297] = (x[40]);
  assign t[298] = (x[43]);
  assign t[299] = (x[43]);
  assign t[29] = ~(t[144]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[46]);
  assign t[301] = (x[46]);
  assign t[302] = (x[49]);
  assign t[303] = (x[49]);
  assign t[304] = (x[54]);
  assign t[305] = (x[54]);
  assign t[306] = (x[67]);
  assign t[307] = (x[67]);
  assign t[308] = (x[70]);
  assign t[309] = (x[70]);
  assign t[30] = ~(t[145]);
  assign t[310] = (x[75]);
  assign t[311] = (x[75]);
  assign t[312] = (x[78]);
  assign t[313] = (x[78]);
  assign t[314] = (x[81]);
  assign t[315] = (x[81]);
  assign t[316] = (x[84]);
  assign t[317] = (x[84]);
  assign t[318] = (x[89]);
  assign t[319] = (x[89]);
  assign t[31] = ~(t[146]);
  assign t[320] = (x[92]);
  assign t[321] = (x[92]);
  assign t[322] = (x[95]);
  assign t[323] = (x[95]);
  assign t[32] = ~(t[49] | t[50]);
  assign t[33] = t[8] ? t[51] : t[147];
  assign t[34] = t[52] ^ t[53];
  assign t[35] = t[54] & t[55];
  assign t[36] = t[56] ? t[57] : t[148];
  assign t[37] = t[56] ? t[58] : t[149];
  assign t[38] = ~(t[59]);
  assign t[39] = t[56] ? t[60] : t[150];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[56] ? t[61] : t[151];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] & t[65];
  assign t[43] = t[56] ? t[66] : t[152];
  assign t[44] = t[67] ^ t[68];
  assign t[45] = t[69] & t[70];
  assign t[46] = ~(t[71] & t[72]);
  assign t[47] = t[153] | t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = ~(t[143]);
  assign t[4] = t[8] ? t[9] : t[142];
  assign t[50] = ~(t[75] & t[154]);
  assign t[51] = t[147] ^ t[76];
  assign t[52] = t[77] & t[78];
  assign t[53] = t[79] & t[80];
  assign t[54] = ~(t[52] ^ t[81]);
  assign t[55] = t[82] ^ t[83];
  assign t[56] = ~(t[15]);
  assign t[57] = t[148] ^ t[84];
  assign t[58] = t[149] ^ t[85];
  assign t[59] = t[56] ? t[86] : t[155];
  assign t[5] = ~(t[10]);
  assign t[60] = t[150] ^ t[87];
  assign t[61] = t[151] ^ t[88];
  assign t[62] = t[89] & t[90];
  assign t[63] = t[91] & t[92];
  assign t[64] = ~(t[93] ^ t[41]);
  assign t[65] = t[94] ^ t[92];
  assign t[66] = t[152] ^ t[95];
  assign t[67] = t[96] & t[97];
  assign t[68] = t[98] & t[99];
  assign t[69] = ~(t[100] ^ t[44]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[101] ^ t[99];
  assign t[71] = ~(t[73] & t[102]);
  assign t[72] = ~(t[156] ^ t[103]);
  assign t[73] = ~(t[104] & t[105]);
  assign t[74] = ~(t[47]);
  assign t[75] = ~(t[157]);
  assign t[76] = t[28] ? x[53] : x[52];
  assign t[77] = ~(t[83]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[33]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[107] : t[158];
  assign t[81] = t[19] ^ t[106];
  assign t[82] = t[106] ^ t[4];
  assign t[83] = t[80] ^ t[33];
  assign t[84] = t[108] ? x[58] : x[57];
  assign t[85] = t[74] ? x[60] : x[59];
  assign t[86] = t[155] ^ t[109];
  assign t[87] = t[108] ? x[62] : x[61];
  assign t[88] = t[110] ? x[64] : x[63];
  assign t[89] = ~(t[111]);
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[112]);
  assign t[91] = ~(t[113]);
  assign t[92] = t[157] ^ t[114];
  assign t[93] = t[112] ^ t[113];
  assign t[94] = t[113] ^ t[23];
  assign t[95] = t[74] ? x[66] : x[65];
  assign t[96] = ~(t[115]);
  assign t[97] = ~(t[116]);
  assign t[98] = ~(t[117]);
  assign t[99] = t[118];
  assign t[9] = t[142] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind42(x, y);
 input [111:0] x;
 output y;

 wire [345:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[41] ^ t[65];
  assign t[101] = t[65] ^ t[25];
  assign t[102] = ~(t[133] & t[134]);
  assign t[103] = t[135] ^ t[183];
  assign t[104] = ~(t[178]);
  assign t[105] = t[136] & t[135];
  assign t[106] = t[137] ? x[67] : x[66];
  assign t[107] = ~(t[138]);
  assign t[108] = ~(t[55]);
  assign t[109] = t[55] ^ t[82];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[82] ^ t[33];
  assign t[111] = t[137] ? x[69] : x[68];
  assign t[112] = t[67] ? t[139] : t[184];
  assign t[113] = t[179] ^ t[140];
  assign t[114] = t[180] ^ t[141];
  assign t[115] = t[181] ^ t[142];
  assign t[116] = t[143] ^ t[144];
  assign t[117] = t[85] ^ t[145];
  assign t[118] = t[67] ? t[146] : t[185];
  assign t[119] = t[28] ? x[77] : x[76];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[147] ^ t[62]);
  assign t[121] = t[39] ^ t[125];
  assign t[122] = ~(t[128]);
  assign t[123] = ~(t[148]);
  assign t[124] = ~(t[4]);
  assign t[125] = t[8] ? t[149] : t[186];
  assign t[126] = t[39] ^ t[148];
  assign t[127] = t[148] ^ t[60];
  assign t[128] = t[125] ^ t[4];
  assign t[129] = t[75] ? x[82] : x[81];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[182] ^ t[150];
  assign t[131] = t[75] ? x[84] : x[83];
  assign t[132] = t[43] ^ t[65];
  assign t[133] = ~(t[136] | t[135]);
  assign t[134] = ~(t[151] | t[104]);
  assign t[135] = ~(t[187]);
  assign t[136] = ~(t[183]);
  assign t[137] = ~(t[49]);
  assign t[138] = t[57] ^ t[82];
  assign t[139] = t[184] ^ t[152];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[137] ? x[89] : x[88];
  assign t[141] = t[153] ? x[91] : x[90];
  assign t[142] = t[153] ? x[93] : x[92];
  assign t[143] = t[154] & t[155];
  assign t[144] = t[156] & t[118];
  assign t[145] = t[67] ? t[157] : t[188];
  assign t[146] = t[185] ^ t[158];
  assign t[147] = t[148] ^ t[4];
  assign t[148] = t[8] ? t[159] : t[189];
  assign t[149] = t[186] ^ t[160];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[137] ? x[101] : x[100];
  assign t[151] = ~(t[170]);
  assign t[152] = t[137] ? x[103] : x[102];
  assign t[153] = ~(t[49]);
  assign t[154] = ~(t[161]);
  assign t[155] = ~(t[84]);
  assign t[156] = ~(t[85]);
  assign t[157] = t[188] ^ t[162];
  assign t[158] = t[153] ? x[105] : x[104];
  assign t[159] = t[189] ^ t[163];
  assign t[15] = ~(t[27]);
  assign t[160] = t[28] ? x[107] : x[106];
  assign t[161] = t[118] ^ t[85];
  assign t[162] = t[75] ? x[109] : x[108];
  assign t[163] = t[28] ? x[111] : x[110];
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = (t[205]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[206]);
  assign t[181] = (t[207]);
  assign t[182] = (t[208]);
  assign t[183] = (t[209]);
  assign t[184] = (t[210]);
  assign t[185] = (t[211]);
  assign t[186] = (t[212]);
  assign t[187] = (t[213]);
  assign t[188] = (t[214]);
  assign t[189] = (t[215]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[4];
  assign t[191] = t[217] ^ x[9];
  assign t[192] = t[218] ^ x[12];
  assign t[193] = t[219] ^ x[15];
  assign t[194] = t[220] ^ x[18];
  assign t[195] = t[221] ^ x[21];
  assign t[196] = t[222] ^ x[24];
  assign t[197] = t[223] ^ x[27];
  assign t[198] = t[224] ^ x[30];
  assign t[199] = t[225] ^ x[33];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[36];
  assign t[201] = t[227] ^ x[39];
  assign t[202] = t[228] ^ x[42];
  assign t[203] = t[229] ^ x[45];
  assign t[204] = t[230] ^ x[48];
  assign t[205] = t[231] ^ x[51];
  assign t[206] = t[232] ^ x[54];
  assign t[207] = t[233] ^ x[57];
  assign t[208] = t[234] ^ x[60];
  assign t[209] = t[235] ^ x[65];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[236] ^ x[72];
  assign t[211] = t[237] ^ x[75];
  assign t[212] = t[238] ^ x[80];
  assign t[213] = t[239] ^ x[87];
  assign t[214] = t[240] ^ x[96];
  assign t[215] = t[241] ^ x[99];
  assign t[216] = (t[242] & ~t[243]);
  assign t[217] = (t[244] & ~t[245]);
  assign t[218] = (t[246] & ~t[247]);
  assign t[219] = (t[248] & ~t[249]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[250] & ~t[251]);
  assign t[221] = (t[252] & ~t[253]);
  assign t[222] = (t[254] & ~t[255]);
  assign t[223] = (t[256] & ~t[257]);
  assign t[224] = (t[258] & ~t[259]);
  assign t[225] = (t[260] & ~t[261]);
  assign t[226] = (t[262] & ~t[263]);
  assign t[227] = (t[264] & ~t[265]);
  assign t[228] = (t[266] & ~t[267]);
  assign t[229] = (t[268] & ~t[269]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[270] & ~t[271]);
  assign t[231] = (t[272] & ~t[273]);
  assign t[232] = (t[274] & ~t[275]);
  assign t[233] = (t[276] & ~t[277]);
  assign t[234] = (t[278] & ~t[279]);
  assign t[235] = (t[280] & ~t[281]);
  assign t[236] = (t[282] & ~t[283]);
  assign t[237] = (t[284] & ~t[285]);
  assign t[238] = (t[286] & ~t[287]);
  assign t[239] = (t[288] & ~t[289]);
  assign t[23] = t[41] ^ t[25];
  assign t[240] = (t[290] & ~t[291]);
  assign t[241] = (t[292] & ~t[293]);
  assign t[242] = t[294] ^ x[4];
  assign t[243] = t[295] ^ x[3];
  assign t[244] = t[296] ^ x[9];
  assign t[245] = t[297] ^ x[8];
  assign t[246] = t[298] ^ x[12];
  assign t[247] = t[299] ^ x[11];
  assign t[248] = t[300] ^ x[15];
  assign t[249] = t[301] ^ x[14];
  assign t[24] = t[42] & t[43];
  assign t[250] = t[302] ^ x[18];
  assign t[251] = t[303] ^ x[17];
  assign t[252] = t[304] ^ x[21];
  assign t[253] = t[305] ^ x[20];
  assign t[254] = t[306] ^ x[24];
  assign t[255] = t[307] ^ x[23];
  assign t[256] = t[308] ^ x[27];
  assign t[257] = t[309] ^ x[26];
  assign t[258] = t[310] ^ x[30];
  assign t[259] = t[311] ^ x[29];
  assign t[25] = t[44];
  assign t[260] = t[312] ^ x[33];
  assign t[261] = t[313] ^ x[32];
  assign t[262] = t[314] ^ x[36];
  assign t[263] = t[315] ^ x[35];
  assign t[264] = t[316] ^ x[39];
  assign t[265] = t[317] ^ x[38];
  assign t[266] = t[318] ^ x[42];
  assign t[267] = t[319] ^ x[41];
  assign t[268] = t[320] ^ x[45];
  assign t[269] = t[321] ^ x[44];
  assign t[26] = t[45] ^ t[46];
  assign t[270] = t[322] ^ x[48];
  assign t[271] = t[323] ^ x[47];
  assign t[272] = t[324] ^ x[51];
  assign t[273] = t[325] ^ x[50];
  assign t[274] = t[326] ^ x[54];
  assign t[275] = t[327] ^ x[53];
  assign t[276] = t[328] ^ x[57];
  assign t[277] = t[329] ^ x[56];
  assign t[278] = t[330] ^ x[60];
  assign t[279] = t[331] ^ x[59];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[332] ^ x[65];
  assign t[281] = t[333] ^ x[64];
  assign t[282] = t[334] ^ x[72];
  assign t[283] = t[335] ^ x[71];
  assign t[284] = t[336] ^ x[75];
  assign t[285] = t[337] ^ x[74];
  assign t[286] = t[338] ^ x[80];
  assign t[287] = t[339] ^ x[79];
  assign t[288] = t[340] ^ x[87];
  assign t[289] = t[341] ^ x[86];
  assign t[28] = ~(t[49]);
  assign t[290] = t[342] ^ x[96];
  assign t[291] = t[343] ^ x[95];
  assign t[292] = t[344] ^ x[99];
  assign t[293] = t[345] ^ x[98];
  assign t[294] = (x[2]);
  assign t[295] = (x[2]);
  assign t[296] = (x[7]);
  assign t[297] = (x[7]);
  assign t[298] = (x[10]);
  assign t[299] = (x[10]);
  assign t[29] = ~(t[165]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[13]);
  assign t[301] = (x[13]);
  assign t[302] = (x[16]);
  assign t[303] = (x[16]);
  assign t[304] = (x[19]);
  assign t[305] = (x[19]);
  assign t[306] = (x[22]);
  assign t[307] = (x[22]);
  assign t[308] = (x[25]);
  assign t[309] = (x[25]);
  assign t[30] = ~(t[166]);
  assign t[310] = (x[28]);
  assign t[311] = (x[28]);
  assign t[312] = (x[31]);
  assign t[313] = (x[31]);
  assign t[314] = (x[34]);
  assign t[315] = (x[34]);
  assign t[316] = (x[37]);
  assign t[317] = (x[37]);
  assign t[318] = (x[40]);
  assign t[319] = (x[40]);
  assign t[31] = ~(t[167]);
  assign t[320] = (x[43]);
  assign t[321] = (x[43]);
  assign t[322] = (x[46]);
  assign t[323] = (x[46]);
  assign t[324] = (x[49]);
  assign t[325] = (x[49]);
  assign t[326] = (x[52]);
  assign t[327] = (x[52]);
  assign t[328] = (x[55]);
  assign t[329] = (x[55]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[58]);
  assign t[331] = (x[58]);
  assign t[332] = (x[63]);
  assign t[333] = (x[63]);
  assign t[334] = (x[70]);
  assign t[335] = (x[70]);
  assign t[336] = (x[73]);
  assign t[337] = (x[73]);
  assign t[338] = (x[78]);
  assign t[339] = (x[78]);
  assign t[33] = t[168] ^ t[52];
  assign t[340] = (x[85]);
  assign t[341] = (x[85]);
  assign t[342] = (x[94]);
  assign t[343] = (x[94]);
  assign t[344] = (x[97]);
  assign t[345] = (x[97]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[55] ^ t[33];
  assign t[36] = t[56] & t[57];
  assign t[37] = t[58] ^ t[59];
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[4] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = t[64];
  assign t[42] = ~(t[65]);
  assign t[43] = t[66];
  assign t[44] = t[67] ? t[68] : t[169];
  assign t[45] = t[69] ^ t[24];
  assign t[46] = t[70] & t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[170] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = t[8] ? t[9] : t[164];
  assign t[50] = ~(t[168]);
  assign t[51] = ~(t[76] & t[171]);
  assign t[52] = t[67] ? t[77] : t[172];
  assign t[53] = t[78] ^ t[36];
  assign t[54] = t[79] & t[80];
  assign t[55] = t[67] ? t[81] : t[173];
  assign t[56] = ~(t[82]);
  assign t[57] = t[174] ^ t[83];
  assign t[58] = t[84] ^ t[85];
  assign t[59] = t[86] & t[87];
  assign t[5] = ~(t[10]);
  assign t[60] = t[8] ? t[88] : t[175];
  assign t[61] = t[62] ^ t[89];
  assign t[62] = t[90] ^ t[91];
  assign t[63] = t[92] & t[93];
  assign t[64] = t[67] ? t[94] : t[176];
  assign t[65] = ~t[95];
  assign t[66] = t[67] ? t[96] : t[177];
  assign t[67] = ~(t[15]);
  assign t[68] = t[169] ^ t[97];
  assign t[69] = t[98] & t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[100] ^ t[45]);
  assign t[71] = t[101] ^ t[43];
  assign t[72] = ~(t[74] & t[102]);
  assign t[73] = ~(t[178] ^ t[103]);
  assign t[74] = ~(t[104] & t[105]);
  assign t[75] = ~(t[48]);
  assign t[76] = ~(t[174]);
  assign t[77] = t[172] ^ t[106];
  assign t[78] = t[107] & t[108];
  assign t[79] = ~(t[109] ^ t[53]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[110] ^ t[57];
  assign t[81] = t[173] ^ t[111];
  assign t[82] = t[167] ^ t[112];
  assign t[83] = t[67] ? t[113] : t[179];
  assign t[84] = t[67] ? t[114] : t[180];
  assign t[85] = t[67] ? t[115] : t[181];
  assign t[86] = ~(t[58] ^ t[116]);
  assign t[87] = t[117] ^ t[118];
  assign t[88] = t[175] ^ t[119];
  assign t[89] = t[120] & t[121];
  assign t[8] = ~(t[15]);
  assign t[90] = t[122] & t[123];
  assign t[91] = t[124] & t[125];
  assign t[92] = ~(t[90] ^ t[126]);
  assign t[93] = t[127] ^ t[128];
  assign t[94] = t[176] ^ t[129];
  assign t[95] = t[67] ? t[130] : t[182];
  assign t[96] = t[177] ^ t[131];
  assign t[97] = t[75] ? x[62] : x[61];
  assign t[98] = ~(t[132]);
  assign t[99] = ~(t[41]);
  assign t[9] = t[164] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind43(x, y);
 input [111:0] x;
 output y;

 wire [345:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[41] ^ t[65];
  assign t[101] = t[65] ^ t[25];
  assign t[102] = ~(t[133] & t[134]);
  assign t[103] = t[135] ^ t[183];
  assign t[104] = ~(t[178]);
  assign t[105] = t[136] & t[135];
  assign t[106] = t[137] ? x[67] : x[66];
  assign t[107] = ~(t[138]);
  assign t[108] = ~(t[55]);
  assign t[109] = t[55] ^ t[82];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[82] ^ t[33];
  assign t[111] = t[137] ? x[69] : x[68];
  assign t[112] = t[67] ? t[139] : t[184];
  assign t[113] = t[179] ^ t[140];
  assign t[114] = t[180] ^ t[141];
  assign t[115] = t[181] ^ t[142];
  assign t[116] = t[143] ^ t[144];
  assign t[117] = t[85] ^ t[145];
  assign t[118] = t[67] ? t[146] : t[185];
  assign t[119] = t[28] ? x[77] : x[76];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[147] ^ t[62]);
  assign t[121] = t[39] ^ t[125];
  assign t[122] = ~(t[128]);
  assign t[123] = ~(t[148]);
  assign t[124] = ~(t[4]);
  assign t[125] = t[8] ? t[149] : t[186];
  assign t[126] = t[39] ^ t[148];
  assign t[127] = t[148] ^ t[60];
  assign t[128] = t[125] ^ t[4];
  assign t[129] = t[75] ? x[82] : x[81];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[182] ^ t[150];
  assign t[131] = t[75] ? x[84] : x[83];
  assign t[132] = t[43] ^ t[65];
  assign t[133] = ~(t[136] | t[135]);
  assign t[134] = ~(t[151] | t[104]);
  assign t[135] = ~(t[187]);
  assign t[136] = ~(t[183]);
  assign t[137] = ~(t[49]);
  assign t[138] = t[57] ^ t[82];
  assign t[139] = t[184] ^ t[152];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[137] ? x[89] : x[88];
  assign t[141] = t[153] ? x[91] : x[90];
  assign t[142] = t[153] ? x[93] : x[92];
  assign t[143] = t[154] & t[155];
  assign t[144] = t[156] & t[118];
  assign t[145] = t[67] ? t[157] : t[188];
  assign t[146] = t[185] ^ t[158];
  assign t[147] = t[148] ^ t[4];
  assign t[148] = t[8] ? t[159] : t[189];
  assign t[149] = t[186] ^ t[160];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[137] ? x[101] : x[100];
  assign t[151] = ~(t[170]);
  assign t[152] = t[137] ? x[103] : x[102];
  assign t[153] = ~(t[49]);
  assign t[154] = ~(t[161]);
  assign t[155] = ~(t[84]);
  assign t[156] = ~(t[85]);
  assign t[157] = t[188] ^ t[162];
  assign t[158] = t[153] ? x[105] : x[104];
  assign t[159] = t[189] ^ t[163];
  assign t[15] = ~(t[27]);
  assign t[160] = t[28] ? x[107] : x[106];
  assign t[161] = t[118] ^ t[85];
  assign t[162] = t[75] ? x[109] : x[108];
  assign t[163] = t[28] ? x[111] : x[110];
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = (t[205]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[206]);
  assign t[181] = (t[207]);
  assign t[182] = (t[208]);
  assign t[183] = (t[209]);
  assign t[184] = (t[210]);
  assign t[185] = (t[211]);
  assign t[186] = (t[212]);
  assign t[187] = (t[213]);
  assign t[188] = (t[214]);
  assign t[189] = (t[215]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[4];
  assign t[191] = t[217] ^ x[9];
  assign t[192] = t[218] ^ x[12];
  assign t[193] = t[219] ^ x[15];
  assign t[194] = t[220] ^ x[18];
  assign t[195] = t[221] ^ x[21];
  assign t[196] = t[222] ^ x[24];
  assign t[197] = t[223] ^ x[27];
  assign t[198] = t[224] ^ x[30];
  assign t[199] = t[225] ^ x[33];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[36];
  assign t[201] = t[227] ^ x[39];
  assign t[202] = t[228] ^ x[42];
  assign t[203] = t[229] ^ x[45];
  assign t[204] = t[230] ^ x[48];
  assign t[205] = t[231] ^ x[51];
  assign t[206] = t[232] ^ x[54];
  assign t[207] = t[233] ^ x[57];
  assign t[208] = t[234] ^ x[60];
  assign t[209] = t[235] ^ x[65];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[236] ^ x[72];
  assign t[211] = t[237] ^ x[75];
  assign t[212] = t[238] ^ x[80];
  assign t[213] = t[239] ^ x[87];
  assign t[214] = t[240] ^ x[96];
  assign t[215] = t[241] ^ x[99];
  assign t[216] = (t[242] & ~t[243]);
  assign t[217] = (t[244] & ~t[245]);
  assign t[218] = (t[246] & ~t[247]);
  assign t[219] = (t[248] & ~t[249]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[250] & ~t[251]);
  assign t[221] = (t[252] & ~t[253]);
  assign t[222] = (t[254] & ~t[255]);
  assign t[223] = (t[256] & ~t[257]);
  assign t[224] = (t[258] & ~t[259]);
  assign t[225] = (t[260] & ~t[261]);
  assign t[226] = (t[262] & ~t[263]);
  assign t[227] = (t[264] & ~t[265]);
  assign t[228] = (t[266] & ~t[267]);
  assign t[229] = (t[268] & ~t[269]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[270] & ~t[271]);
  assign t[231] = (t[272] & ~t[273]);
  assign t[232] = (t[274] & ~t[275]);
  assign t[233] = (t[276] & ~t[277]);
  assign t[234] = (t[278] & ~t[279]);
  assign t[235] = (t[280] & ~t[281]);
  assign t[236] = (t[282] & ~t[283]);
  assign t[237] = (t[284] & ~t[285]);
  assign t[238] = (t[286] & ~t[287]);
  assign t[239] = (t[288] & ~t[289]);
  assign t[23] = t[41] ^ t[25];
  assign t[240] = (t[290] & ~t[291]);
  assign t[241] = (t[292] & ~t[293]);
  assign t[242] = t[294] ^ x[4];
  assign t[243] = t[295] ^ x[3];
  assign t[244] = t[296] ^ x[9];
  assign t[245] = t[297] ^ x[8];
  assign t[246] = t[298] ^ x[12];
  assign t[247] = t[299] ^ x[11];
  assign t[248] = t[300] ^ x[15];
  assign t[249] = t[301] ^ x[14];
  assign t[24] = t[42] & t[43];
  assign t[250] = t[302] ^ x[18];
  assign t[251] = t[303] ^ x[17];
  assign t[252] = t[304] ^ x[21];
  assign t[253] = t[305] ^ x[20];
  assign t[254] = t[306] ^ x[24];
  assign t[255] = t[307] ^ x[23];
  assign t[256] = t[308] ^ x[27];
  assign t[257] = t[309] ^ x[26];
  assign t[258] = t[310] ^ x[30];
  assign t[259] = t[311] ^ x[29];
  assign t[25] = t[44];
  assign t[260] = t[312] ^ x[33];
  assign t[261] = t[313] ^ x[32];
  assign t[262] = t[314] ^ x[36];
  assign t[263] = t[315] ^ x[35];
  assign t[264] = t[316] ^ x[39];
  assign t[265] = t[317] ^ x[38];
  assign t[266] = t[318] ^ x[42];
  assign t[267] = t[319] ^ x[41];
  assign t[268] = t[320] ^ x[45];
  assign t[269] = t[321] ^ x[44];
  assign t[26] = t[45] ^ t[46];
  assign t[270] = t[322] ^ x[48];
  assign t[271] = t[323] ^ x[47];
  assign t[272] = t[324] ^ x[51];
  assign t[273] = t[325] ^ x[50];
  assign t[274] = t[326] ^ x[54];
  assign t[275] = t[327] ^ x[53];
  assign t[276] = t[328] ^ x[57];
  assign t[277] = t[329] ^ x[56];
  assign t[278] = t[330] ^ x[60];
  assign t[279] = t[331] ^ x[59];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[332] ^ x[65];
  assign t[281] = t[333] ^ x[64];
  assign t[282] = t[334] ^ x[72];
  assign t[283] = t[335] ^ x[71];
  assign t[284] = t[336] ^ x[75];
  assign t[285] = t[337] ^ x[74];
  assign t[286] = t[338] ^ x[80];
  assign t[287] = t[339] ^ x[79];
  assign t[288] = t[340] ^ x[87];
  assign t[289] = t[341] ^ x[86];
  assign t[28] = ~(t[49]);
  assign t[290] = t[342] ^ x[96];
  assign t[291] = t[343] ^ x[95];
  assign t[292] = t[344] ^ x[99];
  assign t[293] = t[345] ^ x[98];
  assign t[294] = (x[2]);
  assign t[295] = (x[2]);
  assign t[296] = (x[7]);
  assign t[297] = (x[7]);
  assign t[298] = (x[10]);
  assign t[299] = (x[10]);
  assign t[29] = ~(t[165]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[13]);
  assign t[301] = (x[13]);
  assign t[302] = (x[16]);
  assign t[303] = (x[16]);
  assign t[304] = (x[19]);
  assign t[305] = (x[19]);
  assign t[306] = (x[22]);
  assign t[307] = (x[22]);
  assign t[308] = (x[25]);
  assign t[309] = (x[25]);
  assign t[30] = ~(t[166]);
  assign t[310] = (x[28]);
  assign t[311] = (x[28]);
  assign t[312] = (x[31]);
  assign t[313] = (x[31]);
  assign t[314] = (x[34]);
  assign t[315] = (x[34]);
  assign t[316] = (x[37]);
  assign t[317] = (x[37]);
  assign t[318] = (x[40]);
  assign t[319] = (x[40]);
  assign t[31] = ~(t[167]);
  assign t[320] = (x[43]);
  assign t[321] = (x[43]);
  assign t[322] = (x[46]);
  assign t[323] = (x[46]);
  assign t[324] = (x[49]);
  assign t[325] = (x[49]);
  assign t[326] = (x[52]);
  assign t[327] = (x[52]);
  assign t[328] = (x[55]);
  assign t[329] = (x[55]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[58]);
  assign t[331] = (x[58]);
  assign t[332] = (x[63]);
  assign t[333] = (x[63]);
  assign t[334] = (x[70]);
  assign t[335] = (x[70]);
  assign t[336] = (x[73]);
  assign t[337] = (x[73]);
  assign t[338] = (x[78]);
  assign t[339] = (x[78]);
  assign t[33] = t[168] ^ t[52];
  assign t[340] = (x[85]);
  assign t[341] = (x[85]);
  assign t[342] = (x[94]);
  assign t[343] = (x[94]);
  assign t[344] = (x[97]);
  assign t[345] = (x[97]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[55] ^ t[33];
  assign t[36] = t[56] & t[57];
  assign t[37] = t[58] ^ t[59];
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[4] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = t[64];
  assign t[42] = ~(t[65]);
  assign t[43] = t[66];
  assign t[44] = t[67] ? t[68] : t[169];
  assign t[45] = t[69] ^ t[24];
  assign t[46] = t[70] & t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[170] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = t[8] ? t[9] : t[164];
  assign t[50] = ~(t[168]);
  assign t[51] = ~(t[76] & t[171]);
  assign t[52] = t[67] ? t[77] : t[172];
  assign t[53] = t[78] ^ t[36];
  assign t[54] = t[79] & t[80];
  assign t[55] = t[67] ? t[81] : t[173];
  assign t[56] = ~(t[82]);
  assign t[57] = t[174] ^ t[83];
  assign t[58] = t[84] ^ t[85];
  assign t[59] = t[86] & t[87];
  assign t[5] = ~(t[10]);
  assign t[60] = t[8] ? t[88] : t[175];
  assign t[61] = t[62] ^ t[89];
  assign t[62] = t[90] ^ t[91];
  assign t[63] = t[92] & t[93];
  assign t[64] = t[67] ? t[94] : t[176];
  assign t[65] = ~t[95];
  assign t[66] = t[67] ? t[96] : t[177];
  assign t[67] = ~(t[15]);
  assign t[68] = t[169] ^ t[97];
  assign t[69] = t[98] & t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[100] ^ t[45]);
  assign t[71] = t[101] ^ t[43];
  assign t[72] = ~(t[74] & t[102]);
  assign t[73] = ~(t[178] ^ t[103]);
  assign t[74] = ~(t[104] & t[105]);
  assign t[75] = ~(t[48]);
  assign t[76] = ~(t[174]);
  assign t[77] = t[172] ^ t[106];
  assign t[78] = t[107] & t[108];
  assign t[79] = ~(t[109] ^ t[53]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[110] ^ t[57];
  assign t[81] = t[173] ^ t[111];
  assign t[82] = t[167] ^ t[112];
  assign t[83] = t[67] ? t[113] : t[179];
  assign t[84] = t[67] ? t[114] : t[180];
  assign t[85] = t[67] ? t[115] : t[181];
  assign t[86] = ~(t[58] ^ t[116]);
  assign t[87] = t[117] ^ t[118];
  assign t[88] = t[175] ^ t[119];
  assign t[89] = t[120] & t[121];
  assign t[8] = ~(t[15]);
  assign t[90] = t[122] & t[123];
  assign t[91] = t[124] & t[125];
  assign t[92] = ~(t[90] ^ t[126]);
  assign t[93] = t[127] ^ t[128];
  assign t[94] = t[176] ^ t[129];
  assign t[95] = t[67] ? t[130] : t[182];
  assign t[96] = t[177] ^ t[131];
  assign t[97] = t[75] ? x[62] : x[61];
  assign t[98] = ~(t[132]);
  assign t[99] = ~(t[41]);
  assign t[9] = t[164] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind44(x, y);
 input [111:0] x;
 output y;

 wire [334:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[129] ^ t[172];
  assign t[101] = ~(t[168]);
  assign t[102] = t[130] & t[129];
  assign t[103] = t[28] ? x[71] : x[70];
  assign t[104] = ~(t[48]);
  assign t[105] = t[104] ? x[73] : x[72];
  assign t[106] = ~(t[131]);
  assign t[107] = ~(t[35]);
  assign t[108] = ~(t[36]);
  assign t[109] = t[53] ? t[132] : t[173];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[169] ^ t[133];
  assign t[111] = t[134] ? x[78] : x[77];
  assign t[112] = t[74] ? x[80] : x[79];
  assign t[113] = ~(t[119]);
  assign t[114] = ~(t[135]);
  assign t[115] = ~(t[59]);
  assign t[116] = t[53] ? t[136] : t[174];
  assign t[117] = t[39] ^ t[135];
  assign t[118] = t[135] ^ t[60];
  assign t[119] = t[116] ^ t[59];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[170] ^ t[137];
  assign t[121] = t[171] ^ t[138];
  assign t[122] = t[139] & t[140];
  assign t[123] = t[141] & t[94];
  assign t[124] = t[142];
  assign t[125] = t[53] ? t[143] : t[175];
  assign t[126] = t[4] ^ t[52];
  assign t[127] = ~(t[130] | t[129]);
  assign t[128] = ~(t[144] | t[101]);
  assign t[129] = ~(t[176]);
  assign t[12] = t[21] ^ t[22];
  assign t[130] = ~(t[172]);
  assign t[131] = t[58] ^ t[36];
  assign t[132] = t[173] ^ t[145];
  assign t[133] = t[104] ? x[91] : x[90];
  assign t[134] = ~(t[48]);
  assign t[135] = t[53] ? t[146] : t[177];
  assign t[136] = t[174] ^ t[147];
  assign t[137] = t[74] ? x[96] : x[95];
  assign t[138] = t[104] ? x[98] : x[97];
  assign t[139] = ~(t[148]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[63]);
  assign t[141] = ~(t[64]);
  assign t[142] = t[53] ? t[149] : t[178];
  assign t[143] = t[175] ^ t[150];
  assign t[144] = ~(t[160]);
  assign t[145] = t[104] ? x[103] : x[102];
  assign t[146] = t[177] ^ t[151];
  assign t[147] = t[134] ? x[105] : x[104];
  assign t[148] = t[94] ^ t[64];
  assign t[149] = t[178] ^ t[152];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[74] ? x[107] : x[106];
  assign t[151] = t[134] ? x[109] : x[108];
  assign t[152] = t[74] ? x[111] : x[110];
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = t[205] ^ x[4];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[9];
  assign t[181] = t[207] ^ x[12];
  assign t[182] = t[208] ^ x[15];
  assign t[183] = t[209] ^ x[18];
  assign t[184] = t[210] ^ x[21];
  assign t[185] = t[211] ^ x[24];
  assign t[186] = t[212] ^ x[27];
  assign t[187] = t[213] ^ x[30];
  assign t[188] = t[214] ^ x[33];
  assign t[189] = t[215] ^ x[36];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[39];
  assign t[191] = t[217] ^ x[42];
  assign t[192] = t[218] ^ x[45];
  assign t[193] = t[219] ^ x[48];
  assign t[194] = t[220] ^ x[53];
  assign t[195] = t[221] ^ x[60];
  assign t[196] = t[222] ^ x[63];
  assign t[197] = t[223] ^ x[66];
  assign t[198] = t[224] ^ x[69];
  assign t[199] = t[225] ^ x[76];
  assign t[19] = t[33] ^ t[25];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[83];
  assign t[201] = t[227] ^ x[86];
  assign t[202] = t[228] ^ x[89];
  assign t[203] = t[229] ^ x[94];
  assign t[204] = t[230] ^ x[101];
  assign t[205] = (t[231] & ~t[232]);
  assign t[206] = (t[233] & ~t[234]);
  assign t[207] = (t[235] & ~t[236]);
  assign t[208] = (t[237] & ~t[238]);
  assign t[209] = (t[239] & ~t[240]);
  assign t[20] = t[34] & t[4];
  assign t[210] = (t[241] & ~t[242]);
  assign t[211] = (t[243] & ~t[244]);
  assign t[212] = (t[245] & ~t[246]);
  assign t[213] = (t[247] & ~t[248]);
  assign t[214] = (t[249] & ~t[250]);
  assign t[215] = (t[251] & ~t[252]);
  assign t[216] = (t[253] & ~t[254]);
  assign t[217] = (t[255] & ~t[256]);
  assign t[218] = (t[257] & ~t[258]);
  assign t[219] = (t[259] & ~t[260]);
  assign t[21] = t[35] ^ t[36];
  assign t[220] = (t[261] & ~t[262]);
  assign t[221] = (t[263] & ~t[264]);
  assign t[222] = (t[265] & ~t[266]);
  assign t[223] = (t[267] & ~t[268]);
  assign t[224] = (t[269] & ~t[270]);
  assign t[225] = (t[271] & ~t[272]);
  assign t[226] = (t[273] & ~t[274]);
  assign t[227] = (t[275] & ~t[276]);
  assign t[228] = (t[277] & ~t[278]);
  assign t[229] = (t[279] & ~t[280]);
  assign t[22] = t[37] & t[38];
  assign t[230] = (t[281] & ~t[282]);
  assign t[231] = t[283] ^ x[4];
  assign t[232] = t[284] ^ x[3];
  assign t[233] = t[285] ^ x[9];
  assign t[234] = t[286] ^ x[8];
  assign t[235] = t[287] ^ x[12];
  assign t[236] = t[288] ^ x[11];
  assign t[237] = t[289] ^ x[15];
  assign t[238] = t[290] ^ x[14];
  assign t[239] = t[291] ^ x[18];
  assign t[23] = t[39] ^ t[40];
  assign t[240] = t[292] ^ x[17];
  assign t[241] = t[293] ^ x[21];
  assign t[242] = t[294] ^ x[20];
  assign t[243] = t[295] ^ x[24];
  assign t[244] = t[296] ^ x[23];
  assign t[245] = t[297] ^ x[27];
  assign t[246] = t[298] ^ x[26];
  assign t[247] = t[299] ^ x[30];
  assign t[248] = t[300] ^ x[29];
  assign t[249] = t[301] ^ x[33];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[302] ^ x[32];
  assign t[251] = t[303] ^ x[36];
  assign t[252] = t[304] ^ x[35];
  assign t[253] = t[305] ^ x[39];
  assign t[254] = t[306] ^ x[38];
  assign t[255] = t[307] ^ x[42];
  assign t[256] = t[308] ^ x[41];
  assign t[257] = t[309] ^ x[45];
  assign t[258] = t[310] ^ x[44];
  assign t[259] = t[311] ^ x[48];
  assign t[25] = t[8] ? t[43] : t[154];
  assign t[260] = t[312] ^ x[47];
  assign t[261] = t[313] ^ x[53];
  assign t[262] = t[314] ^ x[52];
  assign t[263] = t[315] ^ x[60];
  assign t[264] = t[316] ^ x[59];
  assign t[265] = t[317] ^ x[63];
  assign t[266] = t[318] ^ x[62];
  assign t[267] = t[319] ^ x[66];
  assign t[268] = t[320] ^ x[65];
  assign t[269] = t[321] ^ x[69];
  assign t[26] = t[44] ^ t[45];
  assign t[270] = t[322] ^ x[68];
  assign t[271] = t[323] ^ x[76];
  assign t[272] = t[324] ^ x[75];
  assign t[273] = t[325] ^ x[83];
  assign t[274] = t[326] ^ x[82];
  assign t[275] = t[327] ^ x[86];
  assign t[276] = t[328] ^ x[85];
  assign t[277] = t[329] ^ x[89];
  assign t[278] = t[330] ^ x[88];
  assign t[279] = t[331] ^ x[94];
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = t[332] ^ x[93];
  assign t[281] = t[333] ^ x[101];
  assign t[282] = t[334] ^ x[100];
  assign t[283] = (x[2]);
  assign t[284] = (x[2]);
  assign t[285] = (x[7]);
  assign t[286] = (x[7]);
  assign t[287] = (x[10]);
  assign t[288] = (x[10]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[48]);
  assign t[290] = (x[13]);
  assign t[291] = (x[16]);
  assign t[292] = (x[16]);
  assign t[293] = (x[19]);
  assign t[294] = (x[19]);
  assign t[295] = (x[22]);
  assign t[296] = (x[22]);
  assign t[297] = (x[25]);
  assign t[298] = (x[25]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[28]);
  assign t[301] = (x[31]);
  assign t[302] = (x[31]);
  assign t[303] = (x[34]);
  assign t[304] = (x[34]);
  assign t[305] = (x[37]);
  assign t[306] = (x[37]);
  assign t[307] = (x[40]);
  assign t[308] = (x[40]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[156]);
  assign t[310] = (x[43]);
  assign t[311] = (x[46]);
  assign t[312] = (x[46]);
  assign t[313] = (x[51]);
  assign t[314] = (x[51]);
  assign t[315] = (x[58]);
  assign t[316] = (x[58]);
  assign t[317] = (x[61]);
  assign t[318] = (x[61]);
  assign t[319] = (x[64]);
  assign t[31] = ~(t[157]);
  assign t[320] = (x[64]);
  assign t[321] = (x[67]);
  assign t[322] = (x[67]);
  assign t[323] = (x[74]);
  assign t[324] = (x[74]);
  assign t[325] = (x[81]);
  assign t[326] = (x[81]);
  assign t[327] = (x[84]);
  assign t[328] = (x[84]);
  assign t[329] = (x[87]);
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = (x[87]);
  assign t[331] = (x[92]);
  assign t[332] = (x[92]);
  assign t[333] = (x[99]);
  assign t[334] = (x[99]);
  assign t[33] = t[8] ? t[51] : t[158];
  assign t[34] = ~(t[52]);
  assign t[35] = t[53] ? t[54] : t[159];
  assign t[36] = t[157] ^ t[55];
  assign t[37] = ~(t[21] ^ t[56]);
  assign t[38] = t[57] ^ t[58];
  assign t[39] = t[59] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[154] ^ t[67];
  assign t[44] = t[68] ^ t[20];
  assign t[45] = t[69] & t[70];
  assign t[46] = ~(t[71] & t[72]);
  assign t[47] = t[160] | t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = ~(t[161]);
  assign t[4] = t[8] ? t[9] : t[153];
  assign t[50] = ~(t[75] & t[162]);
  assign t[51] = t[158] ^ t[76];
  assign t[52] = t[8] ? t[77] : t[163];
  assign t[53] = ~(t[15]);
  assign t[54] = t[159] ^ t[78];
  assign t[55] = t[53] ? t[79] : t[164];
  assign t[56] = t[80] ^ t[81];
  assign t[57] = t[36] ^ t[82];
  assign t[58] = t[165] ^ t[83];
  assign t[59] = t[53] ? t[84] : t[166];
  assign t[5] = ~(t[10]);
  assign t[60] = t[53] ? t[85] : t[167];
  assign t[61] = t[86] ^ t[87];
  assign t[62] = t[88] & t[89];
  assign t[63] = t[90];
  assign t[64] = ~t[91];
  assign t[65] = ~(t[41] ^ t[92]);
  assign t[66] = t[93] ^ t[94];
  assign t[67] = t[28] ? x[50] : x[49];
  assign t[68] = t[95] & t[96];
  assign t[69] = ~(t[97] ^ t[44]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[98] ^ t[4];
  assign t[71] = ~(t[73] & t[99]);
  assign t[72] = ~(t[168] ^ t[100]);
  assign t[73] = ~(t[101] & t[102]);
  assign t[74] = ~(t[47]);
  assign t[75] = ~(t[165]);
  assign t[76] = t[28] ? x[55] : x[54];
  assign t[77] = t[163] ^ t[103];
  assign t[78] = t[104] ? x[57] : x[56];
  assign t[79] = t[164] ^ t[105];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[106] & t[107];
  assign t[81] = t[108] & t[58];
  assign t[82] = t[161] ^ t[109];
  assign t[83] = t[53] ? t[110] : t[169];
  assign t[84] = t[166] ^ t[111];
  assign t[85] = t[167] ^ t[112];
  assign t[86] = t[113] & t[114];
  assign t[87] = t[115] & t[116];
  assign t[88] = ~(t[86] ^ t[117]);
  assign t[89] = t[118] ^ t[119];
  assign t[8] = ~(t[15]);
  assign t[90] = t[53] ? t[120] : t[170];
  assign t[91] = t[53] ? t[121] : t[171];
  assign t[92] = t[122] ^ t[123];
  assign t[93] = t[64] ^ t[124];
  assign t[94] = t[125];
  assign t[95] = ~(t[126]);
  assign t[96] = ~(t[33]);
  assign t[97] = t[33] ^ t[52];
  assign t[98] = t[52] ^ t[25];
  assign t[99] = ~(t[127] & t[128]);
  assign t[9] = t[153] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [111:0] x;
 output y;

 wire [334:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[129] ^ t[172];
  assign t[101] = ~(t[168]);
  assign t[102] = t[130] & t[129];
  assign t[103] = t[28] ? x[71] : x[70];
  assign t[104] = ~(t[48]);
  assign t[105] = t[104] ? x[73] : x[72];
  assign t[106] = ~(t[131]);
  assign t[107] = ~(t[35]);
  assign t[108] = ~(t[36]);
  assign t[109] = t[53] ? t[132] : t[173];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[169] ^ t[133];
  assign t[111] = t[134] ? x[78] : x[77];
  assign t[112] = t[74] ? x[80] : x[79];
  assign t[113] = ~(t[119]);
  assign t[114] = ~(t[135]);
  assign t[115] = ~(t[59]);
  assign t[116] = t[53] ? t[136] : t[174];
  assign t[117] = t[39] ^ t[135];
  assign t[118] = t[135] ^ t[60];
  assign t[119] = t[116] ^ t[59];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[170] ^ t[137];
  assign t[121] = t[171] ^ t[138];
  assign t[122] = t[139] & t[140];
  assign t[123] = t[141] & t[94];
  assign t[124] = t[142];
  assign t[125] = t[53] ? t[143] : t[175];
  assign t[126] = t[4] ^ t[52];
  assign t[127] = ~(t[130] | t[129]);
  assign t[128] = ~(t[144] | t[101]);
  assign t[129] = ~(t[176]);
  assign t[12] = t[21] ^ t[22];
  assign t[130] = ~(t[172]);
  assign t[131] = t[58] ^ t[36];
  assign t[132] = t[173] ^ t[145];
  assign t[133] = t[104] ? x[91] : x[90];
  assign t[134] = ~(t[48]);
  assign t[135] = t[53] ? t[146] : t[177];
  assign t[136] = t[174] ^ t[147];
  assign t[137] = t[74] ? x[96] : x[95];
  assign t[138] = t[104] ? x[98] : x[97];
  assign t[139] = ~(t[148]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[63]);
  assign t[141] = ~(t[64]);
  assign t[142] = t[53] ? t[149] : t[178];
  assign t[143] = t[175] ^ t[150];
  assign t[144] = ~(t[160]);
  assign t[145] = t[104] ? x[103] : x[102];
  assign t[146] = t[177] ^ t[151];
  assign t[147] = t[134] ? x[105] : x[104];
  assign t[148] = t[94] ^ t[64];
  assign t[149] = t[178] ^ t[152];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[74] ? x[107] : x[106];
  assign t[151] = t[134] ? x[109] : x[108];
  assign t[152] = t[74] ? x[111] : x[110];
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = t[205] ^ x[4];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[9];
  assign t[181] = t[207] ^ x[12];
  assign t[182] = t[208] ^ x[15];
  assign t[183] = t[209] ^ x[18];
  assign t[184] = t[210] ^ x[21];
  assign t[185] = t[211] ^ x[24];
  assign t[186] = t[212] ^ x[27];
  assign t[187] = t[213] ^ x[30];
  assign t[188] = t[214] ^ x[33];
  assign t[189] = t[215] ^ x[36];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[39];
  assign t[191] = t[217] ^ x[42];
  assign t[192] = t[218] ^ x[45];
  assign t[193] = t[219] ^ x[48];
  assign t[194] = t[220] ^ x[53];
  assign t[195] = t[221] ^ x[60];
  assign t[196] = t[222] ^ x[63];
  assign t[197] = t[223] ^ x[66];
  assign t[198] = t[224] ^ x[69];
  assign t[199] = t[225] ^ x[76];
  assign t[19] = t[33] ^ t[25];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[83];
  assign t[201] = t[227] ^ x[86];
  assign t[202] = t[228] ^ x[89];
  assign t[203] = t[229] ^ x[94];
  assign t[204] = t[230] ^ x[101];
  assign t[205] = (t[231] & ~t[232]);
  assign t[206] = (t[233] & ~t[234]);
  assign t[207] = (t[235] & ~t[236]);
  assign t[208] = (t[237] & ~t[238]);
  assign t[209] = (t[239] & ~t[240]);
  assign t[20] = t[34] & t[4];
  assign t[210] = (t[241] & ~t[242]);
  assign t[211] = (t[243] & ~t[244]);
  assign t[212] = (t[245] & ~t[246]);
  assign t[213] = (t[247] & ~t[248]);
  assign t[214] = (t[249] & ~t[250]);
  assign t[215] = (t[251] & ~t[252]);
  assign t[216] = (t[253] & ~t[254]);
  assign t[217] = (t[255] & ~t[256]);
  assign t[218] = (t[257] & ~t[258]);
  assign t[219] = (t[259] & ~t[260]);
  assign t[21] = t[35] ^ t[36];
  assign t[220] = (t[261] & ~t[262]);
  assign t[221] = (t[263] & ~t[264]);
  assign t[222] = (t[265] & ~t[266]);
  assign t[223] = (t[267] & ~t[268]);
  assign t[224] = (t[269] & ~t[270]);
  assign t[225] = (t[271] & ~t[272]);
  assign t[226] = (t[273] & ~t[274]);
  assign t[227] = (t[275] & ~t[276]);
  assign t[228] = (t[277] & ~t[278]);
  assign t[229] = (t[279] & ~t[280]);
  assign t[22] = t[37] & t[38];
  assign t[230] = (t[281] & ~t[282]);
  assign t[231] = t[283] ^ x[4];
  assign t[232] = t[284] ^ x[3];
  assign t[233] = t[285] ^ x[9];
  assign t[234] = t[286] ^ x[8];
  assign t[235] = t[287] ^ x[12];
  assign t[236] = t[288] ^ x[11];
  assign t[237] = t[289] ^ x[15];
  assign t[238] = t[290] ^ x[14];
  assign t[239] = t[291] ^ x[18];
  assign t[23] = t[39] ^ t[40];
  assign t[240] = t[292] ^ x[17];
  assign t[241] = t[293] ^ x[21];
  assign t[242] = t[294] ^ x[20];
  assign t[243] = t[295] ^ x[24];
  assign t[244] = t[296] ^ x[23];
  assign t[245] = t[297] ^ x[27];
  assign t[246] = t[298] ^ x[26];
  assign t[247] = t[299] ^ x[30];
  assign t[248] = t[300] ^ x[29];
  assign t[249] = t[301] ^ x[33];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[302] ^ x[32];
  assign t[251] = t[303] ^ x[36];
  assign t[252] = t[304] ^ x[35];
  assign t[253] = t[305] ^ x[39];
  assign t[254] = t[306] ^ x[38];
  assign t[255] = t[307] ^ x[42];
  assign t[256] = t[308] ^ x[41];
  assign t[257] = t[309] ^ x[45];
  assign t[258] = t[310] ^ x[44];
  assign t[259] = t[311] ^ x[48];
  assign t[25] = t[8] ? t[43] : t[154];
  assign t[260] = t[312] ^ x[47];
  assign t[261] = t[313] ^ x[53];
  assign t[262] = t[314] ^ x[52];
  assign t[263] = t[315] ^ x[60];
  assign t[264] = t[316] ^ x[59];
  assign t[265] = t[317] ^ x[63];
  assign t[266] = t[318] ^ x[62];
  assign t[267] = t[319] ^ x[66];
  assign t[268] = t[320] ^ x[65];
  assign t[269] = t[321] ^ x[69];
  assign t[26] = t[44] ^ t[45];
  assign t[270] = t[322] ^ x[68];
  assign t[271] = t[323] ^ x[76];
  assign t[272] = t[324] ^ x[75];
  assign t[273] = t[325] ^ x[83];
  assign t[274] = t[326] ^ x[82];
  assign t[275] = t[327] ^ x[86];
  assign t[276] = t[328] ^ x[85];
  assign t[277] = t[329] ^ x[89];
  assign t[278] = t[330] ^ x[88];
  assign t[279] = t[331] ^ x[94];
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = t[332] ^ x[93];
  assign t[281] = t[333] ^ x[101];
  assign t[282] = t[334] ^ x[100];
  assign t[283] = (x[2]);
  assign t[284] = (x[2]);
  assign t[285] = (x[7]);
  assign t[286] = (x[7]);
  assign t[287] = (x[10]);
  assign t[288] = (x[10]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[48]);
  assign t[290] = (x[13]);
  assign t[291] = (x[16]);
  assign t[292] = (x[16]);
  assign t[293] = (x[19]);
  assign t[294] = (x[19]);
  assign t[295] = (x[22]);
  assign t[296] = (x[22]);
  assign t[297] = (x[25]);
  assign t[298] = (x[25]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[28]);
  assign t[301] = (x[31]);
  assign t[302] = (x[31]);
  assign t[303] = (x[34]);
  assign t[304] = (x[34]);
  assign t[305] = (x[37]);
  assign t[306] = (x[37]);
  assign t[307] = (x[40]);
  assign t[308] = (x[40]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[156]);
  assign t[310] = (x[43]);
  assign t[311] = (x[46]);
  assign t[312] = (x[46]);
  assign t[313] = (x[51]);
  assign t[314] = (x[51]);
  assign t[315] = (x[58]);
  assign t[316] = (x[58]);
  assign t[317] = (x[61]);
  assign t[318] = (x[61]);
  assign t[319] = (x[64]);
  assign t[31] = ~(t[157]);
  assign t[320] = (x[64]);
  assign t[321] = (x[67]);
  assign t[322] = (x[67]);
  assign t[323] = (x[74]);
  assign t[324] = (x[74]);
  assign t[325] = (x[81]);
  assign t[326] = (x[81]);
  assign t[327] = (x[84]);
  assign t[328] = (x[84]);
  assign t[329] = (x[87]);
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = (x[87]);
  assign t[331] = (x[92]);
  assign t[332] = (x[92]);
  assign t[333] = (x[99]);
  assign t[334] = (x[99]);
  assign t[33] = t[8] ? t[51] : t[158];
  assign t[34] = ~(t[52]);
  assign t[35] = t[53] ? t[54] : t[159];
  assign t[36] = t[157] ^ t[55];
  assign t[37] = ~(t[21] ^ t[56]);
  assign t[38] = t[57] ^ t[58];
  assign t[39] = t[59] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[154] ^ t[67];
  assign t[44] = t[68] ^ t[20];
  assign t[45] = t[69] & t[70];
  assign t[46] = ~(t[71] & t[72]);
  assign t[47] = t[160] | t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = ~(t[161]);
  assign t[4] = t[8] ? t[9] : t[153];
  assign t[50] = ~(t[75] & t[162]);
  assign t[51] = t[158] ^ t[76];
  assign t[52] = t[8] ? t[77] : t[163];
  assign t[53] = ~(t[15]);
  assign t[54] = t[159] ^ t[78];
  assign t[55] = t[53] ? t[79] : t[164];
  assign t[56] = t[80] ^ t[81];
  assign t[57] = t[36] ^ t[82];
  assign t[58] = t[165] ^ t[83];
  assign t[59] = t[53] ? t[84] : t[166];
  assign t[5] = ~(t[10]);
  assign t[60] = t[53] ? t[85] : t[167];
  assign t[61] = t[86] ^ t[87];
  assign t[62] = t[88] & t[89];
  assign t[63] = t[90];
  assign t[64] = ~t[91];
  assign t[65] = ~(t[41] ^ t[92]);
  assign t[66] = t[93] ^ t[94];
  assign t[67] = t[28] ? x[50] : x[49];
  assign t[68] = t[95] & t[96];
  assign t[69] = ~(t[97] ^ t[44]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[98] ^ t[4];
  assign t[71] = ~(t[73] & t[99]);
  assign t[72] = ~(t[168] ^ t[100]);
  assign t[73] = ~(t[101] & t[102]);
  assign t[74] = ~(t[47]);
  assign t[75] = ~(t[165]);
  assign t[76] = t[28] ? x[55] : x[54];
  assign t[77] = t[163] ^ t[103];
  assign t[78] = t[104] ? x[57] : x[56];
  assign t[79] = t[164] ^ t[105];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[106] & t[107];
  assign t[81] = t[108] & t[58];
  assign t[82] = t[161] ^ t[109];
  assign t[83] = t[53] ? t[110] : t[169];
  assign t[84] = t[166] ^ t[111];
  assign t[85] = t[167] ^ t[112];
  assign t[86] = t[113] & t[114];
  assign t[87] = t[115] & t[116];
  assign t[88] = ~(t[86] ^ t[117]);
  assign t[89] = t[118] ^ t[119];
  assign t[8] = ~(t[15]);
  assign t[90] = t[53] ? t[120] : t[170];
  assign t[91] = t[53] ? t[121] : t[171];
  assign t[92] = t[122] ^ t[123];
  assign t[93] = t[64] ^ t[124];
  assign t[94] = t[125];
  assign t[95] = ~(t[126]);
  assign t[96] = ~(t[33]);
  assign t[97] = t[33] ^ t[52];
  assign t[98] = t[52] ^ t[25];
  assign t[99] = ~(t[127] & t[128]);
  assign t[9] = t[153] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind46(x, y);
 input [111:0] x;
 output y;

 wire [333:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[127] & t[126];
  assign t[101] = t[166] ^ t[128];
  assign t[102] = t[167] ^ t[129];
  assign t[103] = ~(t[109]);
  assign t[104] = ~(t[130]);
  assign t[105] = ~(t[51]);
  assign t[106] = t[131];
  assign t[107] = t[33] ^ t[130];
  assign t[108] = t[130] ^ t[52];
  assign t[109] = t[106] ^ t[51];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[132]);
  assign t[111] = ~(t[133]);
  assign t[112] = ~(t[134]);
  assign t[113] = t[55] ? t[135] : t[172];
  assign t[114] = t[133] ^ t[134];
  assign t[115] = t[134] ^ t[35];
  assign t[116] = ~(t[136]);
  assign t[117] = ~(t[4]);
  assign t[118] = ~(t[37]);
  assign t[119] = t[168] ^ t[137];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[28] ? x[76] : x[75];
  assign t[121] = ~(t[48]);
  assign t[122] = t[169] ^ t[138];
  assign t[123] = t[170] ^ t[139];
  assign t[124] = ~(t[127] | t[126]);
  assign t[125] = ~(t[140] | t[99]);
  assign t[126] = ~(t[173]);
  assign t[127] = ~(t[171]);
  assign t[128] = t[121] ? x[81] : x[80];
  assign t[129] = t[75] ? x[83] : x[82];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[141];
  assign t[131] = t[55] ? t[142] : t[174];
  assign t[132] = t[113] ^ t[134];
  assign t[133] = t[55] ? t[143] : t[175];
  assign t[134] = t[55] ? t[144] : t[176];
  assign t[135] = t[172] ^ t[145];
  assign t[136] = t[62] ^ t[37];
  assign t[137] = t[28] ? x[94] : x[93];
  assign t[138] = t[121] ? x[96] : x[95];
  assign t[139] = t[121] ? x[98] : x[97];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[161]);
  assign t[141] = t[55] ? t[146] : t[177];
  assign t[142] = t[174] ^ t[147];
  assign t[143] = t[175] ^ t[148];
  assign t[144] = t[176] ^ t[149];
  assign t[145] = t[150] ? x[103] : x[102];
  assign t[146] = t[177] ^ t[151];
  assign t[147] = t[75] ? x[105] : x[104];
  assign t[148] = t[150] ? x[107] : x[106];
  assign t[149] = t[150] ? x[109] : x[108];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = ~(t[48]);
  assign t[151] = t[75] ? x[111] : x[110];
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = t[204] ^ x[4];
  assign t[179] = t[205] ^ x[9];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[12];
  assign t[181] = t[207] ^ x[15];
  assign t[182] = t[208] ^ x[18];
  assign t[183] = t[209] ^ x[21];
  assign t[184] = t[210] ^ x[24];
  assign t[185] = t[211] ^ x[27];
  assign t[186] = t[212] ^ x[30];
  assign t[187] = t[213] ^ x[33];
  assign t[188] = t[214] ^ x[36];
  assign t[189] = t[215] ^ x[39];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[42];
  assign t[191] = t[217] ^ x[45];
  assign t[192] = t[218] ^ x[48];
  assign t[193] = t[219] ^ x[51];
  assign t[194] = t[220] ^ x[58];
  assign t[195] = t[221] ^ x[65];
  assign t[196] = t[222] ^ x[68];
  assign t[197] = t[223] ^ x[71];
  assign t[198] = t[224] ^ x[74];
  assign t[199] = t[225] ^ x[79];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[86];
  assign t[201] = t[227] ^ x[89];
  assign t[202] = t[228] ^ x[92];
  assign t[203] = t[229] ^ x[101];
  assign t[204] = (t[230] & ~t[231]);
  assign t[205] = (t[232] & ~t[233]);
  assign t[206] = (t[234] & ~t[235]);
  assign t[207] = (t[236] & ~t[237]);
  assign t[208] = (t[238] & ~t[239]);
  assign t[209] = (t[240] & ~t[241]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[242] & ~t[243]);
  assign t[211] = (t[244] & ~t[245]);
  assign t[212] = (t[246] & ~t[247]);
  assign t[213] = (t[248] & ~t[249]);
  assign t[214] = (t[250] & ~t[251]);
  assign t[215] = (t[252] & ~t[253]);
  assign t[216] = (t[254] & ~t[255]);
  assign t[217] = (t[256] & ~t[257]);
  assign t[218] = (t[258] & ~t[259]);
  assign t[219] = (t[260] & ~t[261]);
  assign t[21] = t[4] ^ t[37];
  assign t[220] = (t[262] & ~t[263]);
  assign t[221] = (t[264] & ~t[265]);
  assign t[222] = (t[266] & ~t[267]);
  assign t[223] = (t[268] & ~t[269]);
  assign t[224] = (t[270] & ~t[271]);
  assign t[225] = (t[272] & ~t[273]);
  assign t[226] = (t[274] & ~t[275]);
  assign t[227] = (t[276] & ~t[277]);
  assign t[228] = (t[278] & ~t[279]);
  assign t[229] = (t[280] & ~t[281]);
  assign t[22] = t[38] & t[39];
  assign t[230] = t[282] ^ x[4];
  assign t[231] = t[283] ^ x[3];
  assign t[232] = t[284] ^ x[9];
  assign t[233] = t[285] ^ x[8];
  assign t[234] = t[286] ^ x[12];
  assign t[235] = t[287] ^ x[11];
  assign t[236] = t[288] ^ x[15];
  assign t[237] = t[289] ^ x[14];
  assign t[238] = t[290] ^ x[18];
  assign t[239] = t[291] ^ x[17];
  assign t[23] = t[153] ^ t[40];
  assign t[240] = t[292] ^ x[21];
  assign t[241] = t[293] ^ x[20];
  assign t[242] = t[294] ^ x[24];
  assign t[243] = t[295] ^ x[23];
  assign t[244] = t[296] ^ x[27];
  assign t[245] = t[297] ^ x[26];
  assign t[246] = t[298] ^ x[30];
  assign t[247] = t[299] ^ x[29];
  assign t[248] = t[300] ^ x[33];
  assign t[249] = t[301] ^ x[32];
  assign t[24] = t[154] ^ t[41];
  assign t[250] = t[302] ^ x[36];
  assign t[251] = t[303] ^ x[35];
  assign t[252] = t[304] ^ x[39];
  assign t[253] = t[305] ^ x[38];
  assign t[254] = t[306] ^ x[42];
  assign t[255] = t[307] ^ x[41];
  assign t[256] = t[308] ^ x[45];
  assign t[257] = t[309] ^ x[44];
  assign t[258] = t[310] ^ x[48];
  assign t[259] = t[311] ^ x[47];
  assign t[25] = t[42] ^ t[43];
  assign t[260] = t[312] ^ x[51];
  assign t[261] = t[313] ^ x[50];
  assign t[262] = t[314] ^ x[58];
  assign t[263] = t[315] ^ x[57];
  assign t[264] = t[316] ^ x[65];
  assign t[265] = t[317] ^ x[64];
  assign t[266] = t[318] ^ x[68];
  assign t[267] = t[319] ^ x[67];
  assign t[268] = t[320] ^ x[71];
  assign t[269] = t[321] ^ x[70];
  assign t[26] = t[44] & t[45];
  assign t[270] = t[322] ^ x[74];
  assign t[271] = t[323] ^ x[73];
  assign t[272] = t[324] ^ x[79];
  assign t[273] = t[325] ^ x[78];
  assign t[274] = t[326] ^ x[86];
  assign t[275] = t[327] ^ x[85];
  assign t[276] = t[328] ^ x[89];
  assign t[277] = t[329] ^ x[88];
  assign t[278] = t[330] ^ x[92];
  assign t[279] = t[331] ^ x[91];
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = t[332] ^ x[101];
  assign t[281] = t[333] ^ x[100];
  assign t[282] = (x[2]);
  assign t[283] = (x[2]);
  assign t[284] = (x[7]);
  assign t[285] = (x[7]);
  assign t[286] = (x[10]);
  assign t[287] = (x[10]);
  assign t[288] = (x[13]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[48]);
  assign t[290] = (x[16]);
  assign t[291] = (x[16]);
  assign t[292] = (x[19]);
  assign t[293] = (x[19]);
  assign t[294] = (x[22]);
  assign t[295] = (x[22]);
  assign t[296] = (x[25]);
  assign t[297] = (x[25]);
  assign t[298] = (x[28]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[31]);
  assign t[301] = (x[31]);
  assign t[302] = (x[34]);
  assign t[303] = (x[34]);
  assign t[304] = (x[37]);
  assign t[305] = (x[37]);
  assign t[306] = (x[40]);
  assign t[307] = (x[40]);
  assign t[308] = (x[43]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[156]);
  assign t[310] = (x[46]);
  assign t[311] = (x[46]);
  assign t[312] = (x[49]);
  assign t[313] = (x[49]);
  assign t[314] = (x[56]);
  assign t[315] = (x[56]);
  assign t[316] = (x[63]);
  assign t[317] = (x[63]);
  assign t[318] = (x[66]);
  assign t[319] = (x[66]);
  assign t[31] = ~(t[153]);
  assign t[320] = (x[69]);
  assign t[321] = (x[69]);
  assign t[322] = (x[72]);
  assign t[323] = (x[72]);
  assign t[324] = (x[77]);
  assign t[325] = (x[77]);
  assign t[326] = (x[84]);
  assign t[327] = (x[84]);
  assign t[328] = (x[87]);
  assign t[329] = (x[87]);
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = (x[90]);
  assign t[331] = (x[90]);
  assign t[332] = (x[99]);
  assign t[333] = (x[99]);
  assign t[33] = t[51] ^ t[52];
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[55] ? t[56] : t[157];
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[8] ? t[59] : t[158];
  assign t[38] = ~(t[21] ^ t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[55] ? t[63] : t[159];
  assign t[41] = t[55] ? t[64] : t[160];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[67] & t[68];
  assign t[44] = ~(t[42] ^ t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[161] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[154]);
  assign t[4] = t[8] ? t[9] : t[152];
  assign t[50] = ~(t[76] & t[162]);
  assign t[51] = ~t[77];
  assign t[52] = t[78];
  assign t[53] = t[79] ^ t[80];
  assign t[54] = t[81] & t[82];
  assign t[55] = ~(t[15]);
  assign t[56] = t[157] ^ t[83];
  assign t[57] = t[84] ^ t[85];
  assign t[58] = t[86] & t[87];
  assign t[59] = t[158] ^ t[88];
  assign t[5] = ~(t[10]);
  assign t[60] = t[89] ^ t[90];
  assign t[61] = t[37] ^ t[91];
  assign t[62] = t[8] ? t[92] : t[163];
  assign t[63] = t[159] ^ t[93];
  assign t[64] = t[160] ^ t[94];
  assign t[65] = ~(t[71]);
  assign t[66] = ~(t[95]);
  assign t[67] = ~(t[23]);
  assign t[68] = t[164] ^ t[96];
  assign t[69] = t[13] ^ t[95];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[95] ^ t[24];
  assign t[71] = t[68] ^ t[23];
  assign t[72] = ~(t[74] & t[97]);
  assign t[73] = ~(t[165] ^ t[98]);
  assign t[74] = ~(t[99] & t[100]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[164]);
  assign t[77] = t[55] ? t[101] : t[166];
  assign t[78] = t[55] ? t[102] : t[167];
  assign t[79] = t[103] & t[104];
  assign t[7] = t[13] ^ t[14];
  assign t[80] = t[105] & t[106];
  assign t[81] = ~(t[79] ^ t[107]);
  assign t[82] = t[108] ^ t[109];
  assign t[83] = t[75] ? x[53] : x[52];
  assign t[84] = t[110] & t[111];
  assign t[85] = t[112] & t[113];
  assign t[86] = ~(t[114] ^ t[57]);
  assign t[87] = t[115] ^ t[113];
  assign t[88] = t[28] ? x[55] : x[54];
  assign t[89] = t[116] & t[117];
  assign t[8] = ~(t[15]);
  assign t[90] = t[118] & t[62];
  assign t[91] = t[8] ? t[119] : t[168];
  assign t[92] = t[163] ^ t[120];
  assign t[93] = t[121] ? x[60] : x[59];
  assign t[94] = t[121] ? x[62] : x[61];
  assign t[95] = t[55] ? t[122] : t[169];
  assign t[96] = t[55] ? t[123] : t[170];
  assign t[97] = ~(t[124] & t[125]);
  assign t[98] = t[126] ^ t[171];
  assign t[99] = ~(t[165]);
  assign t[9] = t[152] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind47(x, y);
 input [111:0] x;
 output y;

 wire [333:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[127] & t[126];
  assign t[101] = t[166] ^ t[128];
  assign t[102] = t[167] ^ t[129];
  assign t[103] = ~(t[109]);
  assign t[104] = ~(t[130]);
  assign t[105] = ~(t[51]);
  assign t[106] = t[131];
  assign t[107] = t[33] ^ t[130];
  assign t[108] = t[130] ^ t[52];
  assign t[109] = t[106] ^ t[51];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[132]);
  assign t[111] = ~(t[133]);
  assign t[112] = ~(t[134]);
  assign t[113] = t[55] ? t[135] : t[172];
  assign t[114] = t[133] ^ t[134];
  assign t[115] = t[134] ^ t[35];
  assign t[116] = ~(t[136]);
  assign t[117] = ~(t[4]);
  assign t[118] = ~(t[37]);
  assign t[119] = t[168] ^ t[137];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[28] ? x[76] : x[75];
  assign t[121] = ~(t[48]);
  assign t[122] = t[169] ^ t[138];
  assign t[123] = t[170] ^ t[139];
  assign t[124] = ~(t[127] | t[126]);
  assign t[125] = ~(t[140] | t[99]);
  assign t[126] = ~(t[173]);
  assign t[127] = ~(t[171]);
  assign t[128] = t[121] ? x[81] : x[80];
  assign t[129] = t[75] ? x[83] : x[82];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[141];
  assign t[131] = t[55] ? t[142] : t[174];
  assign t[132] = t[113] ^ t[134];
  assign t[133] = t[55] ? t[143] : t[175];
  assign t[134] = t[55] ? t[144] : t[176];
  assign t[135] = t[172] ^ t[145];
  assign t[136] = t[62] ^ t[37];
  assign t[137] = t[28] ? x[94] : x[93];
  assign t[138] = t[121] ? x[96] : x[95];
  assign t[139] = t[121] ? x[98] : x[97];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[161]);
  assign t[141] = t[55] ? t[146] : t[177];
  assign t[142] = t[174] ^ t[147];
  assign t[143] = t[175] ^ t[148];
  assign t[144] = t[176] ^ t[149];
  assign t[145] = t[150] ? x[103] : x[102];
  assign t[146] = t[177] ^ t[151];
  assign t[147] = t[75] ? x[105] : x[104];
  assign t[148] = t[150] ? x[107] : x[106];
  assign t[149] = t[150] ? x[109] : x[108];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = ~(t[48]);
  assign t[151] = t[75] ? x[111] : x[110];
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = t[204] ^ x[4];
  assign t[179] = t[205] ^ x[9];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[12];
  assign t[181] = t[207] ^ x[15];
  assign t[182] = t[208] ^ x[18];
  assign t[183] = t[209] ^ x[21];
  assign t[184] = t[210] ^ x[24];
  assign t[185] = t[211] ^ x[27];
  assign t[186] = t[212] ^ x[30];
  assign t[187] = t[213] ^ x[33];
  assign t[188] = t[214] ^ x[36];
  assign t[189] = t[215] ^ x[39];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[42];
  assign t[191] = t[217] ^ x[45];
  assign t[192] = t[218] ^ x[48];
  assign t[193] = t[219] ^ x[51];
  assign t[194] = t[220] ^ x[58];
  assign t[195] = t[221] ^ x[65];
  assign t[196] = t[222] ^ x[68];
  assign t[197] = t[223] ^ x[71];
  assign t[198] = t[224] ^ x[74];
  assign t[199] = t[225] ^ x[79];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[86];
  assign t[201] = t[227] ^ x[89];
  assign t[202] = t[228] ^ x[92];
  assign t[203] = t[229] ^ x[101];
  assign t[204] = (t[230] & ~t[231]);
  assign t[205] = (t[232] & ~t[233]);
  assign t[206] = (t[234] & ~t[235]);
  assign t[207] = (t[236] & ~t[237]);
  assign t[208] = (t[238] & ~t[239]);
  assign t[209] = (t[240] & ~t[241]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[242] & ~t[243]);
  assign t[211] = (t[244] & ~t[245]);
  assign t[212] = (t[246] & ~t[247]);
  assign t[213] = (t[248] & ~t[249]);
  assign t[214] = (t[250] & ~t[251]);
  assign t[215] = (t[252] & ~t[253]);
  assign t[216] = (t[254] & ~t[255]);
  assign t[217] = (t[256] & ~t[257]);
  assign t[218] = (t[258] & ~t[259]);
  assign t[219] = (t[260] & ~t[261]);
  assign t[21] = t[4] ^ t[37];
  assign t[220] = (t[262] & ~t[263]);
  assign t[221] = (t[264] & ~t[265]);
  assign t[222] = (t[266] & ~t[267]);
  assign t[223] = (t[268] & ~t[269]);
  assign t[224] = (t[270] & ~t[271]);
  assign t[225] = (t[272] & ~t[273]);
  assign t[226] = (t[274] & ~t[275]);
  assign t[227] = (t[276] & ~t[277]);
  assign t[228] = (t[278] & ~t[279]);
  assign t[229] = (t[280] & ~t[281]);
  assign t[22] = t[38] & t[39];
  assign t[230] = t[282] ^ x[4];
  assign t[231] = t[283] ^ x[3];
  assign t[232] = t[284] ^ x[9];
  assign t[233] = t[285] ^ x[8];
  assign t[234] = t[286] ^ x[12];
  assign t[235] = t[287] ^ x[11];
  assign t[236] = t[288] ^ x[15];
  assign t[237] = t[289] ^ x[14];
  assign t[238] = t[290] ^ x[18];
  assign t[239] = t[291] ^ x[17];
  assign t[23] = t[153] ^ t[40];
  assign t[240] = t[292] ^ x[21];
  assign t[241] = t[293] ^ x[20];
  assign t[242] = t[294] ^ x[24];
  assign t[243] = t[295] ^ x[23];
  assign t[244] = t[296] ^ x[27];
  assign t[245] = t[297] ^ x[26];
  assign t[246] = t[298] ^ x[30];
  assign t[247] = t[299] ^ x[29];
  assign t[248] = t[300] ^ x[33];
  assign t[249] = t[301] ^ x[32];
  assign t[24] = t[154] ^ t[41];
  assign t[250] = t[302] ^ x[36];
  assign t[251] = t[303] ^ x[35];
  assign t[252] = t[304] ^ x[39];
  assign t[253] = t[305] ^ x[38];
  assign t[254] = t[306] ^ x[42];
  assign t[255] = t[307] ^ x[41];
  assign t[256] = t[308] ^ x[45];
  assign t[257] = t[309] ^ x[44];
  assign t[258] = t[310] ^ x[48];
  assign t[259] = t[311] ^ x[47];
  assign t[25] = t[42] ^ t[43];
  assign t[260] = t[312] ^ x[51];
  assign t[261] = t[313] ^ x[50];
  assign t[262] = t[314] ^ x[58];
  assign t[263] = t[315] ^ x[57];
  assign t[264] = t[316] ^ x[65];
  assign t[265] = t[317] ^ x[64];
  assign t[266] = t[318] ^ x[68];
  assign t[267] = t[319] ^ x[67];
  assign t[268] = t[320] ^ x[71];
  assign t[269] = t[321] ^ x[70];
  assign t[26] = t[44] & t[45];
  assign t[270] = t[322] ^ x[74];
  assign t[271] = t[323] ^ x[73];
  assign t[272] = t[324] ^ x[79];
  assign t[273] = t[325] ^ x[78];
  assign t[274] = t[326] ^ x[86];
  assign t[275] = t[327] ^ x[85];
  assign t[276] = t[328] ^ x[89];
  assign t[277] = t[329] ^ x[88];
  assign t[278] = t[330] ^ x[92];
  assign t[279] = t[331] ^ x[91];
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = t[332] ^ x[101];
  assign t[281] = t[333] ^ x[100];
  assign t[282] = (x[2]);
  assign t[283] = (x[2]);
  assign t[284] = (x[7]);
  assign t[285] = (x[7]);
  assign t[286] = (x[10]);
  assign t[287] = (x[10]);
  assign t[288] = (x[13]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[48]);
  assign t[290] = (x[16]);
  assign t[291] = (x[16]);
  assign t[292] = (x[19]);
  assign t[293] = (x[19]);
  assign t[294] = (x[22]);
  assign t[295] = (x[22]);
  assign t[296] = (x[25]);
  assign t[297] = (x[25]);
  assign t[298] = (x[28]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[31]);
  assign t[301] = (x[31]);
  assign t[302] = (x[34]);
  assign t[303] = (x[34]);
  assign t[304] = (x[37]);
  assign t[305] = (x[37]);
  assign t[306] = (x[40]);
  assign t[307] = (x[40]);
  assign t[308] = (x[43]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[156]);
  assign t[310] = (x[46]);
  assign t[311] = (x[46]);
  assign t[312] = (x[49]);
  assign t[313] = (x[49]);
  assign t[314] = (x[56]);
  assign t[315] = (x[56]);
  assign t[316] = (x[63]);
  assign t[317] = (x[63]);
  assign t[318] = (x[66]);
  assign t[319] = (x[66]);
  assign t[31] = ~(t[153]);
  assign t[320] = (x[69]);
  assign t[321] = (x[69]);
  assign t[322] = (x[72]);
  assign t[323] = (x[72]);
  assign t[324] = (x[77]);
  assign t[325] = (x[77]);
  assign t[326] = (x[84]);
  assign t[327] = (x[84]);
  assign t[328] = (x[87]);
  assign t[329] = (x[87]);
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = (x[90]);
  assign t[331] = (x[90]);
  assign t[332] = (x[99]);
  assign t[333] = (x[99]);
  assign t[33] = t[51] ^ t[52];
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[55] ? t[56] : t[157];
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[8] ? t[59] : t[158];
  assign t[38] = ~(t[21] ^ t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[55] ? t[63] : t[159];
  assign t[41] = t[55] ? t[64] : t[160];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[67] & t[68];
  assign t[44] = ~(t[42] ^ t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[161] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[154]);
  assign t[4] = t[8] ? t[9] : t[152];
  assign t[50] = ~(t[76] & t[162]);
  assign t[51] = ~t[77];
  assign t[52] = t[78];
  assign t[53] = t[79] ^ t[80];
  assign t[54] = t[81] & t[82];
  assign t[55] = ~(t[15]);
  assign t[56] = t[157] ^ t[83];
  assign t[57] = t[84] ^ t[85];
  assign t[58] = t[86] & t[87];
  assign t[59] = t[158] ^ t[88];
  assign t[5] = ~(t[10]);
  assign t[60] = t[89] ^ t[90];
  assign t[61] = t[37] ^ t[91];
  assign t[62] = t[8] ? t[92] : t[163];
  assign t[63] = t[159] ^ t[93];
  assign t[64] = t[160] ^ t[94];
  assign t[65] = ~(t[71]);
  assign t[66] = ~(t[95]);
  assign t[67] = ~(t[23]);
  assign t[68] = t[164] ^ t[96];
  assign t[69] = t[13] ^ t[95];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[95] ^ t[24];
  assign t[71] = t[68] ^ t[23];
  assign t[72] = ~(t[74] & t[97]);
  assign t[73] = ~(t[165] ^ t[98]);
  assign t[74] = ~(t[99] & t[100]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[164]);
  assign t[77] = t[55] ? t[101] : t[166];
  assign t[78] = t[55] ? t[102] : t[167];
  assign t[79] = t[103] & t[104];
  assign t[7] = t[13] ^ t[14];
  assign t[80] = t[105] & t[106];
  assign t[81] = ~(t[79] ^ t[107]);
  assign t[82] = t[108] ^ t[109];
  assign t[83] = t[75] ? x[53] : x[52];
  assign t[84] = t[110] & t[111];
  assign t[85] = t[112] & t[113];
  assign t[86] = ~(t[114] ^ t[57]);
  assign t[87] = t[115] ^ t[113];
  assign t[88] = t[28] ? x[55] : x[54];
  assign t[89] = t[116] & t[117];
  assign t[8] = ~(t[15]);
  assign t[90] = t[118] & t[62];
  assign t[91] = t[8] ? t[119] : t[168];
  assign t[92] = t[163] ^ t[120];
  assign t[93] = t[121] ? x[60] : x[59];
  assign t[94] = t[121] ? x[62] : x[61];
  assign t[95] = t[55] ? t[122] : t[169];
  assign t[96] = t[55] ? t[123] : t[170];
  assign t[97] = ~(t[124] & t[125]);
  assign t[98] = t[126] ^ t[171];
  assign t[99] = ~(t[165]);
  assign t[9] = t[152] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind48(x, y);
 input [111:0] x;
 output y;

 wire [323:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[117] ^ t[118];
  assign t[101] = t[118] ^ t[25];
  assign t[102] = ~(t[120] & t[121]);
  assign t[103] = t[122] ^ t[160];
  assign t[104] = ~(t[155]);
  assign t[105] = t[123] & t[122];
  assign t[106] = t[8] ? t[124] : t[161];
  assign t[107] = t[157] ^ t[125];
  assign t[108] = t[74] ? x[71] : x[70];
  assign t[109] = t[74] ? x[73] : x[72];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[158] ^ t[126];
  assign t[111] = t[88] ? x[75] : x[74];
  assign t[112] = t[92] ^ t[114];
  assign t[113] = t[40] ? t[127] : t[162];
  assign t[114] = t[40] ? t[128] : t[163];
  assign t[115] = t[159] ^ t[129];
  assign t[116] = t[99] ^ t[118];
  assign t[117] = t[40] ? t[130] : t[164];
  assign t[118] = t[145] ^ t[131];
  assign t[119] = t[40] ? t[132] : t[165];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[123] | t[122]);
  assign t[121] = ~(t[133] | t[104]);
  assign t[122] = ~(t[166]);
  assign t[123] = ~(t[160]);
  assign t[124] = t[161] ^ t[134];
  assign t[125] = t[28] ? x[92] : x[91];
  assign t[126] = t[135] ? x[94] : x[93];
  assign t[127] = t[162] ^ t[136];
  assign t[128] = t[163] ^ t[137];
  assign t[129] = t[88] ? x[96] : x[95];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[164] ^ t[138];
  assign t[131] = t[27] ? t[139] : t[167];
  assign t[132] = t[165] ^ t[140];
  assign t[133] = ~(t[150]);
  assign t[134] = t[28] ? x[101] : x[100];
  assign t[135] = ~(t[49]);
  assign t[136] = t[88] ? x[103] : x[102];
  assign t[137] = t[88] ? x[105] : x[104];
  assign t[138] = t[74] ? x[107] : x[106];
  assign t[139] = t[167] ^ t[141];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[135] ? x[109] : x[108];
  assign t[141] = t[135] ? x[111] : x[110];
  assign t[142] = (t[168]);
  assign t[143] = (t[169]);
  assign t[144] = (t[170]);
  assign t[145] = (t[171]);
  assign t[146] = (t[172]);
  assign t[147] = (t[173]);
  assign t[148] = (t[174]);
  assign t[149] = (t[175]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = (t[176]);
  assign t[151] = (t[177]);
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = t[194] ^ x[4];
  assign t[169] = t[195] ^ x[9];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[196] ^ x[12];
  assign t[171] = t[197] ^ x[15];
  assign t[172] = t[198] ^ x[18];
  assign t[173] = t[199] ^ x[21];
  assign t[174] = t[200] ^ x[24];
  assign t[175] = t[201] ^ x[27];
  assign t[176] = t[202] ^ x[30];
  assign t[177] = t[203] ^ x[33];
  assign t[178] = t[204] ^ x[36];
  assign t[179] = t[205] ^ x[39];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[42];
  assign t[181] = t[207] ^ x[47];
  assign t[182] = t[208] ^ x[50];
  assign t[183] = t[209] ^ x[55];
  assign t[184] = t[210] ^ x[58];
  assign t[185] = t[211] ^ x[61];
  assign t[186] = t[212] ^ x[66];
  assign t[187] = t[213] ^ x[69];
  assign t[188] = t[214] ^ x[78];
  assign t[189] = t[215] ^ x[81];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[84];
  assign t[191] = t[217] ^ x[87];
  assign t[192] = t[218] ^ x[90];
  assign t[193] = t[219] ^ x[99];
  assign t[194] = (t[220] & ~t[221]);
  assign t[195] = (t[222] & ~t[223]);
  assign t[196] = (t[224] & ~t[225]);
  assign t[197] = (t[226] & ~t[227]);
  assign t[198] = (t[228] & ~t[229]);
  assign t[199] = (t[230] & ~t[231]);
  assign t[19] = t[33] ^ t[4];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[232] & ~t[233]);
  assign t[201] = (t[234] & ~t[235]);
  assign t[202] = (t[236] & ~t[237]);
  assign t[203] = (t[238] & ~t[239]);
  assign t[204] = (t[240] & ~t[241]);
  assign t[205] = (t[242] & ~t[243]);
  assign t[206] = (t[244] & ~t[245]);
  assign t[207] = (t[246] & ~t[247]);
  assign t[208] = (t[248] & ~t[249]);
  assign t[209] = (t[250] & ~t[251]);
  assign t[20] = t[34] ^ t[35];
  assign t[210] = (t[252] & ~t[253]);
  assign t[211] = (t[254] & ~t[255]);
  assign t[212] = (t[256] & ~t[257]);
  assign t[213] = (t[258] & ~t[259]);
  assign t[214] = (t[260] & ~t[261]);
  assign t[215] = (t[262] & ~t[263]);
  assign t[216] = (t[264] & ~t[265]);
  assign t[217] = (t[266] & ~t[267]);
  assign t[218] = (t[268] & ~t[269]);
  assign t[219] = (t[270] & ~t[271]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = t[272] ^ x[4];
  assign t[221] = t[273] ^ x[3];
  assign t[222] = t[274] ^ x[9];
  assign t[223] = t[275] ^ x[8];
  assign t[224] = t[276] ^ x[12];
  assign t[225] = t[277] ^ x[11];
  assign t[226] = t[278] ^ x[15];
  assign t[227] = t[279] ^ x[14];
  assign t[228] = t[280] ^ x[18];
  assign t[229] = t[281] ^ x[17];
  assign t[22] = t[38] & t[39];
  assign t[230] = t[282] ^ x[21];
  assign t[231] = t[283] ^ x[20];
  assign t[232] = t[284] ^ x[24];
  assign t[233] = t[285] ^ x[23];
  assign t[234] = t[286] ^ x[27];
  assign t[235] = t[287] ^ x[26];
  assign t[236] = t[288] ^ x[30];
  assign t[237] = t[289] ^ x[29];
  assign t[238] = t[290] ^ x[33];
  assign t[239] = t[291] ^ x[32];
  assign t[23] = t[40] ? t[41] : t[143];
  assign t[240] = t[292] ^ x[36];
  assign t[241] = t[293] ^ x[35];
  assign t[242] = t[294] ^ x[39];
  assign t[243] = t[295] ^ x[38];
  assign t[244] = t[296] ^ x[42];
  assign t[245] = t[297] ^ x[41];
  assign t[246] = t[298] ^ x[47];
  assign t[247] = t[299] ^ x[46];
  assign t[248] = t[300] ^ x[50];
  assign t[249] = t[301] ^ x[49];
  assign t[24] = t[42] ^ t[43];
  assign t[250] = t[302] ^ x[55];
  assign t[251] = t[303] ^ x[54];
  assign t[252] = t[304] ^ x[58];
  assign t[253] = t[305] ^ x[57];
  assign t[254] = t[306] ^ x[61];
  assign t[255] = t[307] ^ x[60];
  assign t[256] = t[308] ^ x[66];
  assign t[257] = t[309] ^ x[65];
  assign t[258] = t[310] ^ x[69];
  assign t[259] = t[311] ^ x[68];
  assign t[25] = t[144] ^ t[44];
  assign t[260] = t[312] ^ x[78];
  assign t[261] = t[313] ^ x[77];
  assign t[262] = t[314] ^ x[81];
  assign t[263] = t[315] ^ x[80];
  assign t[264] = t[316] ^ x[84];
  assign t[265] = t[317] ^ x[83];
  assign t[266] = t[318] ^ x[87];
  assign t[267] = t[319] ^ x[86];
  assign t[268] = t[320] ^ x[90];
  assign t[269] = t[321] ^ x[89];
  assign t[26] = t[45] ^ t[46];
  assign t[270] = t[322] ^ x[99];
  assign t[271] = t[323] ^ x[98];
  assign t[272] = (x[2]);
  assign t[273] = (x[2]);
  assign t[274] = (x[7]);
  assign t[275] = (x[7]);
  assign t[276] = (x[10]);
  assign t[277] = (x[10]);
  assign t[278] = (x[13]);
  assign t[279] = (x[13]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (x[16]);
  assign t[281] = (x[16]);
  assign t[282] = (x[19]);
  assign t[283] = (x[19]);
  assign t[284] = (x[22]);
  assign t[285] = (x[22]);
  assign t[286] = (x[25]);
  assign t[287] = (x[25]);
  assign t[288] = (x[28]);
  assign t[289] = (x[28]);
  assign t[28] = ~(t[49]);
  assign t[290] = (x[31]);
  assign t[291] = (x[31]);
  assign t[292] = (x[34]);
  assign t[293] = (x[34]);
  assign t[294] = (x[37]);
  assign t[295] = (x[37]);
  assign t[296] = (x[40]);
  assign t[297] = (x[40]);
  assign t[298] = (x[45]);
  assign t[299] = (x[45]);
  assign t[29] = ~(t[145]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[48]);
  assign t[301] = (x[48]);
  assign t[302] = (x[53]);
  assign t[303] = (x[53]);
  assign t[304] = (x[56]);
  assign t[305] = (x[56]);
  assign t[306] = (x[59]);
  assign t[307] = (x[59]);
  assign t[308] = (x[64]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[146]);
  assign t[310] = (x[67]);
  assign t[311] = (x[67]);
  assign t[312] = (x[76]);
  assign t[313] = (x[76]);
  assign t[314] = (x[79]);
  assign t[315] = (x[79]);
  assign t[316] = (x[82]);
  assign t[317] = (x[82]);
  assign t[318] = (x[85]);
  assign t[319] = (x[85]);
  assign t[31] = ~(t[147]);
  assign t[320] = (x[88]);
  assign t[321] = (x[88]);
  assign t[322] = (x[97]);
  assign t[323] = (x[97]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[33] = t[8] ? t[52] : t[148];
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[55] & t[56];
  assign t[36] = ~t[57];
  assign t[37] = ~t[58];
  assign t[38] = ~(t[59]);
  assign t[39] = t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[15]);
  assign t[41] = t[143] ^ t[61];
  assign t[42] = t[62] ^ t[63];
  assign t[43] = t[64] & t[65];
  assign t[44] = t[40] ? t[66] : t[149];
  assign t[45] = t[67] ^ t[68];
  assign t[46] = t[69] & t[70];
  assign t[47] = ~(t[71] & t[72]);
  assign t[48] = t[150] | t[73];
  assign t[49] = ~(t[74]);
  assign t[4] = t[8] ? t[9] : t[142];
  assign t[50] = ~(t[151]);
  assign t[51] = ~(t[75] & t[144]);
  assign t[52] = t[148] ^ t[76];
  assign t[53] = t[77] & t[78];
  assign t[54] = t[79] & t[80];
  assign t[55] = ~(t[53] ^ t[81]);
  assign t[56] = t[82] ^ t[83];
  assign t[57] = t[27] ? t[84] : t[152];
  assign t[58] = t[27] ? t[85] : t[153];
  assign t[59] = t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[27] ? t[87] : t[154];
  assign t[61] = t[88] ? x[44] : x[43];
  assign t[62] = t[89] & t[90];
  assign t[63] = t[91] & t[92];
  assign t[64] = ~(t[93] ^ t[42]);
  assign t[65] = t[94] ^ t[92];
  assign t[66] = t[149] ^ t[95];
  assign t[67] = t[96] & t[97];
  assign t[68] = t[98] & t[99];
  assign t[69] = ~(t[100] ^ t[45]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[101] ^ t[99];
  assign t[71] = ~(t[73] & t[102]);
  assign t[72] = ~(t[155] ^ t[103]);
  assign t[73] = ~(t[104] & t[105]);
  assign t[74] = ~(t[48]);
  assign t[75] = ~(t[156]);
  assign t[76] = t[28] ? x[52] : x[51];
  assign t[77] = ~(t[83]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[33]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[107] : t[157];
  assign t[81] = t[19] ^ t[106];
  assign t[82] = t[106] ^ t[4];
  assign t[83] = t[80] ^ t[33];
  assign t[84] = t[152] ^ t[108];
  assign t[85] = t[153] ^ t[109];
  assign t[86] = t[27] ? t[110] : t[158];
  assign t[87] = t[154] ^ t[111];
  assign t[88] = ~(t[49]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[113]);
  assign t[91] = ~(t[114]);
  assign t[92] = t[40] ? t[115] : t[159];
  assign t[93] = t[113] ^ t[114];
  assign t[94] = t[114] ^ t[23];
  assign t[95] = t[74] ? x[63] : x[62];
  assign t[96] = ~(t[116]);
  assign t[97] = ~(t[117]);
  assign t[98] = ~(t[118]);
  assign t[99] = t[146] ^ t[119];
  assign t[9] = t[142] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind49(x, y);
 input [111:0] x;
 output y;

 wire [323:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[117] ^ t[118];
  assign t[101] = t[118] ^ t[25];
  assign t[102] = ~(t[120] & t[121]);
  assign t[103] = t[122] ^ t[160];
  assign t[104] = ~(t[155]);
  assign t[105] = t[123] & t[122];
  assign t[106] = t[8] ? t[124] : t[161];
  assign t[107] = t[157] ^ t[125];
  assign t[108] = t[74] ? x[71] : x[70];
  assign t[109] = t[74] ? x[73] : x[72];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[158] ^ t[126];
  assign t[111] = t[88] ? x[75] : x[74];
  assign t[112] = t[92] ^ t[114];
  assign t[113] = t[40] ? t[127] : t[162];
  assign t[114] = t[40] ? t[128] : t[163];
  assign t[115] = t[159] ^ t[129];
  assign t[116] = t[99] ^ t[118];
  assign t[117] = t[40] ? t[130] : t[164];
  assign t[118] = t[145] ^ t[131];
  assign t[119] = t[40] ? t[132] : t[165];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[123] | t[122]);
  assign t[121] = ~(t[133] | t[104]);
  assign t[122] = ~(t[166]);
  assign t[123] = ~(t[160]);
  assign t[124] = t[161] ^ t[134];
  assign t[125] = t[28] ? x[92] : x[91];
  assign t[126] = t[135] ? x[94] : x[93];
  assign t[127] = t[162] ^ t[136];
  assign t[128] = t[163] ^ t[137];
  assign t[129] = t[88] ? x[96] : x[95];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[164] ^ t[138];
  assign t[131] = t[27] ? t[139] : t[167];
  assign t[132] = t[165] ^ t[140];
  assign t[133] = ~(t[150]);
  assign t[134] = t[28] ? x[101] : x[100];
  assign t[135] = ~(t[49]);
  assign t[136] = t[88] ? x[103] : x[102];
  assign t[137] = t[88] ? x[105] : x[104];
  assign t[138] = t[74] ? x[107] : x[106];
  assign t[139] = t[167] ^ t[141];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[135] ? x[109] : x[108];
  assign t[141] = t[135] ? x[111] : x[110];
  assign t[142] = (t[168]);
  assign t[143] = (t[169]);
  assign t[144] = (t[170]);
  assign t[145] = (t[171]);
  assign t[146] = (t[172]);
  assign t[147] = (t[173]);
  assign t[148] = (t[174]);
  assign t[149] = (t[175]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = (t[176]);
  assign t[151] = (t[177]);
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = t[194] ^ x[4];
  assign t[169] = t[195] ^ x[9];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[196] ^ x[12];
  assign t[171] = t[197] ^ x[15];
  assign t[172] = t[198] ^ x[18];
  assign t[173] = t[199] ^ x[21];
  assign t[174] = t[200] ^ x[24];
  assign t[175] = t[201] ^ x[27];
  assign t[176] = t[202] ^ x[30];
  assign t[177] = t[203] ^ x[33];
  assign t[178] = t[204] ^ x[36];
  assign t[179] = t[205] ^ x[39];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[42];
  assign t[181] = t[207] ^ x[47];
  assign t[182] = t[208] ^ x[50];
  assign t[183] = t[209] ^ x[55];
  assign t[184] = t[210] ^ x[58];
  assign t[185] = t[211] ^ x[61];
  assign t[186] = t[212] ^ x[66];
  assign t[187] = t[213] ^ x[69];
  assign t[188] = t[214] ^ x[78];
  assign t[189] = t[215] ^ x[81];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[84];
  assign t[191] = t[217] ^ x[87];
  assign t[192] = t[218] ^ x[90];
  assign t[193] = t[219] ^ x[99];
  assign t[194] = (t[220] & ~t[221]);
  assign t[195] = (t[222] & ~t[223]);
  assign t[196] = (t[224] & ~t[225]);
  assign t[197] = (t[226] & ~t[227]);
  assign t[198] = (t[228] & ~t[229]);
  assign t[199] = (t[230] & ~t[231]);
  assign t[19] = t[33] ^ t[4];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[232] & ~t[233]);
  assign t[201] = (t[234] & ~t[235]);
  assign t[202] = (t[236] & ~t[237]);
  assign t[203] = (t[238] & ~t[239]);
  assign t[204] = (t[240] & ~t[241]);
  assign t[205] = (t[242] & ~t[243]);
  assign t[206] = (t[244] & ~t[245]);
  assign t[207] = (t[246] & ~t[247]);
  assign t[208] = (t[248] & ~t[249]);
  assign t[209] = (t[250] & ~t[251]);
  assign t[20] = t[34] ^ t[35];
  assign t[210] = (t[252] & ~t[253]);
  assign t[211] = (t[254] & ~t[255]);
  assign t[212] = (t[256] & ~t[257]);
  assign t[213] = (t[258] & ~t[259]);
  assign t[214] = (t[260] & ~t[261]);
  assign t[215] = (t[262] & ~t[263]);
  assign t[216] = (t[264] & ~t[265]);
  assign t[217] = (t[266] & ~t[267]);
  assign t[218] = (t[268] & ~t[269]);
  assign t[219] = (t[270] & ~t[271]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = t[272] ^ x[4];
  assign t[221] = t[273] ^ x[3];
  assign t[222] = t[274] ^ x[9];
  assign t[223] = t[275] ^ x[8];
  assign t[224] = t[276] ^ x[12];
  assign t[225] = t[277] ^ x[11];
  assign t[226] = t[278] ^ x[15];
  assign t[227] = t[279] ^ x[14];
  assign t[228] = t[280] ^ x[18];
  assign t[229] = t[281] ^ x[17];
  assign t[22] = t[38] & t[39];
  assign t[230] = t[282] ^ x[21];
  assign t[231] = t[283] ^ x[20];
  assign t[232] = t[284] ^ x[24];
  assign t[233] = t[285] ^ x[23];
  assign t[234] = t[286] ^ x[27];
  assign t[235] = t[287] ^ x[26];
  assign t[236] = t[288] ^ x[30];
  assign t[237] = t[289] ^ x[29];
  assign t[238] = t[290] ^ x[33];
  assign t[239] = t[291] ^ x[32];
  assign t[23] = t[40] ? t[41] : t[143];
  assign t[240] = t[292] ^ x[36];
  assign t[241] = t[293] ^ x[35];
  assign t[242] = t[294] ^ x[39];
  assign t[243] = t[295] ^ x[38];
  assign t[244] = t[296] ^ x[42];
  assign t[245] = t[297] ^ x[41];
  assign t[246] = t[298] ^ x[47];
  assign t[247] = t[299] ^ x[46];
  assign t[248] = t[300] ^ x[50];
  assign t[249] = t[301] ^ x[49];
  assign t[24] = t[42] ^ t[43];
  assign t[250] = t[302] ^ x[55];
  assign t[251] = t[303] ^ x[54];
  assign t[252] = t[304] ^ x[58];
  assign t[253] = t[305] ^ x[57];
  assign t[254] = t[306] ^ x[61];
  assign t[255] = t[307] ^ x[60];
  assign t[256] = t[308] ^ x[66];
  assign t[257] = t[309] ^ x[65];
  assign t[258] = t[310] ^ x[69];
  assign t[259] = t[311] ^ x[68];
  assign t[25] = t[144] ^ t[44];
  assign t[260] = t[312] ^ x[78];
  assign t[261] = t[313] ^ x[77];
  assign t[262] = t[314] ^ x[81];
  assign t[263] = t[315] ^ x[80];
  assign t[264] = t[316] ^ x[84];
  assign t[265] = t[317] ^ x[83];
  assign t[266] = t[318] ^ x[87];
  assign t[267] = t[319] ^ x[86];
  assign t[268] = t[320] ^ x[90];
  assign t[269] = t[321] ^ x[89];
  assign t[26] = t[45] ^ t[46];
  assign t[270] = t[322] ^ x[99];
  assign t[271] = t[323] ^ x[98];
  assign t[272] = (x[2]);
  assign t[273] = (x[2]);
  assign t[274] = (x[7]);
  assign t[275] = (x[7]);
  assign t[276] = (x[10]);
  assign t[277] = (x[10]);
  assign t[278] = (x[13]);
  assign t[279] = (x[13]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (x[16]);
  assign t[281] = (x[16]);
  assign t[282] = (x[19]);
  assign t[283] = (x[19]);
  assign t[284] = (x[22]);
  assign t[285] = (x[22]);
  assign t[286] = (x[25]);
  assign t[287] = (x[25]);
  assign t[288] = (x[28]);
  assign t[289] = (x[28]);
  assign t[28] = ~(t[49]);
  assign t[290] = (x[31]);
  assign t[291] = (x[31]);
  assign t[292] = (x[34]);
  assign t[293] = (x[34]);
  assign t[294] = (x[37]);
  assign t[295] = (x[37]);
  assign t[296] = (x[40]);
  assign t[297] = (x[40]);
  assign t[298] = (x[45]);
  assign t[299] = (x[45]);
  assign t[29] = ~(t[145]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[48]);
  assign t[301] = (x[48]);
  assign t[302] = (x[53]);
  assign t[303] = (x[53]);
  assign t[304] = (x[56]);
  assign t[305] = (x[56]);
  assign t[306] = (x[59]);
  assign t[307] = (x[59]);
  assign t[308] = (x[64]);
  assign t[309] = (x[64]);
  assign t[30] = ~(t[146]);
  assign t[310] = (x[67]);
  assign t[311] = (x[67]);
  assign t[312] = (x[76]);
  assign t[313] = (x[76]);
  assign t[314] = (x[79]);
  assign t[315] = (x[79]);
  assign t[316] = (x[82]);
  assign t[317] = (x[82]);
  assign t[318] = (x[85]);
  assign t[319] = (x[85]);
  assign t[31] = ~(t[147]);
  assign t[320] = (x[88]);
  assign t[321] = (x[88]);
  assign t[322] = (x[97]);
  assign t[323] = (x[97]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[33] = t[8] ? t[52] : t[148];
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[55] & t[56];
  assign t[36] = ~t[57];
  assign t[37] = ~t[58];
  assign t[38] = ~(t[59]);
  assign t[39] = t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[15]);
  assign t[41] = t[143] ^ t[61];
  assign t[42] = t[62] ^ t[63];
  assign t[43] = t[64] & t[65];
  assign t[44] = t[40] ? t[66] : t[149];
  assign t[45] = t[67] ^ t[68];
  assign t[46] = t[69] & t[70];
  assign t[47] = ~(t[71] & t[72]);
  assign t[48] = t[150] | t[73];
  assign t[49] = ~(t[74]);
  assign t[4] = t[8] ? t[9] : t[142];
  assign t[50] = ~(t[151]);
  assign t[51] = ~(t[75] & t[144]);
  assign t[52] = t[148] ^ t[76];
  assign t[53] = t[77] & t[78];
  assign t[54] = t[79] & t[80];
  assign t[55] = ~(t[53] ^ t[81]);
  assign t[56] = t[82] ^ t[83];
  assign t[57] = t[27] ? t[84] : t[152];
  assign t[58] = t[27] ? t[85] : t[153];
  assign t[59] = t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[27] ? t[87] : t[154];
  assign t[61] = t[88] ? x[44] : x[43];
  assign t[62] = t[89] & t[90];
  assign t[63] = t[91] & t[92];
  assign t[64] = ~(t[93] ^ t[42]);
  assign t[65] = t[94] ^ t[92];
  assign t[66] = t[149] ^ t[95];
  assign t[67] = t[96] & t[97];
  assign t[68] = t[98] & t[99];
  assign t[69] = ~(t[100] ^ t[45]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[101] ^ t[99];
  assign t[71] = ~(t[73] & t[102]);
  assign t[72] = ~(t[155] ^ t[103]);
  assign t[73] = ~(t[104] & t[105]);
  assign t[74] = ~(t[48]);
  assign t[75] = ~(t[156]);
  assign t[76] = t[28] ? x[52] : x[51];
  assign t[77] = ~(t[83]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[33]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[107] : t[157];
  assign t[81] = t[19] ^ t[106];
  assign t[82] = t[106] ^ t[4];
  assign t[83] = t[80] ^ t[33];
  assign t[84] = t[152] ^ t[108];
  assign t[85] = t[153] ^ t[109];
  assign t[86] = t[27] ? t[110] : t[158];
  assign t[87] = t[154] ^ t[111];
  assign t[88] = ~(t[49]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[113]);
  assign t[91] = ~(t[114]);
  assign t[92] = t[40] ? t[115] : t[159];
  assign t[93] = t[113] ^ t[114];
  assign t[94] = t[114] ^ t[23];
  assign t[95] = t[74] ? x[63] : x[62];
  assign t[96] = ~(t[116]);
  assign t[97] = ~(t[117]);
  assign t[98] = ~(t[118]);
  assign t[99] = t[146] ^ t[119];
  assign t[9] = t[142] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [111:0] x;
 output y;

 wire [345:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[41] ^ t[66];
  assign t[101] = t[66] ^ t[25];
  assign t[102] = ~(t[132] & t[133]);
  assign t[103] = t[134] ^ t[182];
  assign t[104] = ~(t[178]);
  assign t[105] = t[135] & t[134];
  assign t[106] = ~(t[49]);
  assign t[107] = ~(t[136]);
  assign t[108] = ~(t[56]);
  assign t[109] = t[56] ^ t[82];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[82] ^ t[33];
  assign t[111] = t[106] ? x[68] : x[67];
  assign t[112] = t[180] ^ t[137];
  assign t[113] = t[106] ? x[70] : x[69];
  assign t[114] = t[27] ? t[138] : t[183];
  assign t[115] = t[27] ? t[139] : t[184];
  assign t[116] = t[140] ^ t[141];
  assign t[117] = t[85] ^ t[142];
  assign t[118] = t[143];
  assign t[119] = t[28] ? x[78] : x[77];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[144] ^ t[63]);
  assign t[121] = t[39] ^ t[125];
  assign t[122] = ~(t[128]);
  assign t[123] = ~(t[145]);
  assign t[124] = ~(t[4]);
  assign t[125] = t[8] ? t[146] : t[185];
  assign t[126] = t[39] ^ t[145];
  assign t[127] = t[145] ^ t[61];
  assign t[128] = t[125] ^ t[4];
  assign t[129] = t[181] ^ t[147];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[148] ? x[83] : x[82];
  assign t[131] = t[43] ^ t[66];
  assign t[132] = ~(t[135] | t[134]);
  assign t[133] = ~(t[149] | t[104]);
  assign t[134] = ~(t[186]);
  assign t[135] = ~(t[182]);
  assign t[136] = t[58] ^ t[82];
  assign t[137] = t[106] ? x[88] : x[87];
  assign t[138] = t[183] ^ t[150];
  assign t[139] = t[184] ^ t[151];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[152] & t[153];
  assign t[141] = t[154] & t[118];
  assign t[142] = ~t[155];
  assign t[143] = t[27] ? t[156] : t[187];
  assign t[144] = t[145] ^ t[4];
  assign t[145] = t[8] ? t[157] : t[188];
  assign t[146] = t[185] ^ t[158];
  assign t[147] = t[148] ? x[96] : x[95];
  assign t[148] = ~(t[49]);
  assign t[149] = ~(t[172]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[75] ? x[98] : x[97];
  assign t[151] = t[148] ? x[100] : x[99];
  assign t[152] = ~(t[159]);
  assign t[153] = ~(t[84]);
  assign t[154] = ~(t[85]);
  assign t[155] = t[27] ? t[160] : t[189];
  assign t[156] = t[187] ^ t[161];
  assign t[157] = t[188] ^ t[162];
  assign t[158] = t[28] ? x[105] : x[104];
  assign t[159] = t[118] ^ t[85];
  assign t[15] = ~(t[27]);
  assign t[160] = t[189] ^ t[163];
  assign t[161] = t[106] ? x[107] : x[106];
  assign t[162] = t[28] ? x[109] : x[108];
  assign t[163] = t[75] ? x[111] : x[110];
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = (t[205]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[206]);
  assign t[181] = (t[207]);
  assign t[182] = (t[208]);
  assign t[183] = (t[209]);
  assign t[184] = (t[210]);
  assign t[185] = (t[211]);
  assign t[186] = (t[212]);
  assign t[187] = (t[213]);
  assign t[188] = (t[214]);
  assign t[189] = (t[215]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[4];
  assign t[191] = t[217] ^ x[9];
  assign t[192] = t[218] ^ x[12];
  assign t[193] = t[219] ^ x[15];
  assign t[194] = t[220] ^ x[18];
  assign t[195] = t[221] ^ x[21];
  assign t[196] = t[222] ^ x[24];
  assign t[197] = t[223] ^ x[27];
  assign t[198] = t[224] ^ x[30];
  assign t[199] = t[225] ^ x[33];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[36];
  assign t[201] = t[227] ^ x[39];
  assign t[202] = t[228] ^ x[42];
  assign t[203] = t[229] ^ x[45];
  assign t[204] = t[230] ^ x[48];
  assign t[205] = t[231] ^ x[51];
  assign t[206] = t[232] ^ x[56];
  assign t[207] = t[233] ^ x[61];
  assign t[208] = t[234] ^ x[66];
  assign t[209] = t[235] ^ x[73];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[236] ^ x[76];
  assign t[211] = t[237] ^ x[81];
  assign t[212] = t[238] ^ x[86];
  assign t[213] = t[239] ^ x[91];
  assign t[214] = t[240] ^ x[94];
  assign t[215] = t[241] ^ x[103];
  assign t[216] = (t[242] & ~t[243]);
  assign t[217] = (t[244] & ~t[245]);
  assign t[218] = (t[246] & ~t[247]);
  assign t[219] = (t[248] & ~t[249]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[250] & ~t[251]);
  assign t[221] = (t[252] & ~t[253]);
  assign t[222] = (t[254] & ~t[255]);
  assign t[223] = (t[256] & ~t[257]);
  assign t[224] = (t[258] & ~t[259]);
  assign t[225] = (t[260] & ~t[261]);
  assign t[226] = (t[262] & ~t[263]);
  assign t[227] = (t[264] & ~t[265]);
  assign t[228] = (t[266] & ~t[267]);
  assign t[229] = (t[268] & ~t[269]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[270] & ~t[271]);
  assign t[231] = (t[272] & ~t[273]);
  assign t[232] = (t[274] & ~t[275]);
  assign t[233] = (t[276] & ~t[277]);
  assign t[234] = (t[278] & ~t[279]);
  assign t[235] = (t[280] & ~t[281]);
  assign t[236] = (t[282] & ~t[283]);
  assign t[237] = (t[284] & ~t[285]);
  assign t[238] = (t[286] & ~t[287]);
  assign t[239] = (t[288] & ~t[289]);
  assign t[23] = t[41] ^ t[25];
  assign t[240] = (t[290] & ~t[291]);
  assign t[241] = (t[292] & ~t[293]);
  assign t[242] = t[294] ^ x[4];
  assign t[243] = t[295] ^ x[3];
  assign t[244] = t[296] ^ x[9];
  assign t[245] = t[297] ^ x[8];
  assign t[246] = t[298] ^ x[12];
  assign t[247] = t[299] ^ x[11];
  assign t[248] = t[300] ^ x[15];
  assign t[249] = t[301] ^ x[14];
  assign t[24] = t[42] & t[43];
  assign t[250] = t[302] ^ x[18];
  assign t[251] = t[303] ^ x[17];
  assign t[252] = t[304] ^ x[21];
  assign t[253] = t[305] ^ x[20];
  assign t[254] = t[306] ^ x[24];
  assign t[255] = t[307] ^ x[23];
  assign t[256] = t[308] ^ x[27];
  assign t[257] = t[309] ^ x[26];
  assign t[258] = t[310] ^ x[30];
  assign t[259] = t[311] ^ x[29];
  assign t[25] = t[165] ^ t[44];
  assign t[260] = t[312] ^ x[33];
  assign t[261] = t[313] ^ x[32];
  assign t[262] = t[314] ^ x[36];
  assign t[263] = t[315] ^ x[35];
  assign t[264] = t[316] ^ x[39];
  assign t[265] = t[317] ^ x[38];
  assign t[266] = t[318] ^ x[42];
  assign t[267] = t[319] ^ x[41];
  assign t[268] = t[320] ^ x[45];
  assign t[269] = t[321] ^ x[44];
  assign t[26] = t[45] ^ t[46];
  assign t[270] = t[322] ^ x[48];
  assign t[271] = t[323] ^ x[47];
  assign t[272] = t[324] ^ x[51];
  assign t[273] = t[325] ^ x[50];
  assign t[274] = t[326] ^ x[56];
  assign t[275] = t[327] ^ x[55];
  assign t[276] = t[328] ^ x[61];
  assign t[277] = t[329] ^ x[60];
  assign t[278] = t[330] ^ x[66];
  assign t[279] = t[331] ^ x[65];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[332] ^ x[73];
  assign t[281] = t[333] ^ x[72];
  assign t[282] = t[334] ^ x[76];
  assign t[283] = t[335] ^ x[75];
  assign t[284] = t[336] ^ x[81];
  assign t[285] = t[337] ^ x[80];
  assign t[286] = t[338] ^ x[86];
  assign t[287] = t[339] ^ x[85];
  assign t[288] = t[340] ^ x[91];
  assign t[289] = t[341] ^ x[90];
  assign t[28] = ~(t[49]);
  assign t[290] = t[342] ^ x[94];
  assign t[291] = t[343] ^ x[93];
  assign t[292] = t[344] ^ x[103];
  assign t[293] = t[345] ^ x[102];
  assign t[294] = (x[2]);
  assign t[295] = (x[2]);
  assign t[296] = (x[7]);
  assign t[297] = (x[7]);
  assign t[298] = (x[10]);
  assign t[299] = (x[10]);
  assign t[29] = ~(t[166]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[13]);
  assign t[301] = (x[13]);
  assign t[302] = (x[16]);
  assign t[303] = (x[16]);
  assign t[304] = (x[19]);
  assign t[305] = (x[19]);
  assign t[306] = (x[22]);
  assign t[307] = (x[22]);
  assign t[308] = (x[25]);
  assign t[309] = (x[25]);
  assign t[30] = ~(t[167]);
  assign t[310] = (x[28]);
  assign t[311] = (x[28]);
  assign t[312] = (x[31]);
  assign t[313] = (x[31]);
  assign t[314] = (x[34]);
  assign t[315] = (x[34]);
  assign t[316] = (x[37]);
  assign t[317] = (x[37]);
  assign t[318] = (x[40]);
  assign t[319] = (x[40]);
  assign t[31] = ~(t[168]);
  assign t[320] = (x[43]);
  assign t[321] = (x[43]);
  assign t[322] = (x[46]);
  assign t[323] = (x[46]);
  assign t[324] = (x[49]);
  assign t[325] = (x[49]);
  assign t[326] = (x[54]);
  assign t[327] = (x[54]);
  assign t[328] = (x[59]);
  assign t[329] = (x[59]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[64]);
  assign t[331] = (x[64]);
  assign t[332] = (x[71]);
  assign t[333] = (x[71]);
  assign t[334] = (x[74]);
  assign t[335] = (x[74]);
  assign t[336] = (x[79]);
  assign t[337] = (x[79]);
  assign t[338] = (x[84]);
  assign t[339] = (x[84]);
  assign t[33] = t[52] ? t[53] : t[169];
  assign t[340] = (x[89]);
  assign t[341] = (x[89]);
  assign t[342] = (x[92]);
  assign t[343] = (x[92]);
  assign t[344] = (x[101]);
  assign t[345] = (x[101]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] ^ t[33];
  assign t[36] = t[57] & t[58];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[4] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[52] ? t[65] : t[170];
  assign t[42] = ~(t[66]);
  assign t[43] = t[167] ^ t[67];
  assign t[44] = t[52] ? t[68] : t[171];
  assign t[45] = t[69] ^ t[24];
  assign t[46] = t[70] & t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[172] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = t[8] ? t[9] : t[164];
  assign t[50] = ~(t[173]);
  assign t[51] = ~(t[76] & t[165]);
  assign t[52] = ~(t[15]);
  assign t[53] = t[169] ^ t[77];
  assign t[54] = t[78] ^ t[36];
  assign t[55] = t[79] & t[80];
  assign t[56] = t[52] ? t[81] : t[174];
  assign t[57] = ~(t[82]);
  assign t[58] = t[52] ? t[83] : t[175];
  assign t[59] = t[84] ^ t[85];
  assign t[5] = ~(t[10]);
  assign t[60] = t[86] & t[87];
  assign t[61] = t[8] ? t[88] : t[176];
  assign t[62] = t[63] ^ t[89];
  assign t[63] = t[90] ^ t[91];
  assign t[64] = t[92] & t[93];
  assign t[65] = t[170] ^ t[94];
  assign t[66] = t[166] ^ t[95];
  assign t[67] = t[52] ? t[96] : t[177];
  assign t[68] = t[171] ^ t[97];
  assign t[69] = t[98] & t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[100] ^ t[45]);
  assign t[71] = t[101] ^ t[43];
  assign t[72] = ~(t[74] & t[102]);
  assign t[73] = ~(t[178] ^ t[103]);
  assign t[74] = ~(t[104] & t[105]);
  assign t[75] = ~(t[48]);
  assign t[76] = ~(t[179]);
  assign t[77] = t[106] ? x[53] : x[52];
  assign t[78] = t[107] & t[108];
  assign t[79] = ~(t[109] ^ t[54]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[110] ^ t[58];
  assign t[81] = t[174] ^ t[111];
  assign t[82] = t[52] ? t[112] : t[180];
  assign t[83] = t[175] ^ t[113];
  assign t[84] = ~t[114];
  assign t[85] = t[115];
  assign t[86] = ~(t[59] ^ t[116]);
  assign t[87] = t[117] ^ t[118];
  assign t[88] = t[176] ^ t[119];
  assign t[89] = t[120] & t[121];
  assign t[8] = ~(t[15]);
  assign t[90] = t[122] & t[123];
  assign t[91] = t[124] & t[125];
  assign t[92] = ~(t[90] ^ t[126]);
  assign t[93] = t[127] ^ t[128];
  assign t[94] = t[75] ? x[58] : x[57];
  assign t[95] = t[27] ? t[129] : t[181];
  assign t[96] = t[177] ^ t[130];
  assign t[97] = t[75] ? x[63] : x[62];
  assign t[98] = ~(t[131]);
  assign t[99] = ~(t[41]);
  assign t[9] = t[164] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind51(x, y);
 input [111:0] x;
 output y;

 wire [345:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[41] ^ t[66];
  assign t[101] = t[66] ^ t[25];
  assign t[102] = ~(t[132] & t[133]);
  assign t[103] = t[134] ^ t[182];
  assign t[104] = ~(t[178]);
  assign t[105] = t[135] & t[134];
  assign t[106] = ~(t[49]);
  assign t[107] = ~(t[136]);
  assign t[108] = ~(t[56]);
  assign t[109] = t[56] ^ t[82];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[82] ^ t[33];
  assign t[111] = t[106] ? x[68] : x[67];
  assign t[112] = t[180] ^ t[137];
  assign t[113] = t[106] ? x[70] : x[69];
  assign t[114] = t[27] ? t[138] : t[183];
  assign t[115] = t[27] ? t[139] : t[184];
  assign t[116] = t[140] ^ t[141];
  assign t[117] = t[85] ^ t[142];
  assign t[118] = t[143];
  assign t[119] = t[28] ? x[78] : x[77];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[144] ^ t[63]);
  assign t[121] = t[39] ^ t[125];
  assign t[122] = ~(t[128]);
  assign t[123] = ~(t[145]);
  assign t[124] = ~(t[4]);
  assign t[125] = t[8] ? t[146] : t[185];
  assign t[126] = t[39] ^ t[145];
  assign t[127] = t[145] ^ t[61];
  assign t[128] = t[125] ^ t[4];
  assign t[129] = t[181] ^ t[147];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[148] ? x[83] : x[82];
  assign t[131] = t[43] ^ t[66];
  assign t[132] = ~(t[135] | t[134]);
  assign t[133] = ~(t[149] | t[104]);
  assign t[134] = ~(t[186]);
  assign t[135] = ~(t[182]);
  assign t[136] = t[58] ^ t[82];
  assign t[137] = t[106] ? x[88] : x[87];
  assign t[138] = t[183] ^ t[150];
  assign t[139] = t[184] ^ t[151];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[152] & t[153];
  assign t[141] = t[154] & t[118];
  assign t[142] = ~t[155];
  assign t[143] = t[27] ? t[156] : t[187];
  assign t[144] = t[145] ^ t[4];
  assign t[145] = t[8] ? t[157] : t[188];
  assign t[146] = t[185] ^ t[158];
  assign t[147] = t[148] ? x[96] : x[95];
  assign t[148] = ~(t[49]);
  assign t[149] = ~(t[172]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[75] ? x[98] : x[97];
  assign t[151] = t[148] ? x[100] : x[99];
  assign t[152] = ~(t[159]);
  assign t[153] = ~(t[84]);
  assign t[154] = ~(t[85]);
  assign t[155] = t[27] ? t[160] : t[189];
  assign t[156] = t[187] ^ t[161];
  assign t[157] = t[188] ^ t[162];
  assign t[158] = t[28] ? x[105] : x[104];
  assign t[159] = t[118] ^ t[85];
  assign t[15] = ~(t[27]);
  assign t[160] = t[189] ^ t[163];
  assign t[161] = t[106] ? x[107] : x[106];
  assign t[162] = t[28] ? x[109] : x[108];
  assign t[163] = t[75] ? x[111] : x[110];
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = (t[205]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[206]);
  assign t[181] = (t[207]);
  assign t[182] = (t[208]);
  assign t[183] = (t[209]);
  assign t[184] = (t[210]);
  assign t[185] = (t[211]);
  assign t[186] = (t[212]);
  assign t[187] = (t[213]);
  assign t[188] = (t[214]);
  assign t[189] = (t[215]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[4];
  assign t[191] = t[217] ^ x[9];
  assign t[192] = t[218] ^ x[12];
  assign t[193] = t[219] ^ x[15];
  assign t[194] = t[220] ^ x[18];
  assign t[195] = t[221] ^ x[21];
  assign t[196] = t[222] ^ x[24];
  assign t[197] = t[223] ^ x[27];
  assign t[198] = t[224] ^ x[30];
  assign t[199] = t[225] ^ x[33];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[36];
  assign t[201] = t[227] ^ x[39];
  assign t[202] = t[228] ^ x[42];
  assign t[203] = t[229] ^ x[45];
  assign t[204] = t[230] ^ x[48];
  assign t[205] = t[231] ^ x[51];
  assign t[206] = t[232] ^ x[56];
  assign t[207] = t[233] ^ x[61];
  assign t[208] = t[234] ^ x[66];
  assign t[209] = t[235] ^ x[73];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[236] ^ x[76];
  assign t[211] = t[237] ^ x[81];
  assign t[212] = t[238] ^ x[86];
  assign t[213] = t[239] ^ x[91];
  assign t[214] = t[240] ^ x[94];
  assign t[215] = t[241] ^ x[103];
  assign t[216] = (t[242] & ~t[243]);
  assign t[217] = (t[244] & ~t[245]);
  assign t[218] = (t[246] & ~t[247]);
  assign t[219] = (t[248] & ~t[249]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[250] & ~t[251]);
  assign t[221] = (t[252] & ~t[253]);
  assign t[222] = (t[254] & ~t[255]);
  assign t[223] = (t[256] & ~t[257]);
  assign t[224] = (t[258] & ~t[259]);
  assign t[225] = (t[260] & ~t[261]);
  assign t[226] = (t[262] & ~t[263]);
  assign t[227] = (t[264] & ~t[265]);
  assign t[228] = (t[266] & ~t[267]);
  assign t[229] = (t[268] & ~t[269]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[270] & ~t[271]);
  assign t[231] = (t[272] & ~t[273]);
  assign t[232] = (t[274] & ~t[275]);
  assign t[233] = (t[276] & ~t[277]);
  assign t[234] = (t[278] & ~t[279]);
  assign t[235] = (t[280] & ~t[281]);
  assign t[236] = (t[282] & ~t[283]);
  assign t[237] = (t[284] & ~t[285]);
  assign t[238] = (t[286] & ~t[287]);
  assign t[239] = (t[288] & ~t[289]);
  assign t[23] = t[41] ^ t[25];
  assign t[240] = (t[290] & ~t[291]);
  assign t[241] = (t[292] & ~t[293]);
  assign t[242] = t[294] ^ x[4];
  assign t[243] = t[295] ^ x[3];
  assign t[244] = t[296] ^ x[9];
  assign t[245] = t[297] ^ x[8];
  assign t[246] = t[298] ^ x[12];
  assign t[247] = t[299] ^ x[11];
  assign t[248] = t[300] ^ x[15];
  assign t[249] = t[301] ^ x[14];
  assign t[24] = t[42] & t[43];
  assign t[250] = t[302] ^ x[18];
  assign t[251] = t[303] ^ x[17];
  assign t[252] = t[304] ^ x[21];
  assign t[253] = t[305] ^ x[20];
  assign t[254] = t[306] ^ x[24];
  assign t[255] = t[307] ^ x[23];
  assign t[256] = t[308] ^ x[27];
  assign t[257] = t[309] ^ x[26];
  assign t[258] = t[310] ^ x[30];
  assign t[259] = t[311] ^ x[29];
  assign t[25] = t[165] ^ t[44];
  assign t[260] = t[312] ^ x[33];
  assign t[261] = t[313] ^ x[32];
  assign t[262] = t[314] ^ x[36];
  assign t[263] = t[315] ^ x[35];
  assign t[264] = t[316] ^ x[39];
  assign t[265] = t[317] ^ x[38];
  assign t[266] = t[318] ^ x[42];
  assign t[267] = t[319] ^ x[41];
  assign t[268] = t[320] ^ x[45];
  assign t[269] = t[321] ^ x[44];
  assign t[26] = t[45] ^ t[46];
  assign t[270] = t[322] ^ x[48];
  assign t[271] = t[323] ^ x[47];
  assign t[272] = t[324] ^ x[51];
  assign t[273] = t[325] ^ x[50];
  assign t[274] = t[326] ^ x[56];
  assign t[275] = t[327] ^ x[55];
  assign t[276] = t[328] ^ x[61];
  assign t[277] = t[329] ^ x[60];
  assign t[278] = t[330] ^ x[66];
  assign t[279] = t[331] ^ x[65];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[332] ^ x[73];
  assign t[281] = t[333] ^ x[72];
  assign t[282] = t[334] ^ x[76];
  assign t[283] = t[335] ^ x[75];
  assign t[284] = t[336] ^ x[81];
  assign t[285] = t[337] ^ x[80];
  assign t[286] = t[338] ^ x[86];
  assign t[287] = t[339] ^ x[85];
  assign t[288] = t[340] ^ x[91];
  assign t[289] = t[341] ^ x[90];
  assign t[28] = ~(t[49]);
  assign t[290] = t[342] ^ x[94];
  assign t[291] = t[343] ^ x[93];
  assign t[292] = t[344] ^ x[103];
  assign t[293] = t[345] ^ x[102];
  assign t[294] = (x[2]);
  assign t[295] = (x[2]);
  assign t[296] = (x[7]);
  assign t[297] = (x[7]);
  assign t[298] = (x[10]);
  assign t[299] = (x[10]);
  assign t[29] = ~(t[166]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[13]);
  assign t[301] = (x[13]);
  assign t[302] = (x[16]);
  assign t[303] = (x[16]);
  assign t[304] = (x[19]);
  assign t[305] = (x[19]);
  assign t[306] = (x[22]);
  assign t[307] = (x[22]);
  assign t[308] = (x[25]);
  assign t[309] = (x[25]);
  assign t[30] = ~(t[167]);
  assign t[310] = (x[28]);
  assign t[311] = (x[28]);
  assign t[312] = (x[31]);
  assign t[313] = (x[31]);
  assign t[314] = (x[34]);
  assign t[315] = (x[34]);
  assign t[316] = (x[37]);
  assign t[317] = (x[37]);
  assign t[318] = (x[40]);
  assign t[319] = (x[40]);
  assign t[31] = ~(t[168]);
  assign t[320] = (x[43]);
  assign t[321] = (x[43]);
  assign t[322] = (x[46]);
  assign t[323] = (x[46]);
  assign t[324] = (x[49]);
  assign t[325] = (x[49]);
  assign t[326] = (x[54]);
  assign t[327] = (x[54]);
  assign t[328] = (x[59]);
  assign t[329] = (x[59]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[64]);
  assign t[331] = (x[64]);
  assign t[332] = (x[71]);
  assign t[333] = (x[71]);
  assign t[334] = (x[74]);
  assign t[335] = (x[74]);
  assign t[336] = (x[79]);
  assign t[337] = (x[79]);
  assign t[338] = (x[84]);
  assign t[339] = (x[84]);
  assign t[33] = t[52] ? t[53] : t[169];
  assign t[340] = (x[89]);
  assign t[341] = (x[89]);
  assign t[342] = (x[92]);
  assign t[343] = (x[92]);
  assign t[344] = (x[101]);
  assign t[345] = (x[101]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[56] ^ t[33];
  assign t[36] = t[57] & t[58];
  assign t[37] = t[59] ^ t[60];
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[4] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[52] ? t[65] : t[170];
  assign t[42] = ~(t[66]);
  assign t[43] = t[167] ^ t[67];
  assign t[44] = t[52] ? t[68] : t[171];
  assign t[45] = t[69] ^ t[24];
  assign t[46] = t[70] & t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[172] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = t[8] ? t[9] : t[164];
  assign t[50] = ~(t[173]);
  assign t[51] = ~(t[76] & t[165]);
  assign t[52] = ~(t[15]);
  assign t[53] = t[169] ^ t[77];
  assign t[54] = t[78] ^ t[36];
  assign t[55] = t[79] & t[80];
  assign t[56] = t[52] ? t[81] : t[174];
  assign t[57] = ~(t[82]);
  assign t[58] = t[52] ? t[83] : t[175];
  assign t[59] = t[84] ^ t[85];
  assign t[5] = ~(t[10]);
  assign t[60] = t[86] & t[87];
  assign t[61] = t[8] ? t[88] : t[176];
  assign t[62] = t[63] ^ t[89];
  assign t[63] = t[90] ^ t[91];
  assign t[64] = t[92] & t[93];
  assign t[65] = t[170] ^ t[94];
  assign t[66] = t[166] ^ t[95];
  assign t[67] = t[52] ? t[96] : t[177];
  assign t[68] = t[171] ^ t[97];
  assign t[69] = t[98] & t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[100] ^ t[45]);
  assign t[71] = t[101] ^ t[43];
  assign t[72] = ~(t[74] & t[102]);
  assign t[73] = ~(t[178] ^ t[103]);
  assign t[74] = ~(t[104] & t[105]);
  assign t[75] = ~(t[48]);
  assign t[76] = ~(t[179]);
  assign t[77] = t[106] ? x[53] : x[52];
  assign t[78] = t[107] & t[108];
  assign t[79] = ~(t[109] ^ t[54]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[110] ^ t[58];
  assign t[81] = t[174] ^ t[111];
  assign t[82] = t[52] ? t[112] : t[180];
  assign t[83] = t[175] ^ t[113];
  assign t[84] = ~t[114];
  assign t[85] = t[115];
  assign t[86] = ~(t[59] ^ t[116]);
  assign t[87] = t[117] ^ t[118];
  assign t[88] = t[176] ^ t[119];
  assign t[89] = t[120] & t[121];
  assign t[8] = ~(t[15]);
  assign t[90] = t[122] & t[123];
  assign t[91] = t[124] & t[125];
  assign t[92] = ~(t[90] ^ t[126]);
  assign t[93] = t[127] ^ t[128];
  assign t[94] = t[75] ? x[58] : x[57];
  assign t[95] = t[27] ? t[129] : t[181];
  assign t[96] = t[177] ^ t[130];
  assign t[97] = t[75] ? x[63] : x[62];
  assign t[98] = ~(t[131]);
  assign t[99] = ~(t[41]);
  assign t[9] = t[164] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind52(x, y);
 input [111:0] x;
 output y;

 wire [334:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[128] ^ t[173];
  assign t[101] = ~(t[167]);
  assign t[102] = t[129] & t[128];
  assign t[103] = t[28] ? x[76] : x[75];
  assign t[104] = ~(t[48]);
  assign t[105] = ~(t[130]);
  assign t[106] = ~(t[35]);
  assign t[107] = ~(t[36]);
  assign t[108] = t[169] ^ t[131];
  assign t[109] = t[104] ? x[78] : x[77];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[170] ^ t[132];
  assign t[111] = t[171] ^ t[133];
  assign t[112] = ~(t[118]);
  assign t[113] = ~(t[134]);
  assign t[114] = ~(t[59]);
  assign t[115] = t[135];
  assign t[116] = t[39] ^ t[134];
  assign t[117] = t[134] ^ t[60];
  assign t[118] = t[115] ^ t[59];
  assign t[119] = t[74] ? x[80] : x[79];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[172] ^ t[136];
  assign t[121] = t[137] & t[138];
  assign t[122] = t[139] & t[94];
  assign t[123] = t[163] ^ t[140];
  assign t[124] = t[53] ? t[141] : t[174];
  assign t[125] = t[4] ^ t[52];
  assign t[126] = ~(t[129] | t[128]);
  assign t[127] = ~(t[142] | t[101]);
  assign t[128] = ~(t[175]);
  assign t[129] = ~(t[173]);
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[58] ^ t[36];
  assign t[131] = t[104] ? x[88] : x[87];
  assign t[132] = t[143] ? x[90] : x[89];
  assign t[133] = t[74] ? x[92] : x[91];
  assign t[134] = ~t[144];
  assign t[135] = t[27] ? t[145] : t[176];
  assign t[136] = t[143] ? x[97] : x[96];
  assign t[137] = ~(t[146]);
  assign t[138] = ~(t[63]);
  assign t[139] = ~(t[64]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[53] ? t[147] : t[177];
  assign t[141] = t[174] ^ t[148];
  assign t[142] = ~(t[161]);
  assign t[143] = ~(t[48]);
  assign t[144] = t[27] ? t[149] : t[178];
  assign t[145] = t[176] ^ t[150];
  assign t[146] = t[94] ^ t[64];
  assign t[147] = t[177] ^ t[151];
  assign t[148] = t[143] ? x[105] : x[104];
  assign t[149] = t[178] ^ t[152];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[104] ? x[107] : x[106];
  assign t[151] = t[74] ? x[109] : x[108];
  assign t[152] = t[74] ? x[111] : x[110];
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = t[205] ^ x[4];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[9];
  assign t[181] = t[207] ^ x[12];
  assign t[182] = t[208] ^ x[15];
  assign t[183] = t[209] ^ x[18];
  assign t[184] = t[210] ^ x[21];
  assign t[185] = t[211] ^ x[24];
  assign t[186] = t[212] ^ x[27];
  assign t[187] = t[213] ^ x[30];
  assign t[188] = t[214] ^ x[33];
  assign t[189] = t[215] ^ x[36];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[39];
  assign t[191] = t[217] ^ x[42];
  assign t[192] = t[218] ^ x[45];
  assign t[193] = t[219] ^ x[50];
  assign t[194] = t[220] ^ x[53];
  assign t[195] = t[221] ^ x[62];
  assign t[196] = t[222] ^ x[65];
  assign t[197] = t[223] ^ x[68];
  assign t[198] = t[224] ^ x[71];
  assign t[199] = t[225] ^ x[74];
  assign t[19] = t[33] ^ t[25];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[83];
  assign t[201] = t[227] ^ x[86];
  assign t[202] = t[228] ^ x[95];
  assign t[203] = t[229] ^ x[100];
  assign t[204] = t[230] ^ x[103];
  assign t[205] = (t[231] & ~t[232]);
  assign t[206] = (t[233] & ~t[234]);
  assign t[207] = (t[235] & ~t[236]);
  assign t[208] = (t[237] & ~t[238]);
  assign t[209] = (t[239] & ~t[240]);
  assign t[20] = t[34] & t[4];
  assign t[210] = (t[241] & ~t[242]);
  assign t[211] = (t[243] & ~t[244]);
  assign t[212] = (t[245] & ~t[246]);
  assign t[213] = (t[247] & ~t[248]);
  assign t[214] = (t[249] & ~t[250]);
  assign t[215] = (t[251] & ~t[252]);
  assign t[216] = (t[253] & ~t[254]);
  assign t[217] = (t[255] & ~t[256]);
  assign t[218] = (t[257] & ~t[258]);
  assign t[219] = (t[259] & ~t[260]);
  assign t[21] = t[35] ^ t[36];
  assign t[220] = (t[261] & ~t[262]);
  assign t[221] = (t[263] & ~t[264]);
  assign t[222] = (t[265] & ~t[266]);
  assign t[223] = (t[267] & ~t[268]);
  assign t[224] = (t[269] & ~t[270]);
  assign t[225] = (t[271] & ~t[272]);
  assign t[226] = (t[273] & ~t[274]);
  assign t[227] = (t[275] & ~t[276]);
  assign t[228] = (t[277] & ~t[278]);
  assign t[229] = (t[279] & ~t[280]);
  assign t[22] = t[37] & t[38];
  assign t[230] = (t[281] & ~t[282]);
  assign t[231] = t[283] ^ x[4];
  assign t[232] = t[284] ^ x[3];
  assign t[233] = t[285] ^ x[9];
  assign t[234] = t[286] ^ x[8];
  assign t[235] = t[287] ^ x[12];
  assign t[236] = t[288] ^ x[11];
  assign t[237] = t[289] ^ x[15];
  assign t[238] = t[290] ^ x[14];
  assign t[239] = t[291] ^ x[18];
  assign t[23] = t[39] ^ t[40];
  assign t[240] = t[292] ^ x[17];
  assign t[241] = t[293] ^ x[21];
  assign t[242] = t[294] ^ x[20];
  assign t[243] = t[295] ^ x[24];
  assign t[244] = t[296] ^ x[23];
  assign t[245] = t[297] ^ x[27];
  assign t[246] = t[298] ^ x[26];
  assign t[247] = t[299] ^ x[30];
  assign t[248] = t[300] ^ x[29];
  assign t[249] = t[301] ^ x[33];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[302] ^ x[32];
  assign t[251] = t[303] ^ x[36];
  assign t[252] = t[304] ^ x[35];
  assign t[253] = t[305] ^ x[39];
  assign t[254] = t[306] ^ x[38];
  assign t[255] = t[307] ^ x[42];
  assign t[256] = t[308] ^ x[41];
  assign t[257] = t[309] ^ x[45];
  assign t[258] = t[310] ^ x[44];
  assign t[259] = t[311] ^ x[50];
  assign t[25] = t[8] ? t[43] : t[154];
  assign t[260] = t[312] ^ x[49];
  assign t[261] = t[313] ^ x[53];
  assign t[262] = t[314] ^ x[52];
  assign t[263] = t[315] ^ x[62];
  assign t[264] = t[316] ^ x[61];
  assign t[265] = t[317] ^ x[65];
  assign t[266] = t[318] ^ x[64];
  assign t[267] = t[319] ^ x[68];
  assign t[268] = t[320] ^ x[67];
  assign t[269] = t[321] ^ x[71];
  assign t[26] = t[44] ^ t[45];
  assign t[270] = t[322] ^ x[70];
  assign t[271] = t[323] ^ x[74];
  assign t[272] = t[324] ^ x[73];
  assign t[273] = t[325] ^ x[83];
  assign t[274] = t[326] ^ x[82];
  assign t[275] = t[327] ^ x[86];
  assign t[276] = t[328] ^ x[85];
  assign t[277] = t[329] ^ x[95];
  assign t[278] = t[330] ^ x[94];
  assign t[279] = t[331] ^ x[100];
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = t[332] ^ x[99];
  assign t[281] = t[333] ^ x[103];
  assign t[282] = t[334] ^ x[102];
  assign t[283] = (x[2]);
  assign t[284] = (x[2]);
  assign t[285] = (x[7]);
  assign t[286] = (x[7]);
  assign t[287] = (x[10]);
  assign t[288] = (x[10]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[48]);
  assign t[290] = (x[13]);
  assign t[291] = (x[16]);
  assign t[292] = (x[16]);
  assign t[293] = (x[19]);
  assign t[294] = (x[19]);
  assign t[295] = (x[22]);
  assign t[296] = (x[22]);
  assign t[297] = (x[25]);
  assign t[298] = (x[25]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[28]);
  assign t[301] = (x[31]);
  assign t[302] = (x[31]);
  assign t[303] = (x[34]);
  assign t[304] = (x[34]);
  assign t[305] = (x[37]);
  assign t[306] = (x[37]);
  assign t[307] = (x[40]);
  assign t[308] = (x[40]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[156]);
  assign t[310] = (x[43]);
  assign t[311] = (x[48]);
  assign t[312] = (x[48]);
  assign t[313] = (x[51]);
  assign t[314] = (x[51]);
  assign t[315] = (x[60]);
  assign t[316] = (x[60]);
  assign t[317] = (x[63]);
  assign t[318] = (x[63]);
  assign t[319] = (x[66]);
  assign t[31] = ~(t[157]);
  assign t[320] = (x[66]);
  assign t[321] = (x[69]);
  assign t[322] = (x[69]);
  assign t[323] = (x[72]);
  assign t[324] = (x[72]);
  assign t[325] = (x[81]);
  assign t[326] = (x[81]);
  assign t[327] = (x[84]);
  assign t[328] = (x[84]);
  assign t[329] = (x[93]);
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = (x[93]);
  assign t[331] = (x[98]);
  assign t[332] = (x[98]);
  assign t[333] = (x[101]);
  assign t[334] = (x[101]);
  assign t[33] = t[8] ? t[51] : t[158];
  assign t[34] = ~(t[52]);
  assign t[35] = t[53] ? t[54] : t[159];
  assign t[36] = t[53] ? t[55] : t[160];
  assign t[37] = ~(t[21] ^ t[56]);
  assign t[38] = t[57] ^ t[58];
  assign t[39] = t[59] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[154] ^ t[67];
  assign t[44] = t[68] ^ t[20];
  assign t[45] = t[69] & t[70];
  assign t[46] = ~(t[71] & t[72]);
  assign t[47] = t[161] | t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = ~(t[162]);
  assign t[4] = t[8] ? t[9] : t[153];
  assign t[50] = ~(t[75] & t[163]);
  assign t[51] = t[158] ^ t[76];
  assign t[52] = t[8] ? t[77] : t[164];
  assign t[53] = ~(t[15]);
  assign t[54] = t[159] ^ t[78];
  assign t[55] = t[160] ^ t[79];
  assign t[56] = t[80] ^ t[81];
  assign t[57] = t[36] ^ t[82];
  assign t[58] = t[53] ? t[83] : t[165];
  assign t[59] = t[84];
  assign t[5] = ~(t[10]);
  assign t[60] = ~t[85];
  assign t[61] = t[86] ^ t[87];
  assign t[62] = t[88] & t[89];
  assign t[63] = t[53] ? t[90] : t[166];
  assign t[64] = t[155] ^ t[91];
  assign t[65] = ~(t[41] ^ t[92]);
  assign t[66] = t[93] ^ t[94];
  assign t[67] = t[28] ? x[47] : x[46];
  assign t[68] = t[95] & t[96];
  assign t[69] = ~(t[97] ^ t[44]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[98] ^ t[4];
  assign t[71] = ~(t[73] & t[99]);
  assign t[72] = ~(t[167] ^ t[100]);
  assign t[73] = ~(t[101] & t[102]);
  assign t[74] = ~(t[47]);
  assign t[75] = ~(t[168]);
  assign t[76] = t[28] ? x[55] : x[54];
  assign t[77] = t[164] ^ t[103];
  assign t[78] = t[104] ? x[57] : x[56];
  assign t[79] = t[104] ? x[59] : x[58];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[105] & t[106];
  assign t[81] = t[107] & t[58];
  assign t[82] = t[53] ? t[108] : t[169];
  assign t[83] = t[165] ^ t[109];
  assign t[84] = t[27] ? t[110] : t[170];
  assign t[85] = t[27] ? t[111] : t[171];
  assign t[86] = t[112] & t[113];
  assign t[87] = t[114] & t[115];
  assign t[88] = ~(t[86] ^ t[116]);
  assign t[89] = t[117] ^ t[118];
  assign t[8] = ~(t[15]);
  assign t[90] = t[166] ^ t[119];
  assign t[91] = t[27] ? t[120] : t[172];
  assign t[92] = t[121] ^ t[122];
  assign t[93] = t[64] ^ t[123];
  assign t[94] = t[156] ^ t[124];
  assign t[95] = ~(t[125]);
  assign t[96] = ~(t[33]);
  assign t[97] = t[33] ^ t[52];
  assign t[98] = t[52] ^ t[25];
  assign t[99] = ~(t[126] & t[127]);
  assign t[9] = t[153] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind53(x, y);
 input [111:0] x;
 output y;

 wire [334:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[128] ^ t[173];
  assign t[101] = ~(t[167]);
  assign t[102] = t[129] & t[128];
  assign t[103] = t[28] ? x[76] : x[75];
  assign t[104] = ~(t[48]);
  assign t[105] = ~(t[130]);
  assign t[106] = ~(t[35]);
  assign t[107] = ~(t[36]);
  assign t[108] = t[169] ^ t[131];
  assign t[109] = t[104] ? x[78] : x[77];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[170] ^ t[132];
  assign t[111] = t[171] ^ t[133];
  assign t[112] = ~(t[118]);
  assign t[113] = ~(t[134]);
  assign t[114] = ~(t[59]);
  assign t[115] = t[135];
  assign t[116] = t[39] ^ t[134];
  assign t[117] = t[134] ^ t[60];
  assign t[118] = t[115] ^ t[59];
  assign t[119] = t[74] ? x[80] : x[79];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[172] ^ t[136];
  assign t[121] = t[137] & t[138];
  assign t[122] = t[139] & t[94];
  assign t[123] = t[163] ^ t[140];
  assign t[124] = t[53] ? t[141] : t[174];
  assign t[125] = t[4] ^ t[52];
  assign t[126] = ~(t[129] | t[128]);
  assign t[127] = ~(t[142] | t[101]);
  assign t[128] = ~(t[175]);
  assign t[129] = ~(t[173]);
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[58] ^ t[36];
  assign t[131] = t[104] ? x[88] : x[87];
  assign t[132] = t[143] ? x[90] : x[89];
  assign t[133] = t[74] ? x[92] : x[91];
  assign t[134] = ~t[144];
  assign t[135] = t[27] ? t[145] : t[176];
  assign t[136] = t[143] ? x[97] : x[96];
  assign t[137] = ~(t[146]);
  assign t[138] = ~(t[63]);
  assign t[139] = ~(t[64]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[53] ? t[147] : t[177];
  assign t[141] = t[174] ^ t[148];
  assign t[142] = ~(t[161]);
  assign t[143] = ~(t[48]);
  assign t[144] = t[27] ? t[149] : t[178];
  assign t[145] = t[176] ^ t[150];
  assign t[146] = t[94] ^ t[64];
  assign t[147] = t[177] ^ t[151];
  assign t[148] = t[143] ? x[105] : x[104];
  assign t[149] = t[178] ^ t[152];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[104] ? x[107] : x[106];
  assign t[151] = t[74] ? x[109] : x[108];
  assign t[152] = t[74] ? x[111] : x[110];
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = (t[204]);
  assign t[179] = t[205] ^ x[4];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[9];
  assign t[181] = t[207] ^ x[12];
  assign t[182] = t[208] ^ x[15];
  assign t[183] = t[209] ^ x[18];
  assign t[184] = t[210] ^ x[21];
  assign t[185] = t[211] ^ x[24];
  assign t[186] = t[212] ^ x[27];
  assign t[187] = t[213] ^ x[30];
  assign t[188] = t[214] ^ x[33];
  assign t[189] = t[215] ^ x[36];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[39];
  assign t[191] = t[217] ^ x[42];
  assign t[192] = t[218] ^ x[45];
  assign t[193] = t[219] ^ x[50];
  assign t[194] = t[220] ^ x[53];
  assign t[195] = t[221] ^ x[62];
  assign t[196] = t[222] ^ x[65];
  assign t[197] = t[223] ^ x[68];
  assign t[198] = t[224] ^ x[71];
  assign t[199] = t[225] ^ x[74];
  assign t[19] = t[33] ^ t[25];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[83];
  assign t[201] = t[227] ^ x[86];
  assign t[202] = t[228] ^ x[95];
  assign t[203] = t[229] ^ x[100];
  assign t[204] = t[230] ^ x[103];
  assign t[205] = (t[231] & ~t[232]);
  assign t[206] = (t[233] & ~t[234]);
  assign t[207] = (t[235] & ~t[236]);
  assign t[208] = (t[237] & ~t[238]);
  assign t[209] = (t[239] & ~t[240]);
  assign t[20] = t[34] & t[4];
  assign t[210] = (t[241] & ~t[242]);
  assign t[211] = (t[243] & ~t[244]);
  assign t[212] = (t[245] & ~t[246]);
  assign t[213] = (t[247] & ~t[248]);
  assign t[214] = (t[249] & ~t[250]);
  assign t[215] = (t[251] & ~t[252]);
  assign t[216] = (t[253] & ~t[254]);
  assign t[217] = (t[255] & ~t[256]);
  assign t[218] = (t[257] & ~t[258]);
  assign t[219] = (t[259] & ~t[260]);
  assign t[21] = t[35] ^ t[36];
  assign t[220] = (t[261] & ~t[262]);
  assign t[221] = (t[263] & ~t[264]);
  assign t[222] = (t[265] & ~t[266]);
  assign t[223] = (t[267] & ~t[268]);
  assign t[224] = (t[269] & ~t[270]);
  assign t[225] = (t[271] & ~t[272]);
  assign t[226] = (t[273] & ~t[274]);
  assign t[227] = (t[275] & ~t[276]);
  assign t[228] = (t[277] & ~t[278]);
  assign t[229] = (t[279] & ~t[280]);
  assign t[22] = t[37] & t[38];
  assign t[230] = (t[281] & ~t[282]);
  assign t[231] = t[283] ^ x[4];
  assign t[232] = t[284] ^ x[3];
  assign t[233] = t[285] ^ x[9];
  assign t[234] = t[286] ^ x[8];
  assign t[235] = t[287] ^ x[12];
  assign t[236] = t[288] ^ x[11];
  assign t[237] = t[289] ^ x[15];
  assign t[238] = t[290] ^ x[14];
  assign t[239] = t[291] ^ x[18];
  assign t[23] = t[39] ^ t[40];
  assign t[240] = t[292] ^ x[17];
  assign t[241] = t[293] ^ x[21];
  assign t[242] = t[294] ^ x[20];
  assign t[243] = t[295] ^ x[24];
  assign t[244] = t[296] ^ x[23];
  assign t[245] = t[297] ^ x[27];
  assign t[246] = t[298] ^ x[26];
  assign t[247] = t[299] ^ x[30];
  assign t[248] = t[300] ^ x[29];
  assign t[249] = t[301] ^ x[33];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[302] ^ x[32];
  assign t[251] = t[303] ^ x[36];
  assign t[252] = t[304] ^ x[35];
  assign t[253] = t[305] ^ x[39];
  assign t[254] = t[306] ^ x[38];
  assign t[255] = t[307] ^ x[42];
  assign t[256] = t[308] ^ x[41];
  assign t[257] = t[309] ^ x[45];
  assign t[258] = t[310] ^ x[44];
  assign t[259] = t[311] ^ x[50];
  assign t[25] = t[8] ? t[43] : t[154];
  assign t[260] = t[312] ^ x[49];
  assign t[261] = t[313] ^ x[53];
  assign t[262] = t[314] ^ x[52];
  assign t[263] = t[315] ^ x[62];
  assign t[264] = t[316] ^ x[61];
  assign t[265] = t[317] ^ x[65];
  assign t[266] = t[318] ^ x[64];
  assign t[267] = t[319] ^ x[68];
  assign t[268] = t[320] ^ x[67];
  assign t[269] = t[321] ^ x[71];
  assign t[26] = t[44] ^ t[45];
  assign t[270] = t[322] ^ x[70];
  assign t[271] = t[323] ^ x[74];
  assign t[272] = t[324] ^ x[73];
  assign t[273] = t[325] ^ x[83];
  assign t[274] = t[326] ^ x[82];
  assign t[275] = t[327] ^ x[86];
  assign t[276] = t[328] ^ x[85];
  assign t[277] = t[329] ^ x[95];
  assign t[278] = t[330] ^ x[94];
  assign t[279] = t[331] ^ x[100];
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = t[332] ^ x[99];
  assign t[281] = t[333] ^ x[103];
  assign t[282] = t[334] ^ x[102];
  assign t[283] = (x[2]);
  assign t[284] = (x[2]);
  assign t[285] = (x[7]);
  assign t[286] = (x[7]);
  assign t[287] = (x[10]);
  assign t[288] = (x[10]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[48]);
  assign t[290] = (x[13]);
  assign t[291] = (x[16]);
  assign t[292] = (x[16]);
  assign t[293] = (x[19]);
  assign t[294] = (x[19]);
  assign t[295] = (x[22]);
  assign t[296] = (x[22]);
  assign t[297] = (x[25]);
  assign t[298] = (x[25]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[28]);
  assign t[301] = (x[31]);
  assign t[302] = (x[31]);
  assign t[303] = (x[34]);
  assign t[304] = (x[34]);
  assign t[305] = (x[37]);
  assign t[306] = (x[37]);
  assign t[307] = (x[40]);
  assign t[308] = (x[40]);
  assign t[309] = (x[43]);
  assign t[30] = ~(t[156]);
  assign t[310] = (x[43]);
  assign t[311] = (x[48]);
  assign t[312] = (x[48]);
  assign t[313] = (x[51]);
  assign t[314] = (x[51]);
  assign t[315] = (x[60]);
  assign t[316] = (x[60]);
  assign t[317] = (x[63]);
  assign t[318] = (x[63]);
  assign t[319] = (x[66]);
  assign t[31] = ~(t[157]);
  assign t[320] = (x[66]);
  assign t[321] = (x[69]);
  assign t[322] = (x[69]);
  assign t[323] = (x[72]);
  assign t[324] = (x[72]);
  assign t[325] = (x[81]);
  assign t[326] = (x[81]);
  assign t[327] = (x[84]);
  assign t[328] = (x[84]);
  assign t[329] = (x[93]);
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = (x[93]);
  assign t[331] = (x[98]);
  assign t[332] = (x[98]);
  assign t[333] = (x[101]);
  assign t[334] = (x[101]);
  assign t[33] = t[8] ? t[51] : t[158];
  assign t[34] = ~(t[52]);
  assign t[35] = t[53] ? t[54] : t[159];
  assign t[36] = t[53] ? t[55] : t[160];
  assign t[37] = ~(t[21] ^ t[56]);
  assign t[38] = t[57] ^ t[58];
  assign t[39] = t[59] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] & t[66];
  assign t[43] = t[154] ^ t[67];
  assign t[44] = t[68] ^ t[20];
  assign t[45] = t[69] & t[70];
  assign t[46] = ~(t[71] & t[72]);
  assign t[47] = t[161] | t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = ~(t[162]);
  assign t[4] = t[8] ? t[9] : t[153];
  assign t[50] = ~(t[75] & t[163]);
  assign t[51] = t[158] ^ t[76];
  assign t[52] = t[8] ? t[77] : t[164];
  assign t[53] = ~(t[15]);
  assign t[54] = t[159] ^ t[78];
  assign t[55] = t[160] ^ t[79];
  assign t[56] = t[80] ^ t[81];
  assign t[57] = t[36] ^ t[82];
  assign t[58] = t[53] ? t[83] : t[165];
  assign t[59] = t[84];
  assign t[5] = ~(t[10]);
  assign t[60] = ~t[85];
  assign t[61] = t[86] ^ t[87];
  assign t[62] = t[88] & t[89];
  assign t[63] = t[53] ? t[90] : t[166];
  assign t[64] = t[155] ^ t[91];
  assign t[65] = ~(t[41] ^ t[92]);
  assign t[66] = t[93] ^ t[94];
  assign t[67] = t[28] ? x[47] : x[46];
  assign t[68] = t[95] & t[96];
  assign t[69] = ~(t[97] ^ t[44]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[98] ^ t[4];
  assign t[71] = ~(t[73] & t[99]);
  assign t[72] = ~(t[167] ^ t[100]);
  assign t[73] = ~(t[101] & t[102]);
  assign t[74] = ~(t[47]);
  assign t[75] = ~(t[168]);
  assign t[76] = t[28] ? x[55] : x[54];
  assign t[77] = t[164] ^ t[103];
  assign t[78] = t[104] ? x[57] : x[56];
  assign t[79] = t[104] ? x[59] : x[58];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[105] & t[106];
  assign t[81] = t[107] & t[58];
  assign t[82] = t[53] ? t[108] : t[169];
  assign t[83] = t[165] ^ t[109];
  assign t[84] = t[27] ? t[110] : t[170];
  assign t[85] = t[27] ? t[111] : t[171];
  assign t[86] = t[112] & t[113];
  assign t[87] = t[114] & t[115];
  assign t[88] = ~(t[86] ^ t[116]);
  assign t[89] = t[117] ^ t[118];
  assign t[8] = ~(t[15]);
  assign t[90] = t[166] ^ t[119];
  assign t[91] = t[27] ? t[120] : t[172];
  assign t[92] = t[121] ^ t[122];
  assign t[93] = t[64] ^ t[123];
  assign t[94] = t[156] ^ t[124];
  assign t[95] = ~(t[125]);
  assign t[96] = ~(t[33]);
  assign t[97] = t[33] ^ t[52];
  assign t[98] = t[52] ^ t[25];
  assign t[99] = ~(t[126] & t[127]);
  assign t[9] = t[153] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind54(x, y);
 input [111:0] x;
 output y;

 wire [333:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[167] ^ t[127];
  assign t[101] = t[168] ^ t[128];
  assign t[102] = ~(t[108]);
  assign t[103] = ~(t[129]);
  assign t[104] = ~(t[52]);
  assign t[105] = t[156] ^ t[130];
  assign t[106] = t[33] ^ t[129];
  assign t[107] = t[129] ^ t[53];
  assign t[108] = t[105] ^ t[52];
  assign t[109] = t[75] ? x[71] : x[70];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[131]);
  assign t[111] = ~(t[132]);
  assign t[112] = ~(t[133]);
  assign t[113] = t[134];
  assign t[114] = t[132] ^ t[133];
  assign t[115] = t[133] ^ t[35];
  assign t[116] = ~(t[135]);
  assign t[117] = ~(t[4]);
  assign t[118] = ~(t[37]);
  assign t[119] = t[169] ^ t[136];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[28] ? x[73] : x[72];
  assign t[121] = t[170] ^ t[137];
  assign t[122] = t[93] ? x[75] : x[74];
  assign t[123] = ~(t[126] | t[125]);
  assign t[124] = ~(t[138] | t[98]);
  assign t[125] = ~(t[172]);
  assign t[126] = ~(t[171]);
  assign t[127] = t[139] ? x[80] : x[79];
  assign t[128] = t[75] ? x[82] : x[81];
  assign t[129] = t[40] ? t[140] : t[173];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[40] ? t[141] : t[174];
  assign t[131] = t[113] ^ t[133];
  assign t[132] = ~t[142];
  assign t[133] = t[143];
  assign t[134] = t[27] ? t[144] : t[175];
  assign t[135] = t[62] ^ t[37];
  assign t[136] = t[28] ? x[93] : x[92];
  assign t[137] = t[93] ? x[95] : x[94];
  assign t[138] = ~(t[159]);
  assign t[139] = ~(t[49]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[173] ^ t[145];
  assign t[141] = t[174] ^ t[146];
  assign t[142] = t[27] ? t[147] : t[176];
  assign t[143] = t[27] ? t[148] : t[177];
  assign t[144] = t[175] ^ t[149];
  assign t[145] = t[75] ? x[103] : x[102];
  assign t[146] = t[139] ? x[105] : x[104];
  assign t[147] = t[176] ^ t[150];
  assign t[148] = t[177] ^ t[151];
  assign t[149] = t[93] ? x[107] : x[106];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[75] ? x[109] : x[108];
  assign t[151] = t[139] ? x[111] : x[110];
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = t[204] ^ x[4];
  assign t[179] = t[205] ^ x[9];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[12];
  assign t[181] = t[207] ^ x[15];
  assign t[182] = t[208] ^ x[18];
  assign t[183] = t[209] ^ x[21];
  assign t[184] = t[210] ^ x[24];
  assign t[185] = t[211] ^ x[27];
  assign t[186] = t[212] ^ x[30];
  assign t[187] = t[213] ^ x[33];
  assign t[188] = t[214] ^ x[36];
  assign t[189] = t[215] ^ x[39];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[46];
  assign t[191] = t[217] ^ x[49];
  assign t[192] = t[218] ^ x[52];
  assign t[193] = t[219] ^ x[55];
  assign t[194] = t[220] ^ x[58];
  assign t[195] = t[221] ^ x[63];
  assign t[196] = t[222] ^ x[66];
  assign t[197] = t[223] ^ x[69];
  assign t[198] = t[224] ^ x[78];
  assign t[199] = t[225] ^ x[85];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[88];
  assign t[201] = t[227] ^ x[91];
  assign t[202] = t[228] ^ x[98];
  assign t[203] = t[229] ^ x[101];
  assign t[204] = (t[230] & ~t[231]);
  assign t[205] = (t[232] & ~t[233]);
  assign t[206] = (t[234] & ~t[235]);
  assign t[207] = (t[236] & ~t[237]);
  assign t[208] = (t[238] & ~t[239]);
  assign t[209] = (t[240] & ~t[241]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[242] & ~t[243]);
  assign t[211] = (t[244] & ~t[245]);
  assign t[212] = (t[246] & ~t[247]);
  assign t[213] = (t[248] & ~t[249]);
  assign t[214] = (t[250] & ~t[251]);
  assign t[215] = (t[252] & ~t[253]);
  assign t[216] = (t[254] & ~t[255]);
  assign t[217] = (t[256] & ~t[257]);
  assign t[218] = (t[258] & ~t[259]);
  assign t[219] = (t[260] & ~t[261]);
  assign t[21] = t[4] ^ t[37];
  assign t[220] = (t[262] & ~t[263]);
  assign t[221] = (t[264] & ~t[265]);
  assign t[222] = (t[266] & ~t[267]);
  assign t[223] = (t[268] & ~t[269]);
  assign t[224] = (t[270] & ~t[271]);
  assign t[225] = (t[272] & ~t[273]);
  assign t[226] = (t[274] & ~t[275]);
  assign t[227] = (t[276] & ~t[277]);
  assign t[228] = (t[278] & ~t[279]);
  assign t[229] = (t[280] & ~t[281]);
  assign t[22] = t[38] & t[39];
  assign t[230] = t[282] ^ x[4];
  assign t[231] = t[283] ^ x[3];
  assign t[232] = t[284] ^ x[9];
  assign t[233] = t[285] ^ x[8];
  assign t[234] = t[286] ^ x[12];
  assign t[235] = t[287] ^ x[11];
  assign t[236] = t[288] ^ x[15];
  assign t[237] = t[289] ^ x[14];
  assign t[238] = t[290] ^ x[18];
  assign t[239] = t[291] ^ x[17];
  assign t[23] = t[40] ? t[41] : t[153];
  assign t[240] = t[292] ^ x[21];
  assign t[241] = t[293] ^ x[20];
  assign t[242] = t[294] ^ x[24];
  assign t[243] = t[295] ^ x[23];
  assign t[244] = t[296] ^ x[27];
  assign t[245] = t[297] ^ x[26];
  assign t[246] = t[298] ^ x[30];
  assign t[247] = t[299] ^ x[29];
  assign t[248] = t[300] ^ x[33];
  assign t[249] = t[301] ^ x[32];
  assign t[24] = t[40] ? t[42] : t[154];
  assign t[250] = t[302] ^ x[36];
  assign t[251] = t[303] ^ x[35];
  assign t[252] = t[304] ^ x[39];
  assign t[253] = t[305] ^ x[38];
  assign t[254] = t[306] ^ x[46];
  assign t[255] = t[307] ^ x[45];
  assign t[256] = t[308] ^ x[49];
  assign t[257] = t[309] ^ x[48];
  assign t[258] = t[310] ^ x[52];
  assign t[259] = t[311] ^ x[51];
  assign t[25] = t[43] ^ t[44];
  assign t[260] = t[312] ^ x[55];
  assign t[261] = t[313] ^ x[54];
  assign t[262] = t[314] ^ x[58];
  assign t[263] = t[315] ^ x[57];
  assign t[264] = t[316] ^ x[63];
  assign t[265] = t[317] ^ x[62];
  assign t[266] = t[318] ^ x[66];
  assign t[267] = t[319] ^ x[65];
  assign t[268] = t[320] ^ x[69];
  assign t[269] = t[321] ^ x[68];
  assign t[26] = t[45] & t[46];
  assign t[270] = t[322] ^ x[78];
  assign t[271] = t[323] ^ x[77];
  assign t[272] = t[324] ^ x[85];
  assign t[273] = t[325] ^ x[84];
  assign t[274] = t[326] ^ x[88];
  assign t[275] = t[327] ^ x[87];
  assign t[276] = t[328] ^ x[91];
  assign t[277] = t[329] ^ x[90];
  assign t[278] = t[330] ^ x[98];
  assign t[279] = t[331] ^ x[97];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[332] ^ x[101];
  assign t[281] = t[333] ^ x[100];
  assign t[282] = (x[2]);
  assign t[283] = (x[2]);
  assign t[284] = (x[7]);
  assign t[285] = (x[7]);
  assign t[286] = (x[10]);
  assign t[287] = (x[10]);
  assign t[288] = (x[13]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[49]);
  assign t[290] = (x[16]);
  assign t[291] = (x[16]);
  assign t[292] = (x[19]);
  assign t[293] = (x[19]);
  assign t[294] = (x[22]);
  assign t[295] = (x[22]);
  assign t[296] = (x[25]);
  assign t[297] = (x[25]);
  assign t[298] = (x[28]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[31]);
  assign t[301] = (x[31]);
  assign t[302] = (x[34]);
  assign t[303] = (x[34]);
  assign t[304] = (x[37]);
  assign t[305] = (x[37]);
  assign t[306] = (x[44]);
  assign t[307] = (x[44]);
  assign t[308] = (x[47]);
  assign t[309] = (x[47]);
  assign t[30] = ~(t[156]);
  assign t[310] = (x[50]);
  assign t[311] = (x[50]);
  assign t[312] = (x[53]);
  assign t[313] = (x[53]);
  assign t[314] = (x[56]);
  assign t[315] = (x[56]);
  assign t[316] = (x[61]);
  assign t[317] = (x[61]);
  assign t[318] = (x[64]);
  assign t[319] = (x[64]);
  assign t[31] = ~(t[157]);
  assign t[320] = (x[67]);
  assign t[321] = (x[67]);
  assign t[322] = (x[76]);
  assign t[323] = (x[76]);
  assign t[324] = (x[83]);
  assign t[325] = (x[83]);
  assign t[326] = (x[86]);
  assign t[327] = (x[86]);
  assign t[328] = (x[89]);
  assign t[329] = (x[89]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[96]);
  assign t[331] = (x[96]);
  assign t[332] = (x[99]);
  assign t[333] = (x[99]);
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[54] ^ t[55];
  assign t[35] = ~t[56];
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[8] ? t[59] : t[158];
  assign t[38] = ~(t[21] ^ t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[15]);
  assign t[41] = t[153] ^ t[63];
  assign t[42] = t[154] ^ t[64];
  assign t[43] = t[65] & t[66];
  assign t[44] = t[67] & t[68];
  assign t[45] = ~(t[43] ^ t[69]);
  assign t[46] = t[70] ^ t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[159] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = t[8] ? t[9] : t[152];
  assign t[50] = ~(t[160]);
  assign t[51] = ~(t[76] & t[161]);
  assign t[52] = t[155] ^ t[77];
  assign t[53] = t[161] ^ t[78];
  assign t[54] = t[79] ^ t[80];
  assign t[55] = t[81] & t[82];
  assign t[56] = t[27] ? t[83] : t[162];
  assign t[57] = t[84] ^ t[85];
  assign t[58] = t[86] & t[87];
  assign t[59] = t[158] ^ t[88];
  assign t[5] = ~(t[10]);
  assign t[60] = t[89] ^ t[90];
  assign t[61] = t[37] ^ t[91];
  assign t[62] = t[8] ? t[92] : t[163];
  assign t[63] = t[93] ? x[41] : x[40];
  assign t[64] = t[93] ? x[43] : x[42];
  assign t[65] = ~(t[71]);
  assign t[66] = ~(t[94]);
  assign t[67] = ~(t[23]);
  assign t[68] = t[40] ? t[95] : t[164];
  assign t[69] = t[13] ^ t[94];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[94] ^ t[24];
  assign t[71] = t[68] ^ t[23];
  assign t[72] = ~(t[74] & t[96]);
  assign t[73] = ~(t[165] ^ t[97]);
  assign t[74] = ~(t[98] & t[99]);
  assign t[75] = ~(t[48]);
  assign t[76] = ~(t[166]);
  assign t[77] = t[27] ? t[100] : t[167];
  assign t[78] = t[40] ? t[101] : t[168];
  assign t[79] = t[102] & t[103];
  assign t[7] = t[13] ^ t[14];
  assign t[80] = t[104] & t[105];
  assign t[81] = ~(t[79] ^ t[106]);
  assign t[82] = t[107] ^ t[108];
  assign t[83] = t[162] ^ t[109];
  assign t[84] = t[110] & t[111];
  assign t[85] = t[112] & t[113];
  assign t[86] = ~(t[114] ^ t[57]);
  assign t[87] = t[115] ^ t[113];
  assign t[88] = t[28] ? x[60] : x[59];
  assign t[89] = t[116] & t[117];
  assign t[8] = ~(t[15]);
  assign t[90] = t[118] & t[62];
  assign t[91] = t[8] ? t[119] : t[169];
  assign t[92] = t[163] ^ t[120];
  assign t[93] = ~(t[49]);
  assign t[94] = t[40] ? t[121] : t[170];
  assign t[95] = t[164] ^ t[122];
  assign t[96] = ~(t[123] & t[124]);
  assign t[97] = t[125] ^ t[171];
  assign t[98] = ~(t[165]);
  assign t[99] = t[126] & t[125];
  assign t[9] = t[152] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [111:0] x;
 output y;

 wire [333:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[167] ^ t[127];
  assign t[101] = t[168] ^ t[128];
  assign t[102] = ~(t[108]);
  assign t[103] = ~(t[129]);
  assign t[104] = ~(t[52]);
  assign t[105] = t[156] ^ t[130];
  assign t[106] = t[33] ^ t[129];
  assign t[107] = t[129] ^ t[53];
  assign t[108] = t[105] ^ t[52];
  assign t[109] = t[75] ? x[71] : x[70];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[131]);
  assign t[111] = ~(t[132]);
  assign t[112] = ~(t[133]);
  assign t[113] = t[134];
  assign t[114] = t[132] ^ t[133];
  assign t[115] = t[133] ^ t[35];
  assign t[116] = ~(t[135]);
  assign t[117] = ~(t[4]);
  assign t[118] = ~(t[37]);
  assign t[119] = t[169] ^ t[136];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[28] ? x[73] : x[72];
  assign t[121] = t[170] ^ t[137];
  assign t[122] = t[93] ? x[75] : x[74];
  assign t[123] = ~(t[126] | t[125]);
  assign t[124] = ~(t[138] | t[98]);
  assign t[125] = ~(t[172]);
  assign t[126] = ~(t[171]);
  assign t[127] = t[139] ? x[80] : x[79];
  assign t[128] = t[75] ? x[82] : x[81];
  assign t[129] = t[40] ? t[140] : t[173];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[40] ? t[141] : t[174];
  assign t[131] = t[113] ^ t[133];
  assign t[132] = ~t[142];
  assign t[133] = t[143];
  assign t[134] = t[27] ? t[144] : t[175];
  assign t[135] = t[62] ^ t[37];
  assign t[136] = t[28] ? x[93] : x[92];
  assign t[137] = t[93] ? x[95] : x[94];
  assign t[138] = ~(t[159]);
  assign t[139] = ~(t[49]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[173] ^ t[145];
  assign t[141] = t[174] ^ t[146];
  assign t[142] = t[27] ? t[147] : t[176];
  assign t[143] = t[27] ? t[148] : t[177];
  assign t[144] = t[175] ^ t[149];
  assign t[145] = t[75] ? x[103] : x[102];
  assign t[146] = t[139] ? x[105] : x[104];
  assign t[147] = t[176] ^ t[150];
  assign t[148] = t[177] ^ t[151];
  assign t[149] = t[93] ? x[107] : x[106];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[75] ? x[109] : x[108];
  assign t[151] = t[139] ? x[111] : x[110];
  assign t[152] = (t[178]);
  assign t[153] = (t[179]);
  assign t[154] = (t[180]);
  assign t[155] = (t[181]);
  assign t[156] = (t[182]);
  assign t[157] = (t[183]);
  assign t[158] = (t[184]);
  assign t[159] = (t[185]);
  assign t[15] = ~(t[27]);
  assign t[160] = (t[186]);
  assign t[161] = (t[187]);
  assign t[162] = (t[188]);
  assign t[163] = (t[189]);
  assign t[164] = (t[190]);
  assign t[165] = (t[191]);
  assign t[166] = (t[192]);
  assign t[167] = (t[193]);
  assign t[168] = (t[194]);
  assign t[169] = (t[195]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = (t[196]);
  assign t[171] = (t[197]);
  assign t[172] = (t[198]);
  assign t[173] = (t[199]);
  assign t[174] = (t[200]);
  assign t[175] = (t[201]);
  assign t[176] = (t[202]);
  assign t[177] = (t[203]);
  assign t[178] = t[204] ^ x[4];
  assign t[179] = t[205] ^ x[9];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[206] ^ x[12];
  assign t[181] = t[207] ^ x[15];
  assign t[182] = t[208] ^ x[18];
  assign t[183] = t[209] ^ x[21];
  assign t[184] = t[210] ^ x[24];
  assign t[185] = t[211] ^ x[27];
  assign t[186] = t[212] ^ x[30];
  assign t[187] = t[213] ^ x[33];
  assign t[188] = t[214] ^ x[36];
  assign t[189] = t[215] ^ x[39];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[216] ^ x[46];
  assign t[191] = t[217] ^ x[49];
  assign t[192] = t[218] ^ x[52];
  assign t[193] = t[219] ^ x[55];
  assign t[194] = t[220] ^ x[58];
  assign t[195] = t[221] ^ x[63];
  assign t[196] = t[222] ^ x[66];
  assign t[197] = t[223] ^ x[69];
  assign t[198] = t[224] ^ x[78];
  assign t[199] = t[225] ^ x[85];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[226] ^ x[88];
  assign t[201] = t[227] ^ x[91];
  assign t[202] = t[228] ^ x[98];
  assign t[203] = t[229] ^ x[101];
  assign t[204] = (t[230] & ~t[231]);
  assign t[205] = (t[232] & ~t[233]);
  assign t[206] = (t[234] & ~t[235]);
  assign t[207] = (t[236] & ~t[237]);
  assign t[208] = (t[238] & ~t[239]);
  assign t[209] = (t[240] & ~t[241]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[242] & ~t[243]);
  assign t[211] = (t[244] & ~t[245]);
  assign t[212] = (t[246] & ~t[247]);
  assign t[213] = (t[248] & ~t[249]);
  assign t[214] = (t[250] & ~t[251]);
  assign t[215] = (t[252] & ~t[253]);
  assign t[216] = (t[254] & ~t[255]);
  assign t[217] = (t[256] & ~t[257]);
  assign t[218] = (t[258] & ~t[259]);
  assign t[219] = (t[260] & ~t[261]);
  assign t[21] = t[4] ^ t[37];
  assign t[220] = (t[262] & ~t[263]);
  assign t[221] = (t[264] & ~t[265]);
  assign t[222] = (t[266] & ~t[267]);
  assign t[223] = (t[268] & ~t[269]);
  assign t[224] = (t[270] & ~t[271]);
  assign t[225] = (t[272] & ~t[273]);
  assign t[226] = (t[274] & ~t[275]);
  assign t[227] = (t[276] & ~t[277]);
  assign t[228] = (t[278] & ~t[279]);
  assign t[229] = (t[280] & ~t[281]);
  assign t[22] = t[38] & t[39];
  assign t[230] = t[282] ^ x[4];
  assign t[231] = t[283] ^ x[3];
  assign t[232] = t[284] ^ x[9];
  assign t[233] = t[285] ^ x[8];
  assign t[234] = t[286] ^ x[12];
  assign t[235] = t[287] ^ x[11];
  assign t[236] = t[288] ^ x[15];
  assign t[237] = t[289] ^ x[14];
  assign t[238] = t[290] ^ x[18];
  assign t[239] = t[291] ^ x[17];
  assign t[23] = t[40] ? t[41] : t[153];
  assign t[240] = t[292] ^ x[21];
  assign t[241] = t[293] ^ x[20];
  assign t[242] = t[294] ^ x[24];
  assign t[243] = t[295] ^ x[23];
  assign t[244] = t[296] ^ x[27];
  assign t[245] = t[297] ^ x[26];
  assign t[246] = t[298] ^ x[30];
  assign t[247] = t[299] ^ x[29];
  assign t[248] = t[300] ^ x[33];
  assign t[249] = t[301] ^ x[32];
  assign t[24] = t[40] ? t[42] : t[154];
  assign t[250] = t[302] ^ x[36];
  assign t[251] = t[303] ^ x[35];
  assign t[252] = t[304] ^ x[39];
  assign t[253] = t[305] ^ x[38];
  assign t[254] = t[306] ^ x[46];
  assign t[255] = t[307] ^ x[45];
  assign t[256] = t[308] ^ x[49];
  assign t[257] = t[309] ^ x[48];
  assign t[258] = t[310] ^ x[52];
  assign t[259] = t[311] ^ x[51];
  assign t[25] = t[43] ^ t[44];
  assign t[260] = t[312] ^ x[55];
  assign t[261] = t[313] ^ x[54];
  assign t[262] = t[314] ^ x[58];
  assign t[263] = t[315] ^ x[57];
  assign t[264] = t[316] ^ x[63];
  assign t[265] = t[317] ^ x[62];
  assign t[266] = t[318] ^ x[66];
  assign t[267] = t[319] ^ x[65];
  assign t[268] = t[320] ^ x[69];
  assign t[269] = t[321] ^ x[68];
  assign t[26] = t[45] & t[46];
  assign t[270] = t[322] ^ x[78];
  assign t[271] = t[323] ^ x[77];
  assign t[272] = t[324] ^ x[85];
  assign t[273] = t[325] ^ x[84];
  assign t[274] = t[326] ^ x[88];
  assign t[275] = t[327] ^ x[87];
  assign t[276] = t[328] ^ x[91];
  assign t[277] = t[329] ^ x[90];
  assign t[278] = t[330] ^ x[98];
  assign t[279] = t[331] ^ x[97];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[332] ^ x[101];
  assign t[281] = t[333] ^ x[100];
  assign t[282] = (x[2]);
  assign t[283] = (x[2]);
  assign t[284] = (x[7]);
  assign t[285] = (x[7]);
  assign t[286] = (x[10]);
  assign t[287] = (x[10]);
  assign t[288] = (x[13]);
  assign t[289] = (x[13]);
  assign t[28] = ~(t[49]);
  assign t[290] = (x[16]);
  assign t[291] = (x[16]);
  assign t[292] = (x[19]);
  assign t[293] = (x[19]);
  assign t[294] = (x[22]);
  assign t[295] = (x[22]);
  assign t[296] = (x[25]);
  assign t[297] = (x[25]);
  assign t[298] = (x[28]);
  assign t[299] = (x[28]);
  assign t[29] = ~(t[155]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[31]);
  assign t[301] = (x[31]);
  assign t[302] = (x[34]);
  assign t[303] = (x[34]);
  assign t[304] = (x[37]);
  assign t[305] = (x[37]);
  assign t[306] = (x[44]);
  assign t[307] = (x[44]);
  assign t[308] = (x[47]);
  assign t[309] = (x[47]);
  assign t[30] = ~(t[156]);
  assign t[310] = (x[50]);
  assign t[311] = (x[50]);
  assign t[312] = (x[53]);
  assign t[313] = (x[53]);
  assign t[314] = (x[56]);
  assign t[315] = (x[56]);
  assign t[316] = (x[61]);
  assign t[317] = (x[61]);
  assign t[318] = (x[64]);
  assign t[319] = (x[64]);
  assign t[31] = ~(t[157]);
  assign t[320] = (x[67]);
  assign t[321] = (x[67]);
  assign t[322] = (x[76]);
  assign t[323] = (x[76]);
  assign t[324] = (x[83]);
  assign t[325] = (x[83]);
  assign t[326] = (x[86]);
  assign t[327] = (x[86]);
  assign t[328] = (x[89]);
  assign t[329] = (x[89]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[96]);
  assign t[331] = (x[96]);
  assign t[332] = (x[99]);
  assign t[333] = (x[99]);
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[54] ^ t[55];
  assign t[35] = ~t[56];
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[8] ? t[59] : t[158];
  assign t[38] = ~(t[21] ^ t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[15]);
  assign t[41] = t[153] ^ t[63];
  assign t[42] = t[154] ^ t[64];
  assign t[43] = t[65] & t[66];
  assign t[44] = t[67] & t[68];
  assign t[45] = ~(t[43] ^ t[69]);
  assign t[46] = t[70] ^ t[71];
  assign t[47] = ~(t[72] & t[73]);
  assign t[48] = t[159] | t[74];
  assign t[49] = ~(t[75]);
  assign t[4] = t[8] ? t[9] : t[152];
  assign t[50] = ~(t[160]);
  assign t[51] = ~(t[76] & t[161]);
  assign t[52] = t[155] ^ t[77];
  assign t[53] = t[161] ^ t[78];
  assign t[54] = t[79] ^ t[80];
  assign t[55] = t[81] & t[82];
  assign t[56] = t[27] ? t[83] : t[162];
  assign t[57] = t[84] ^ t[85];
  assign t[58] = t[86] & t[87];
  assign t[59] = t[158] ^ t[88];
  assign t[5] = ~(t[10]);
  assign t[60] = t[89] ^ t[90];
  assign t[61] = t[37] ^ t[91];
  assign t[62] = t[8] ? t[92] : t[163];
  assign t[63] = t[93] ? x[41] : x[40];
  assign t[64] = t[93] ? x[43] : x[42];
  assign t[65] = ~(t[71]);
  assign t[66] = ~(t[94]);
  assign t[67] = ~(t[23]);
  assign t[68] = t[40] ? t[95] : t[164];
  assign t[69] = t[13] ^ t[94];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[94] ^ t[24];
  assign t[71] = t[68] ^ t[23];
  assign t[72] = ~(t[74] & t[96]);
  assign t[73] = ~(t[165] ^ t[97]);
  assign t[74] = ~(t[98] & t[99]);
  assign t[75] = ~(t[48]);
  assign t[76] = ~(t[166]);
  assign t[77] = t[27] ? t[100] : t[167];
  assign t[78] = t[40] ? t[101] : t[168];
  assign t[79] = t[102] & t[103];
  assign t[7] = t[13] ^ t[14];
  assign t[80] = t[104] & t[105];
  assign t[81] = ~(t[79] ^ t[106]);
  assign t[82] = t[107] ^ t[108];
  assign t[83] = t[162] ^ t[109];
  assign t[84] = t[110] & t[111];
  assign t[85] = t[112] & t[113];
  assign t[86] = ~(t[114] ^ t[57]);
  assign t[87] = t[115] ^ t[113];
  assign t[88] = t[28] ? x[60] : x[59];
  assign t[89] = t[116] & t[117];
  assign t[8] = ~(t[15]);
  assign t[90] = t[118] & t[62];
  assign t[91] = t[8] ? t[119] : t[169];
  assign t[92] = t[163] ^ t[120];
  assign t[93] = ~(t[49]);
  assign t[94] = t[40] ? t[121] : t[170];
  assign t[95] = t[164] ^ t[122];
  assign t[96] = ~(t[123] & t[124]);
  assign t[97] = t[125] ^ t[171];
  assign t[98] = ~(t[165]);
  assign t[99] = t[126] & t[125];
  assign t[9] = t[152] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind56(x, y);
 input [116:0] x;
 output y;

 wire [360:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[122] ^ t[123];
  assign t[101] = t[42] ^ t[124];
  assign t[102] = ~t[125];
  assign t[103] = t[126];
  assign t[104] = ~(t[70] ^ t[127]);
  assign t[105] = t[128] ^ t[129];
  assign t[106] = t[188] ^ t[130];
  assign t[107] = ~(t[76] ^ t[131]);
  assign t[108] = t[132] ^ t[133];
  assign t[109] = ~(t[134]);
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[133]);
  assign t[111] = ~(t[135]);
  assign t[112] = ~(t[72]);
  assign t[113] = t[48] ? t[136] : t[191];
  assign t[114] = t[135] ^ t[72];
  assign t[115] = ~(t[173]);
  assign t[116] = ~(t[134]);
  assign t[117] = t[116] ? x[73] : x[72];
  assign t[118] = t[109] ? x[75] : x[74];
  assign t[119] = t[137] ? x[77] : x[76];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[8] ? t[138] : t[192];
  assign t[121] = t[8] ? t[139] : t[193];
  assign t[122] = t[140] ^ t[21];
  assign t[123] = t[141] & t[142];
  assign t[124] = t[143] & t[144];
  assign t[125] = t[8] ? t[145] : t[194];
  assign t[126] = t[8] ? t[146] : t[195];
  assign t[127] = t[147] ^ t[148];
  assign t[128] = t[103] ^ t[149];
  assign t[129] = t[150];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[109] ? x[91] : x[90];
  assign t[131] = t[46] ^ t[135];
  assign t[132] = t[135] ^ t[26];
  assign t[133] = t[113] ^ t[72];
  assign t[134] = ~(t[31]);
  assign t[135] = t[48] ? t[151] : t[196];
  assign t[136] = t[191] ^ t[152];
  assign t[137] = ~(t[134]);
  assign t[138] = t[192] ^ t[153];
  assign t[139] = t[193] ^ t[154];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[155] & t[156];
  assign t[141] = ~(t[140] ^ t[157]);
  assign t[142] = t[20] ^ t[158];
  assign t[143] = ~(t[159] ^ t[42]);
  assign t[144] = t[22] ^ t[95];
  assign t[145] = t[194] ^ t[160];
  assign t[146] = t[195] ^ t[161];
  assign t[147] = t[162] & t[163];
  assign t[148] = t[164] & t[129];
  assign t[149] = t[165];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[8] ? t[166] : t[197];
  assign t[151] = t[196] ^ t[167];
  assign t[152] = t[109] ? x[99] : x[98];
  assign t[153] = t[109] ? x[101] : x[100];
  assign t[154] = t[31] ? x[103] : x[102];
  assign t[155] = ~(t[158]);
  assign t[156] = ~(t[36]);
  assign t[157] = t[99] ^ t[36];
  assign t[158] = t[39] ^ t[60];
  assign t[159] = t[120] ^ t[40];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[31] ? x[105] : x[104];
  assign t[161] = t[137] ? x[107] : x[106];
  assign t[162] = ~(t[168]);
  assign t[163] = ~(t[102]);
  assign t[164] = ~(t[103]);
  assign t[165] = t[8] ? t[169] : t[198];
  assign t[166] = t[197] ^ t[170];
  assign t[167] = t[109] ? x[112] : x[111];
  assign t[168] = t[129] ^ t[103];
  assign t[169] = t[198] ^ t[171];
  assign t[16] = t[173] | t[30];
  assign t[170] = t[137] ? x[114] : x[113];
  assign t[171] = t[31] ? x[116] : x[115];
  assign t[172] = (t[199]);
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = t[226] ^ x[4];
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[7];
  assign t[201] = t[228] ^ x[12];
  assign t[202] = t[229] ^ x[15];
  assign t[203] = t[230] ^ x[18];
  assign t[204] = t[231] ^ x[21];
  assign t[205] = t[232] ^ x[24];
  assign t[206] = t[233] ^ x[27];
  assign t[207] = t[234] ^ x[30];
  assign t[208] = t[235] ^ x[33];
  assign t[209] = t[236] ^ x[36];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[39];
  assign t[211] = t[238] ^ x[42];
  assign t[212] = t[239] ^ x[45];
  assign t[213] = t[240] ^ x[48];
  assign t[214] = t[241] ^ x[51];
  assign t[215] = t[242] ^ x[54];
  assign t[216] = t[243] ^ x[59];
  assign t[217] = t[244] ^ x[62];
  assign t[218] = t[245] ^ x[71];
  assign t[219] = t[246] ^ x[80];
  assign t[21] = t[38] & t[39];
  assign t[220] = t[247] ^ x[83];
  assign t[221] = t[248] ^ x[86];
  assign t[222] = t[249] ^ x[89];
  assign t[223] = t[250] ^ x[94];
  assign t[224] = t[251] ^ x[97];
  assign t[225] = t[252] ^ x[110];
  assign t[226] = (t[253] & ~t[254]);
  assign t[227] = (t[255] & ~t[256]);
  assign t[228] = (t[257] & ~t[258]);
  assign t[229] = (t[259] & ~t[260]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[261] & ~t[262]);
  assign t[231] = (t[263] & ~t[264]);
  assign t[232] = (t[265] & ~t[266]);
  assign t[233] = (t[267] & ~t[268]);
  assign t[234] = (t[269] & ~t[270]);
  assign t[235] = (t[271] & ~t[272]);
  assign t[236] = (t[273] & ~t[274]);
  assign t[237] = (t[275] & ~t[276]);
  assign t[238] = (t[277] & ~t[278]);
  assign t[239] = (t[279] & ~t[280]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (t[281] & ~t[282]);
  assign t[241] = (t[283] & ~t[284]);
  assign t[242] = (t[285] & ~t[286]);
  assign t[243] = (t[287] & ~t[288]);
  assign t[244] = (t[289] & ~t[290]);
  assign t[245] = (t[291] & ~t[292]);
  assign t[246] = (t[293] & ~t[294]);
  assign t[247] = (t[295] & ~t[296]);
  assign t[248] = (t[297] & ~t[298]);
  assign t[249] = (t[299] & ~t[300]);
  assign t[24] = ~(t[44] ^ t[45]);
  assign t[250] = (t[301] & ~t[302]);
  assign t[251] = (t[303] & ~t[304]);
  assign t[252] = (t[305] & ~t[306]);
  assign t[253] = t[307] ^ x[4];
  assign t[254] = t[308] ^ x[3];
  assign t[255] = t[309] ^ x[7];
  assign t[256] = t[310] ^ x[6];
  assign t[257] = t[311] ^ x[12];
  assign t[258] = t[312] ^ x[11];
  assign t[259] = t[313] ^ x[15];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[314] ^ x[14];
  assign t[261] = t[315] ^ x[18];
  assign t[262] = t[316] ^ x[17];
  assign t[263] = t[317] ^ x[21];
  assign t[264] = t[318] ^ x[20];
  assign t[265] = t[319] ^ x[24];
  assign t[266] = t[320] ^ x[23];
  assign t[267] = t[321] ^ x[27];
  assign t[268] = t[322] ^ x[26];
  assign t[269] = t[323] ^ x[30];
  assign t[26] = t[48] ? t[49] : t[174];
  assign t[270] = t[324] ^ x[29];
  assign t[271] = t[325] ^ x[33];
  assign t[272] = t[326] ^ x[32];
  assign t[273] = t[327] ^ x[36];
  assign t[274] = t[328] ^ x[35];
  assign t[275] = t[329] ^ x[39];
  assign t[276] = t[330] ^ x[38];
  assign t[277] = t[331] ^ x[42];
  assign t[278] = t[332] ^ x[41];
  assign t[279] = t[333] ^ x[45];
  assign t[27] = t[50] ^ t[51];
  assign t[280] = t[334] ^ x[44];
  assign t[281] = t[335] ^ x[48];
  assign t[282] = t[336] ^ x[47];
  assign t[283] = t[337] ^ x[51];
  assign t[284] = t[338] ^ x[50];
  assign t[285] = t[339] ^ x[54];
  assign t[286] = t[340] ^ x[53];
  assign t[287] = t[341] ^ x[59];
  assign t[288] = t[342] ^ x[58];
  assign t[289] = t[343] ^ x[62];
  assign t[28] = ~(t[30] & t[52]);
  assign t[290] = t[344] ^ x[61];
  assign t[291] = t[345] ^ x[71];
  assign t[292] = t[346] ^ x[70];
  assign t[293] = t[347] ^ x[80];
  assign t[294] = t[348] ^ x[79];
  assign t[295] = t[349] ^ x[83];
  assign t[296] = t[350] ^ x[82];
  assign t[297] = t[351] ^ x[86];
  assign t[298] = t[352] ^ x[85];
  assign t[299] = t[353] ^ x[89];
  assign t[29] = ~(t[175] ^ t[53]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[88];
  assign t[301] = t[355] ^ x[94];
  assign t[302] = t[356] ^ x[93];
  assign t[303] = t[357] ^ x[97];
  assign t[304] = t[358] ^ x[96];
  assign t[305] = t[359] ^ x[110];
  assign t[306] = t[360] ^ x[109];
  assign t[307] = (x[2]);
  assign t[308] = (x[2]);
  assign t[309] = (x[5]);
  assign t[30] = ~(t[54] & t[55]);
  assign t[310] = (x[5]);
  assign t[311] = (x[10]);
  assign t[312] = (x[10]);
  assign t[313] = (x[13]);
  assign t[314] = (x[13]);
  assign t[315] = (x[16]);
  assign t[316] = (x[16]);
  assign t[317] = (x[19]);
  assign t[318] = (x[19]);
  assign t[319] = (x[22]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[22]);
  assign t[321] = (x[25]);
  assign t[322] = (x[25]);
  assign t[323] = (x[28]);
  assign t[324] = (x[28]);
  assign t[325] = (x[31]);
  assign t[326] = (x[31]);
  assign t[327] = (x[34]);
  assign t[328] = (x[34]);
  assign t[329] = (x[37]);
  assign t[32] = ~(t[176]);
  assign t[330] = (x[37]);
  assign t[331] = (x[40]);
  assign t[332] = (x[40]);
  assign t[333] = (x[43]);
  assign t[334] = (x[43]);
  assign t[335] = (x[46]);
  assign t[336] = (x[46]);
  assign t[337] = (x[49]);
  assign t[338] = (x[49]);
  assign t[339] = (x[52]);
  assign t[33] = ~(t[177]);
  assign t[340] = (x[52]);
  assign t[341] = (x[57]);
  assign t[342] = (x[57]);
  assign t[343] = (x[60]);
  assign t[344] = (x[60]);
  assign t[345] = (x[69]);
  assign t[346] = (x[69]);
  assign t[347] = (x[78]);
  assign t[348] = (x[78]);
  assign t[349] = (x[81]);
  assign t[34] = ~(t[178]);
  assign t[350] = (x[81]);
  assign t[351] = (x[84]);
  assign t[352] = (x[84]);
  assign t[353] = (x[87]);
  assign t[354] = (x[87]);
  assign t[355] = (x[92]);
  assign t[356] = (x[92]);
  assign t[357] = (x[95]);
  assign t[358] = (x[95]);
  assign t[359] = (x[108]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = (x[108]);
  assign t[36] = t[48] ? t[58] : t[179];
  assign t[37] = t[48] ? t[59] : t[180];
  assign t[38] = ~(t[60]);
  assign t[39] = t[48] ? t[61] : t[181];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[178] ^ t[62];
  assign t[41] = t[182] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] ^ t[26];
  assign t[47] = t[50] ^ t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = t[174] ^ t[75];
  assign t[4] = t[8] ? t[9] : t[172];
  assign t[50] = t[76] ^ t[77];
  assign t[51] = t[78] & t[79];
  assign t[52] = ~(t[80] & t[81]);
  assign t[53] = t[82] ^ t[183];
  assign t[54] = ~(t[175]);
  assign t[55] = t[83] & t[82];
  assign t[56] = ~(t[182]);
  assign t[57] = ~(t[84] & t[184]);
  assign t[58] = t[179] ^ t[85];
  assign t[59] = t[180] ^ t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[48] ? t[87] : t[185];
  assign t[61] = t[181] ^ t[88];
  assign t[62] = t[8] ? t[89] : t[186];
  assign t[63] = t[90] ? t[91] : t[187];
  assign t[64] = t[92] & t[93];
  assign t[65] = t[94] & t[95];
  assign t[66] = ~(t[64] ^ t[96]);
  assign t[67] = t[97] ^ t[98];
  assign t[68] = t[99] ^ t[100];
  assign t[69] = t[41] ^ t[101];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[102] ^ t[103];
  assign t[71] = t[104] & t[105];
  assign t[72] = t[48] ? t[106] : t[188];
  assign t[73] = t[107] & t[108];
  assign t[74] = ~(t[8]);
  assign t[75] = t[109] ? x[56] : x[55];
  assign t[76] = t[110] & t[111];
  assign t[77] = t[112] & t[113];
  assign t[78] = ~(t[114] ^ t[50]);
  assign t[79] = t[46] ^ t[113];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[83] | t[82]);
  assign t[81] = ~(t[115] | t[54]);
  assign t[82] = ~(t[189]);
  assign t[83] = ~(t[183]);
  assign t[84] = ~(t[190]);
  assign t[85] = t[116] ? x[64] : x[63];
  assign t[86] = t[116] ? x[66] : x[65];
  assign t[87] = t[185] ^ t[117];
  assign t[88] = t[116] ? x[68] : x[67];
  assign t[89] = t[186] ^ t[118];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = ~(t[74]);
  assign t[91] = t[187] ^ t[119];
  assign t[92] = ~(t[98]);
  assign t[93] = ~(t[120]);
  assign t[94] = ~(t[40]);
  assign t[95] = t[190] ^ t[121];
  assign t[96] = t[22] ^ t[120];
  assign t[97] = t[120] ^ t[41];
  assign t[98] = t[95] ^ t[40];
  assign t[99] = t[60] ^ t[37];
  assign t[9] = t[172] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind57(x, y);
 input [116:0] x;
 output y;

 wire [360:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[122] ^ t[123];
  assign t[101] = t[42] ^ t[124];
  assign t[102] = ~t[125];
  assign t[103] = t[126];
  assign t[104] = ~(t[70] ^ t[127]);
  assign t[105] = t[128] ^ t[129];
  assign t[106] = t[188] ^ t[130];
  assign t[107] = ~(t[76] ^ t[131]);
  assign t[108] = t[132] ^ t[133];
  assign t[109] = ~(t[134]);
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[133]);
  assign t[111] = ~(t[135]);
  assign t[112] = ~(t[72]);
  assign t[113] = t[48] ? t[136] : t[191];
  assign t[114] = t[135] ^ t[72];
  assign t[115] = ~(t[173]);
  assign t[116] = ~(t[134]);
  assign t[117] = t[116] ? x[73] : x[72];
  assign t[118] = t[109] ? x[75] : x[74];
  assign t[119] = t[137] ? x[77] : x[76];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[8] ? t[138] : t[192];
  assign t[121] = t[8] ? t[139] : t[193];
  assign t[122] = t[140] ^ t[21];
  assign t[123] = t[141] & t[142];
  assign t[124] = t[143] & t[144];
  assign t[125] = t[8] ? t[145] : t[194];
  assign t[126] = t[8] ? t[146] : t[195];
  assign t[127] = t[147] ^ t[148];
  assign t[128] = t[103] ^ t[149];
  assign t[129] = t[150];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[109] ? x[91] : x[90];
  assign t[131] = t[46] ^ t[135];
  assign t[132] = t[135] ^ t[26];
  assign t[133] = t[113] ^ t[72];
  assign t[134] = ~(t[31]);
  assign t[135] = t[48] ? t[151] : t[196];
  assign t[136] = t[191] ^ t[152];
  assign t[137] = ~(t[134]);
  assign t[138] = t[192] ^ t[153];
  assign t[139] = t[193] ^ t[154];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[155] & t[156];
  assign t[141] = ~(t[140] ^ t[157]);
  assign t[142] = t[20] ^ t[158];
  assign t[143] = ~(t[159] ^ t[42]);
  assign t[144] = t[22] ^ t[95];
  assign t[145] = t[194] ^ t[160];
  assign t[146] = t[195] ^ t[161];
  assign t[147] = t[162] & t[163];
  assign t[148] = t[164] & t[129];
  assign t[149] = t[165];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[8] ? t[166] : t[197];
  assign t[151] = t[196] ^ t[167];
  assign t[152] = t[109] ? x[99] : x[98];
  assign t[153] = t[109] ? x[101] : x[100];
  assign t[154] = t[31] ? x[103] : x[102];
  assign t[155] = ~(t[158]);
  assign t[156] = ~(t[36]);
  assign t[157] = t[99] ^ t[36];
  assign t[158] = t[39] ^ t[60];
  assign t[159] = t[120] ^ t[40];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[31] ? x[105] : x[104];
  assign t[161] = t[137] ? x[107] : x[106];
  assign t[162] = ~(t[168]);
  assign t[163] = ~(t[102]);
  assign t[164] = ~(t[103]);
  assign t[165] = t[8] ? t[169] : t[198];
  assign t[166] = t[197] ^ t[170];
  assign t[167] = t[109] ? x[112] : x[111];
  assign t[168] = t[129] ^ t[103];
  assign t[169] = t[198] ^ t[171];
  assign t[16] = t[173] | t[30];
  assign t[170] = t[137] ? x[114] : x[113];
  assign t[171] = t[31] ? x[116] : x[115];
  assign t[172] = (t[199]);
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = t[226] ^ x[4];
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[7];
  assign t[201] = t[228] ^ x[12];
  assign t[202] = t[229] ^ x[15];
  assign t[203] = t[230] ^ x[18];
  assign t[204] = t[231] ^ x[21];
  assign t[205] = t[232] ^ x[24];
  assign t[206] = t[233] ^ x[27];
  assign t[207] = t[234] ^ x[30];
  assign t[208] = t[235] ^ x[33];
  assign t[209] = t[236] ^ x[36];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[39];
  assign t[211] = t[238] ^ x[42];
  assign t[212] = t[239] ^ x[45];
  assign t[213] = t[240] ^ x[48];
  assign t[214] = t[241] ^ x[51];
  assign t[215] = t[242] ^ x[54];
  assign t[216] = t[243] ^ x[59];
  assign t[217] = t[244] ^ x[62];
  assign t[218] = t[245] ^ x[71];
  assign t[219] = t[246] ^ x[80];
  assign t[21] = t[38] & t[39];
  assign t[220] = t[247] ^ x[83];
  assign t[221] = t[248] ^ x[86];
  assign t[222] = t[249] ^ x[89];
  assign t[223] = t[250] ^ x[94];
  assign t[224] = t[251] ^ x[97];
  assign t[225] = t[252] ^ x[110];
  assign t[226] = (t[253] & ~t[254]);
  assign t[227] = (t[255] & ~t[256]);
  assign t[228] = (t[257] & ~t[258]);
  assign t[229] = (t[259] & ~t[260]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[261] & ~t[262]);
  assign t[231] = (t[263] & ~t[264]);
  assign t[232] = (t[265] & ~t[266]);
  assign t[233] = (t[267] & ~t[268]);
  assign t[234] = (t[269] & ~t[270]);
  assign t[235] = (t[271] & ~t[272]);
  assign t[236] = (t[273] & ~t[274]);
  assign t[237] = (t[275] & ~t[276]);
  assign t[238] = (t[277] & ~t[278]);
  assign t[239] = (t[279] & ~t[280]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (t[281] & ~t[282]);
  assign t[241] = (t[283] & ~t[284]);
  assign t[242] = (t[285] & ~t[286]);
  assign t[243] = (t[287] & ~t[288]);
  assign t[244] = (t[289] & ~t[290]);
  assign t[245] = (t[291] & ~t[292]);
  assign t[246] = (t[293] & ~t[294]);
  assign t[247] = (t[295] & ~t[296]);
  assign t[248] = (t[297] & ~t[298]);
  assign t[249] = (t[299] & ~t[300]);
  assign t[24] = ~(t[44] ^ t[45]);
  assign t[250] = (t[301] & ~t[302]);
  assign t[251] = (t[303] & ~t[304]);
  assign t[252] = (t[305] & ~t[306]);
  assign t[253] = t[307] ^ x[4];
  assign t[254] = t[308] ^ x[3];
  assign t[255] = t[309] ^ x[7];
  assign t[256] = t[310] ^ x[6];
  assign t[257] = t[311] ^ x[12];
  assign t[258] = t[312] ^ x[11];
  assign t[259] = t[313] ^ x[15];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[314] ^ x[14];
  assign t[261] = t[315] ^ x[18];
  assign t[262] = t[316] ^ x[17];
  assign t[263] = t[317] ^ x[21];
  assign t[264] = t[318] ^ x[20];
  assign t[265] = t[319] ^ x[24];
  assign t[266] = t[320] ^ x[23];
  assign t[267] = t[321] ^ x[27];
  assign t[268] = t[322] ^ x[26];
  assign t[269] = t[323] ^ x[30];
  assign t[26] = t[48] ? t[49] : t[174];
  assign t[270] = t[324] ^ x[29];
  assign t[271] = t[325] ^ x[33];
  assign t[272] = t[326] ^ x[32];
  assign t[273] = t[327] ^ x[36];
  assign t[274] = t[328] ^ x[35];
  assign t[275] = t[329] ^ x[39];
  assign t[276] = t[330] ^ x[38];
  assign t[277] = t[331] ^ x[42];
  assign t[278] = t[332] ^ x[41];
  assign t[279] = t[333] ^ x[45];
  assign t[27] = t[50] ^ t[51];
  assign t[280] = t[334] ^ x[44];
  assign t[281] = t[335] ^ x[48];
  assign t[282] = t[336] ^ x[47];
  assign t[283] = t[337] ^ x[51];
  assign t[284] = t[338] ^ x[50];
  assign t[285] = t[339] ^ x[54];
  assign t[286] = t[340] ^ x[53];
  assign t[287] = t[341] ^ x[59];
  assign t[288] = t[342] ^ x[58];
  assign t[289] = t[343] ^ x[62];
  assign t[28] = ~(t[30] & t[52]);
  assign t[290] = t[344] ^ x[61];
  assign t[291] = t[345] ^ x[71];
  assign t[292] = t[346] ^ x[70];
  assign t[293] = t[347] ^ x[80];
  assign t[294] = t[348] ^ x[79];
  assign t[295] = t[349] ^ x[83];
  assign t[296] = t[350] ^ x[82];
  assign t[297] = t[351] ^ x[86];
  assign t[298] = t[352] ^ x[85];
  assign t[299] = t[353] ^ x[89];
  assign t[29] = ~(t[175] ^ t[53]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[88];
  assign t[301] = t[355] ^ x[94];
  assign t[302] = t[356] ^ x[93];
  assign t[303] = t[357] ^ x[97];
  assign t[304] = t[358] ^ x[96];
  assign t[305] = t[359] ^ x[110];
  assign t[306] = t[360] ^ x[109];
  assign t[307] = (x[2]);
  assign t[308] = (x[2]);
  assign t[309] = (x[5]);
  assign t[30] = ~(t[54] & t[55]);
  assign t[310] = (x[5]);
  assign t[311] = (x[10]);
  assign t[312] = (x[10]);
  assign t[313] = (x[13]);
  assign t[314] = (x[13]);
  assign t[315] = (x[16]);
  assign t[316] = (x[16]);
  assign t[317] = (x[19]);
  assign t[318] = (x[19]);
  assign t[319] = (x[22]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[22]);
  assign t[321] = (x[25]);
  assign t[322] = (x[25]);
  assign t[323] = (x[28]);
  assign t[324] = (x[28]);
  assign t[325] = (x[31]);
  assign t[326] = (x[31]);
  assign t[327] = (x[34]);
  assign t[328] = (x[34]);
  assign t[329] = (x[37]);
  assign t[32] = ~(t[176]);
  assign t[330] = (x[37]);
  assign t[331] = (x[40]);
  assign t[332] = (x[40]);
  assign t[333] = (x[43]);
  assign t[334] = (x[43]);
  assign t[335] = (x[46]);
  assign t[336] = (x[46]);
  assign t[337] = (x[49]);
  assign t[338] = (x[49]);
  assign t[339] = (x[52]);
  assign t[33] = ~(t[177]);
  assign t[340] = (x[52]);
  assign t[341] = (x[57]);
  assign t[342] = (x[57]);
  assign t[343] = (x[60]);
  assign t[344] = (x[60]);
  assign t[345] = (x[69]);
  assign t[346] = (x[69]);
  assign t[347] = (x[78]);
  assign t[348] = (x[78]);
  assign t[349] = (x[81]);
  assign t[34] = ~(t[178]);
  assign t[350] = (x[81]);
  assign t[351] = (x[84]);
  assign t[352] = (x[84]);
  assign t[353] = (x[87]);
  assign t[354] = (x[87]);
  assign t[355] = (x[92]);
  assign t[356] = (x[92]);
  assign t[357] = (x[95]);
  assign t[358] = (x[95]);
  assign t[359] = (x[108]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = (x[108]);
  assign t[36] = t[48] ? t[58] : t[179];
  assign t[37] = t[48] ? t[59] : t[180];
  assign t[38] = ~(t[60]);
  assign t[39] = t[48] ? t[61] : t[181];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[178] ^ t[62];
  assign t[41] = t[182] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] ^ t[26];
  assign t[47] = t[50] ^ t[73];
  assign t[48] = ~(t[74]);
  assign t[49] = t[174] ^ t[75];
  assign t[4] = t[8] ? t[9] : t[172];
  assign t[50] = t[76] ^ t[77];
  assign t[51] = t[78] & t[79];
  assign t[52] = ~(t[80] & t[81]);
  assign t[53] = t[82] ^ t[183];
  assign t[54] = ~(t[175]);
  assign t[55] = t[83] & t[82];
  assign t[56] = ~(t[182]);
  assign t[57] = ~(t[84] & t[184]);
  assign t[58] = t[179] ^ t[85];
  assign t[59] = t[180] ^ t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[48] ? t[87] : t[185];
  assign t[61] = t[181] ^ t[88];
  assign t[62] = t[8] ? t[89] : t[186];
  assign t[63] = t[90] ? t[91] : t[187];
  assign t[64] = t[92] & t[93];
  assign t[65] = t[94] & t[95];
  assign t[66] = ~(t[64] ^ t[96]);
  assign t[67] = t[97] ^ t[98];
  assign t[68] = t[99] ^ t[100];
  assign t[69] = t[41] ^ t[101];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[102] ^ t[103];
  assign t[71] = t[104] & t[105];
  assign t[72] = t[48] ? t[106] : t[188];
  assign t[73] = t[107] & t[108];
  assign t[74] = ~(t[8]);
  assign t[75] = t[109] ? x[56] : x[55];
  assign t[76] = t[110] & t[111];
  assign t[77] = t[112] & t[113];
  assign t[78] = ~(t[114] ^ t[50]);
  assign t[79] = t[46] ^ t[113];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[83] | t[82]);
  assign t[81] = ~(t[115] | t[54]);
  assign t[82] = ~(t[189]);
  assign t[83] = ~(t[183]);
  assign t[84] = ~(t[190]);
  assign t[85] = t[116] ? x[64] : x[63];
  assign t[86] = t[116] ? x[66] : x[65];
  assign t[87] = t[185] ^ t[117];
  assign t[88] = t[116] ? x[68] : x[67];
  assign t[89] = t[186] ^ t[118];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = ~(t[74]);
  assign t[91] = t[187] ^ t[119];
  assign t[92] = ~(t[98]);
  assign t[93] = ~(t[120]);
  assign t[94] = ~(t[40]);
  assign t[95] = t[190] ^ t[121];
  assign t[96] = t[22] ^ t[120];
  assign t[97] = t[120] ^ t[41];
  assign t[98] = t[95] ^ t[40];
  assign t[99] = t[60] ^ t[37];
  assign t[9] = t[172] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind58(x, y);
 input [116:0] x;
 output y;

 wire [381:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] & t[125];
  assign t[101] = t[36] ? t[126] : t[209];
  assign t[102] = t[36] ? t[127] : t[210];
  assign t[103] = ~(t[71] ^ t[128]);
  assign t[104] = t[129] ^ t[130];
  assign t[105] = t[129] ^ t[131];
  assign t[106] = t[132] ^ t[133];
  assign t[107] = t[134] & t[135];
  assign t[108] = t[136] & t[137];
  assign t[109] = t[133] ^ t[138];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[139] ^ t[140];
  assign t[111] = t[141] ^ t[43];
  assign t[112] = t[36] ? t[142] : t[211];
  assign t[113] = t[128] ^ t[72];
  assign t[114] = ~(t[194]);
  assign t[115] = t[42] ^ t[64];
  assign t[116] = t[86] ? x[68] : x[67];
  assign t[117] = t[143] ? x[70] : x[69];
  assign t[118] = ~(t[144]);
  assign t[119] = ~(t[141]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = ~(t[99]);
  assign t[121] = t[208] ^ t[145];
  assign t[122] = t[141] ^ t[99];
  assign t[123] = t[8] ? t[146] : t[212];
  assign t[124] = ~(t[95] ^ t[147]);
  assign t[125] = t[111] ^ t[144];
  assign t[126] = t[209] ^ t[148];
  assign t[127] = t[210] ^ t[149];
  assign t[128] = t[150] ^ t[151];
  assign t[129] = t[102] ^ t[112];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[36] ? t[152] : t[213];
  assign t[131] = t[128] ^ t[153];
  assign t[132] = ~t[154];
  assign t[133] = t[155];
  assign t[134] = ~(t[106] ^ t[139]);
  assign t[135] = t[109] ^ t[156];
  assign t[136] = ~(t[60] ^ t[157]);
  assign t[137] = t[22] ^ t[115];
  assign t[138] = t[158];
  assign t[139] = t[159] ^ t[160];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[161] & t[162];
  assign t[141] = t[8] ? t[163] : t[214];
  assign t[142] = t[211] ^ t[164];
  assign t[143] = ~(t[55]);
  assign t[144] = t[121] ^ t[99];
  assign t[145] = t[8] ? t[165] : t[215];
  assign t[146] = t[212] ^ t[166];
  assign t[147] = t[69] ^ t[141];
  assign t[148] = t[31] ? x[84] : x[83];
  assign t[149] = t[31] ? x[86] : x[85];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[167] & t[168];
  assign t[151] = t[169] & t[130];
  assign t[152] = t[213] ^ t[170];
  assign t[153] = t[171] & t[172];
  assign t[154] = t[8] ? t[173] : t[216];
  assign t[155] = t[8] ? t[174] : t[217];
  assign t[156] = t[175];
  assign t[157] = t[75] ^ t[40];
  assign t[158] = t[8] ? t[176] : t[218];
  assign t[159] = t[177] & t[178];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[179] & t[156];
  assign t[161] = ~(t[159] ^ t[180]);
  assign t[162] = t[181] ^ t[182];
  assign t[163] = t[214] ^ t[183];
  assign t[164] = t[31] ? x[97] : x[96];
  assign t[165] = t[215] ^ t[184];
  assign t[166] = t[86] ? x[99] : x[98];
  assign t[167] = ~(t[185]);
  assign t[168] = ~(t[101]);
  assign t[169] = ~(t[102]);
  assign t[16] = t[194] | t[30];
  assign t[170] = t[31] ? x[101] : x[100];
  assign t[171] = ~(t[150] ^ t[186]);
  assign t[172] = t[187] ^ t[185];
  assign t[173] = t[216] ^ t[188];
  assign t[174] = t[217] ^ t[189];
  assign t[175] = t[8] ? t[190] : t[219];
  assign t[176] = t[218] ^ t[191];
  assign t[177] = ~(t[182]);
  assign t[178] = ~(t[132]);
  assign t[179] = ~(t[133]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[109] ^ t[132];
  assign t[181] = t[132] ^ t[138];
  assign t[182] = t[156] ^ t[133];
  assign t[183] = t[86] ? x[106] : x[105];
  assign t[184] = t[84] ? x[108] : x[107];
  assign t[185] = t[130] ^ t[102];
  assign t[186] = t[129] ^ t[101];
  assign t[187] = t[101] ^ t[112];
  assign t[188] = t[84] ? x[110] : x[109];
  assign t[189] = t[143] ? x[112] : x[111];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[219] ^ t[192];
  assign t[191] = t[84] ? x[114] : x[113];
  assign t[192] = t[143] ? x[116] : x[115];
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[36] ? t[37] : t[195];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[247] ^ x[4];
  assign t[221] = t[248] ^ x[7];
  assign t[222] = t[249] ^ x[12];
  assign t[223] = t[250] ^ x[15];
  assign t[224] = t[251] ^ x[18];
  assign t[225] = t[252] ^ x[21];
  assign t[226] = t[253] ^ x[24];
  assign t[227] = t[254] ^ x[27];
  assign t[228] = t[255] ^ x[30];
  assign t[229] = t[256] ^ x[33];
  assign t[22] = t[40] ^ t[20];
  assign t[230] = t[257] ^ x[36];
  assign t[231] = t[258] ^ x[39];
  assign t[232] = t[259] ^ x[44];
  assign t[233] = t[260] ^ x[47];
  assign t[234] = t[261] ^ x[50];
  assign t[235] = t[262] ^ x[53];
  assign t[236] = t[263] ^ x[60];
  assign t[237] = t[264] ^ x[63];
  assign t[238] = t[265] ^ x[66];
  assign t[239] = t[266] ^ x[73];
  assign t[23] = t[41] & t[42];
  assign t[240] = t[267] ^ x[76];
  assign t[241] = t[268] ^ x[79];
  assign t[242] = t[269] ^ x[82];
  assign t[243] = t[270] ^ x[89];
  assign t[244] = t[271] ^ x[92];
  assign t[245] = t[272] ^ x[95];
  assign t[246] = t[273] ^ x[104];
  assign t[247] = (t[274] & ~t[275]);
  assign t[248] = (t[276] & ~t[277]);
  assign t[249] = (t[278] & ~t[279]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (t[280] & ~t[281]);
  assign t[251] = (t[282] & ~t[283]);
  assign t[252] = (t[284] & ~t[285]);
  assign t[253] = (t[286] & ~t[287]);
  assign t[254] = (t[288] & ~t[289]);
  assign t[255] = (t[290] & ~t[291]);
  assign t[256] = (t[292] & ~t[293]);
  assign t[257] = (t[294] & ~t[295]);
  assign t[258] = (t[296] & ~t[297]);
  assign t[259] = (t[298] & ~t[299]);
  assign t[25] = t[45] ^ t[46];
  assign t[260] = (t[300] & ~t[301]);
  assign t[261] = (t[302] & ~t[303]);
  assign t[262] = (t[304] & ~t[305]);
  assign t[263] = (t[306] & ~t[307]);
  assign t[264] = (t[308] & ~t[309]);
  assign t[265] = (t[310] & ~t[311]);
  assign t[266] = (t[312] & ~t[313]);
  assign t[267] = (t[314] & ~t[315]);
  assign t[268] = (t[316] & ~t[317]);
  assign t[269] = (t[318] & ~t[319]);
  assign t[26] = ~(t[47] ^ t[48]);
  assign t[270] = (t[320] & ~t[321]);
  assign t[271] = (t[322] & ~t[323]);
  assign t[272] = (t[324] & ~t[325]);
  assign t[273] = (t[326] & ~t[327]);
  assign t[274] = t[328] ^ x[4];
  assign t[275] = t[329] ^ x[3];
  assign t[276] = t[330] ^ x[7];
  assign t[277] = t[331] ^ x[6];
  assign t[278] = t[332] ^ x[12];
  assign t[279] = t[333] ^ x[11];
  assign t[27] = ~(t[49] ^ t[50]);
  assign t[280] = t[334] ^ x[15];
  assign t[281] = t[335] ^ x[14];
  assign t[282] = t[336] ^ x[18];
  assign t[283] = t[337] ^ x[17];
  assign t[284] = t[338] ^ x[21];
  assign t[285] = t[339] ^ x[20];
  assign t[286] = t[340] ^ x[24];
  assign t[287] = t[341] ^ x[23];
  assign t[288] = t[342] ^ x[27];
  assign t[289] = t[343] ^ x[26];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[30];
  assign t[291] = t[345] ^ x[29];
  assign t[292] = t[346] ^ x[33];
  assign t[293] = t[347] ^ x[32];
  assign t[294] = t[348] ^ x[36];
  assign t[295] = t[349] ^ x[35];
  assign t[296] = t[350] ^ x[39];
  assign t[297] = t[351] ^ x[38];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[43];
  assign t[29] = ~(t[196] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[47];
  assign t[301] = t[355] ^ x[46];
  assign t[302] = t[356] ^ x[50];
  assign t[303] = t[357] ^ x[49];
  assign t[304] = t[358] ^ x[53];
  assign t[305] = t[359] ^ x[52];
  assign t[306] = t[360] ^ x[60];
  assign t[307] = t[361] ^ x[59];
  assign t[308] = t[362] ^ x[63];
  assign t[309] = t[363] ^ x[62];
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = t[364] ^ x[66];
  assign t[311] = t[365] ^ x[65];
  assign t[312] = t[366] ^ x[73];
  assign t[313] = t[367] ^ x[72];
  assign t[314] = t[368] ^ x[76];
  assign t[315] = t[369] ^ x[75];
  assign t[316] = t[370] ^ x[79];
  assign t[317] = t[371] ^ x[78];
  assign t[318] = t[372] ^ x[82];
  assign t[319] = t[373] ^ x[81];
  assign t[31] = ~(t[55]);
  assign t[320] = t[374] ^ x[89];
  assign t[321] = t[375] ^ x[88];
  assign t[322] = t[376] ^ x[92];
  assign t[323] = t[377] ^ x[91];
  assign t[324] = t[378] ^ x[95];
  assign t[325] = t[379] ^ x[94];
  assign t[326] = t[380] ^ x[104];
  assign t[327] = t[381] ^ x[103];
  assign t[328] = (x[2]);
  assign t[329] = (x[2]);
  assign t[32] = ~(t[197]);
  assign t[330] = (x[5]);
  assign t[331] = (x[5]);
  assign t[332] = (x[10]);
  assign t[333] = (x[10]);
  assign t[334] = (x[13]);
  assign t[335] = (x[13]);
  assign t[336] = (x[16]);
  assign t[337] = (x[16]);
  assign t[338] = (x[19]);
  assign t[339] = (x[19]);
  assign t[33] = ~(t[198]);
  assign t[340] = (x[22]);
  assign t[341] = (x[22]);
  assign t[342] = (x[25]);
  assign t[343] = (x[25]);
  assign t[344] = (x[28]);
  assign t[345] = (x[28]);
  assign t[346] = (x[31]);
  assign t[347] = (x[31]);
  assign t[348] = (x[34]);
  assign t[349] = (x[34]);
  assign t[34] = ~(t[199]);
  assign t[350] = (x[37]);
  assign t[351] = (x[37]);
  assign t[352] = (x[42]);
  assign t[353] = (x[42]);
  assign t[354] = (x[45]);
  assign t[355] = (x[45]);
  assign t[356] = (x[48]);
  assign t[357] = (x[48]);
  assign t[358] = (x[51]);
  assign t[359] = (x[51]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = (x[58]);
  assign t[361] = (x[58]);
  assign t[362] = (x[61]);
  assign t[363] = (x[61]);
  assign t[364] = (x[64]);
  assign t[365] = (x[64]);
  assign t[366] = (x[71]);
  assign t[367] = (x[71]);
  assign t[368] = (x[74]);
  assign t[369] = (x[74]);
  assign t[36] = ~(t[58]);
  assign t[370] = (x[77]);
  assign t[371] = (x[77]);
  assign t[372] = (x[80]);
  assign t[373] = (x[80]);
  assign t[374] = (x[87]);
  assign t[375] = (x[87]);
  assign t[376] = (x[90]);
  assign t[377] = (x[90]);
  assign t[378] = (x[93]);
  assign t[379] = (x[93]);
  assign t[37] = t[195] ^ t[59];
  assign t[380] = (x[102]);
  assign t[381] = (x[102]);
  assign t[38] = t[60] ^ t[23];
  assign t[39] = t[61] & t[62];
  assign t[3] = t[6] ^ t[7];
  assign t[40] = t[36] ? t[63] : t[200];
  assign t[41] = ~(t[64]);
  assign t[42] = t[36] ? t[65] : t[201];
  assign t[43] = t[202] ^ t[66];
  assign t[44] = t[67] ^ t[68];
  assign t[45] = t[69] ^ t[70];
  assign t[46] = t[71] ^ t[72];
  assign t[47] = ~(t[73] ^ t[74]);
  assign t[48] = t[75] ^ t[76];
  assign t[49] = t[77] ^ t[78];
  assign t[4] = t[8] ? t[9] : t[193];
  assign t[50] = ~(t[11] ^ t[79]);
  assign t[51] = ~(t[80] & t[81]);
  assign t[52] = t[82] ^ t[203];
  assign t[53] = ~(t[196]);
  assign t[54] = t[83] & t[82];
  assign t[55] = ~(t[84]);
  assign t[56] = ~(t[202]);
  assign t[57] = ~(t[85] & t[204]);
  assign t[58] = ~(t[8]);
  assign t[59] = t[86] ? x[41] : x[40];
  assign t[5] = ~(t[10]);
  assign t[60] = t[87] & t[88];
  assign t[61] = ~(t[89] ^ t[38]);
  assign t[62] = t[75] ^ t[42];
  assign t[63] = t[200] ^ t[90];
  assign t[64] = t[36] ? t[91] : t[205];
  assign t[65] = t[201] ^ t[92];
  assign t[66] = t[93] ? t[94] : t[206];
  assign t[67] = t[95] ^ t[96];
  assign t[68] = t[97] & t[98];
  assign t[69] = t[99] ^ t[43];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[67] ^ t[100];
  assign t[71] = t[101] ^ t[102];
  assign t[72] = t[103] & t[104];
  assign t[73] = t[105] ^ t[24];
  assign t[74] = t[106] ^ t[107];
  assign t[75] = t[64] ^ t[20];
  assign t[76] = t[38] ^ t[108];
  assign t[77] = t[109] ^ t[110];
  assign t[78] = t[111] ^ t[96];
  assign t[79] = t[112] ^ t[113];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[83] | t[82]);
  assign t[81] = ~(t[114] | t[53]);
  assign t[82] = ~(t[207]);
  assign t[83] = ~(t[203]);
  assign t[84] = ~(t[16]);
  assign t[85] = ~(t[208]);
  assign t[86] = ~(t[55]);
  assign t[87] = ~(t[115]);
  assign t[88] = ~(t[40]);
  assign t[89] = t[40] ^ t[64];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[86] ? x[55] : x[54];
  assign t[91] = t[205] ^ t[116];
  assign t[92] = t[86] ? x[57] : x[56];
  assign t[93] = ~(t[58]);
  assign t[94] = t[206] ^ t[117];
  assign t[95] = t[118] & t[119];
  assign t[96] = t[120] & t[121];
  assign t[97] = ~(t[122] ^ t[67]);
  assign t[98] = t[69] ^ t[121];
  assign t[99] = t[199] ^ t[123];
  assign t[9] = t[193] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind59(x, y);
 input [116:0] x;
 output y;

 wire [381:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] & t[125];
  assign t[101] = t[36] ? t[126] : t[209];
  assign t[102] = t[36] ? t[127] : t[210];
  assign t[103] = ~(t[71] ^ t[128]);
  assign t[104] = t[129] ^ t[130];
  assign t[105] = t[129] ^ t[131];
  assign t[106] = t[132] ^ t[133];
  assign t[107] = t[134] & t[135];
  assign t[108] = t[136] & t[137];
  assign t[109] = t[133] ^ t[138];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[139] ^ t[140];
  assign t[111] = t[141] ^ t[43];
  assign t[112] = t[36] ? t[142] : t[211];
  assign t[113] = t[128] ^ t[72];
  assign t[114] = ~(t[194]);
  assign t[115] = t[42] ^ t[64];
  assign t[116] = t[86] ? x[68] : x[67];
  assign t[117] = t[143] ? x[70] : x[69];
  assign t[118] = ~(t[144]);
  assign t[119] = ~(t[141]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = ~(t[99]);
  assign t[121] = t[208] ^ t[145];
  assign t[122] = t[141] ^ t[99];
  assign t[123] = t[8] ? t[146] : t[212];
  assign t[124] = ~(t[95] ^ t[147]);
  assign t[125] = t[111] ^ t[144];
  assign t[126] = t[209] ^ t[148];
  assign t[127] = t[210] ^ t[149];
  assign t[128] = t[150] ^ t[151];
  assign t[129] = t[102] ^ t[112];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[36] ? t[152] : t[213];
  assign t[131] = t[128] ^ t[153];
  assign t[132] = ~t[154];
  assign t[133] = t[155];
  assign t[134] = ~(t[106] ^ t[139]);
  assign t[135] = t[109] ^ t[156];
  assign t[136] = ~(t[60] ^ t[157]);
  assign t[137] = t[22] ^ t[115];
  assign t[138] = t[158];
  assign t[139] = t[159] ^ t[160];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[161] & t[162];
  assign t[141] = t[8] ? t[163] : t[214];
  assign t[142] = t[211] ^ t[164];
  assign t[143] = ~(t[55]);
  assign t[144] = t[121] ^ t[99];
  assign t[145] = t[8] ? t[165] : t[215];
  assign t[146] = t[212] ^ t[166];
  assign t[147] = t[69] ^ t[141];
  assign t[148] = t[31] ? x[84] : x[83];
  assign t[149] = t[31] ? x[86] : x[85];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[167] & t[168];
  assign t[151] = t[169] & t[130];
  assign t[152] = t[213] ^ t[170];
  assign t[153] = t[171] & t[172];
  assign t[154] = t[8] ? t[173] : t[216];
  assign t[155] = t[8] ? t[174] : t[217];
  assign t[156] = t[175];
  assign t[157] = t[75] ^ t[40];
  assign t[158] = t[8] ? t[176] : t[218];
  assign t[159] = t[177] & t[178];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[179] & t[156];
  assign t[161] = ~(t[159] ^ t[180]);
  assign t[162] = t[181] ^ t[182];
  assign t[163] = t[214] ^ t[183];
  assign t[164] = t[31] ? x[97] : x[96];
  assign t[165] = t[215] ^ t[184];
  assign t[166] = t[86] ? x[99] : x[98];
  assign t[167] = ~(t[185]);
  assign t[168] = ~(t[101]);
  assign t[169] = ~(t[102]);
  assign t[16] = t[194] | t[30];
  assign t[170] = t[31] ? x[101] : x[100];
  assign t[171] = ~(t[150] ^ t[186]);
  assign t[172] = t[187] ^ t[185];
  assign t[173] = t[216] ^ t[188];
  assign t[174] = t[217] ^ t[189];
  assign t[175] = t[8] ? t[190] : t[219];
  assign t[176] = t[218] ^ t[191];
  assign t[177] = ~(t[182]);
  assign t[178] = ~(t[132]);
  assign t[179] = ~(t[133]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[109] ^ t[132];
  assign t[181] = t[132] ^ t[138];
  assign t[182] = t[156] ^ t[133];
  assign t[183] = t[86] ? x[106] : x[105];
  assign t[184] = t[84] ? x[108] : x[107];
  assign t[185] = t[130] ^ t[102];
  assign t[186] = t[129] ^ t[101];
  assign t[187] = t[101] ^ t[112];
  assign t[188] = t[84] ? x[110] : x[109];
  assign t[189] = t[143] ? x[112] : x[111];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[219] ^ t[192];
  assign t[191] = t[84] ? x[114] : x[113];
  assign t[192] = t[143] ? x[116] : x[115];
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[36] ? t[37] : t[195];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = t[247] ^ x[4];
  assign t[221] = t[248] ^ x[7];
  assign t[222] = t[249] ^ x[12];
  assign t[223] = t[250] ^ x[15];
  assign t[224] = t[251] ^ x[18];
  assign t[225] = t[252] ^ x[21];
  assign t[226] = t[253] ^ x[24];
  assign t[227] = t[254] ^ x[27];
  assign t[228] = t[255] ^ x[30];
  assign t[229] = t[256] ^ x[33];
  assign t[22] = t[40] ^ t[20];
  assign t[230] = t[257] ^ x[36];
  assign t[231] = t[258] ^ x[39];
  assign t[232] = t[259] ^ x[44];
  assign t[233] = t[260] ^ x[47];
  assign t[234] = t[261] ^ x[50];
  assign t[235] = t[262] ^ x[53];
  assign t[236] = t[263] ^ x[60];
  assign t[237] = t[264] ^ x[63];
  assign t[238] = t[265] ^ x[66];
  assign t[239] = t[266] ^ x[73];
  assign t[23] = t[41] & t[42];
  assign t[240] = t[267] ^ x[76];
  assign t[241] = t[268] ^ x[79];
  assign t[242] = t[269] ^ x[82];
  assign t[243] = t[270] ^ x[89];
  assign t[244] = t[271] ^ x[92];
  assign t[245] = t[272] ^ x[95];
  assign t[246] = t[273] ^ x[104];
  assign t[247] = (t[274] & ~t[275]);
  assign t[248] = (t[276] & ~t[277]);
  assign t[249] = (t[278] & ~t[279]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (t[280] & ~t[281]);
  assign t[251] = (t[282] & ~t[283]);
  assign t[252] = (t[284] & ~t[285]);
  assign t[253] = (t[286] & ~t[287]);
  assign t[254] = (t[288] & ~t[289]);
  assign t[255] = (t[290] & ~t[291]);
  assign t[256] = (t[292] & ~t[293]);
  assign t[257] = (t[294] & ~t[295]);
  assign t[258] = (t[296] & ~t[297]);
  assign t[259] = (t[298] & ~t[299]);
  assign t[25] = t[45] ^ t[46];
  assign t[260] = (t[300] & ~t[301]);
  assign t[261] = (t[302] & ~t[303]);
  assign t[262] = (t[304] & ~t[305]);
  assign t[263] = (t[306] & ~t[307]);
  assign t[264] = (t[308] & ~t[309]);
  assign t[265] = (t[310] & ~t[311]);
  assign t[266] = (t[312] & ~t[313]);
  assign t[267] = (t[314] & ~t[315]);
  assign t[268] = (t[316] & ~t[317]);
  assign t[269] = (t[318] & ~t[319]);
  assign t[26] = ~(t[47] ^ t[48]);
  assign t[270] = (t[320] & ~t[321]);
  assign t[271] = (t[322] & ~t[323]);
  assign t[272] = (t[324] & ~t[325]);
  assign t[273] = (t[326] & ~t[327]);
  assign t[274] = t[328] ^ x[4];
  assign t[275] = t[329] ^ x[3];
  assign t[276] = t[330] ^ x[7];
  assign t[277] = t[331] ^ x[6];
  assign t[278] = t[332] ^ x[12];
  assign t[279] = t[333] ^ x[11];
  assign t[27] = ~(t[49] ^ t[50]);
  assign t[280] = t[334] ^ x[15];
  assign t[281] = t[335] ^ x[14];
  assign t[282] = t[336] ^ x[18];
  assign t[283] = t[337] ^ x[17];
  assign t[284] = t[338] ^ x[21];
  assign t[285] = t[339] ^ x[20];
  assign t[286] = t[340] ^ x[24];
  assign t[287] = t[341] ^ x[23];
  assign t[288] = t[342] ^ x[27];
  assign t[289] = t[343] ^ x[26];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[30];
  assign t[291] = t[345] ^ x[29];
  assign t[292] = t[346] ^ x[33];
  assign t[293] = t[347] ^ x[32];
  assign t[294] = t[348] ^ x[36];
  assign t[295] = t[349] ^ x[35];
  assign t[296] = t[350] ^ x[39];
  assign t[297] = t[351] ^ x[38];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[43];
  assign t[29] = ~(t[196] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[47];
  assign t[301] = t[355] ^ x[46];
  assign t[302] = t[356] ^ x[50];
  assign t[303] = t[357] ^ x[49];
  assign t[304] = t[358] ^ x[53];
  assign t[305] = t[359] ^ x[52];
  assign t[306] = t[360] ^ x[60];
  assign t[307] = t[361] ^ x[59];
  assign t[308] = t[362] ^ x[63];
  assign t[309] = t[363] ^ x[62];
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = t[364] ^ x[66];
  assign t[311] = t[365] ^ x[65];
  assign t[312] = t[366] ^ x[73];
  assign t[313] = t[367] ^ x[72];
  assign t[314] = t[368] ^ x[76];
  assign t[315] = t[369] ^ x[75];
  assign t[316] = t[370] ^ x[79];
  assign t[317] = t[371] ^ x[78];
  assign t[318] = t[372] ^ x[82];
  assign t[319] = t[373] ^ x[81];
  assign t[31] = ~(t[55]);
  assign t[320] = t[374] ^ x[89];
  assign t[321] = t[375] ^ x[88];
  assign t[322] = t[376] ^ x[92];
  assign t[323] = t[377] ^ x[91];
  assign t[324] = t[378] ^ x[95];
  assign t[325] = t[379] ^ x[94];
  assign t[326] = t[380] ^ x[104];
  assign t[327] = t[381] ^ x[103];
  assign t[328] = (x[2]);
  assign t[329] = (x[2]);
  assign t[32] = ~(t[197]);
  assign t[330] = (x[5]);
  assign t[331] = (x[5]);
  assign t[332] = (x[10]);
  assign t[333] = (x[10]);
  assign t[334] = (x[13]);
  assign t[335] = (x[13]);
  assign t[336] = (x[16]);
  assign t[337] = (x[16]);
  assign t[338] = (x[19]);
  assign t[339] = (x[19]);
  assign t[33] = ~(t[198]);
  assign t[340] = (x[22]);
  assign t[341] = (x[22]);
  assign t[342] = (x[25]);
  assign t[343] = (x[25]);
  assign t[344] = (x[28]);
  assign t[345] = (x[28]);
  assign t[346] = (x[31]);
  assign t[347] = (x[31]);
  assign t[348] = (x[34]);
  assign t[349] = (x[34]);
  assign t[34] = ~(t[199]);
  assign t[350] = (x[37]);
  assign t[351] = (x[37]);
  assign t[352] = (x[42]);
  assign t[353] = (x[42]);
  assign t[354] = (x[45]);
  assign t[355] = (x[45]);
  assign t[356] = (x[48]);
  assign t[357] = (x[48]);
  assign t[358] = (x[51]);
  assign t[359] = (x[51]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = (x[58]);
  assign t[361] = (x[58]);
  assign t[362] = (x[61]);
  assign t[363] = (x[61]);
  assign t[364] = (x[64]);
  assign t[365] = (x[64]);
  assign t[366] = (x[71]);
  assign t[367] = (x[71]);
  assign t[368] = (x[74]);
  assign t[369] = (x[74]);
  assign t[36] = ~(t[58]);
  assign t[370] = (x[77]);
  assign t[371] = (x[77]);
  assign t[372] = (x[80]);
  assign t[373] = (x[80]);
  assign t[374] = (x[87]);
  assign t[375] = (x[87]);
  assign t[376] = (x[90]);
  assign t[377] = (x[90]);
  assign t[378] = (x[93]);
  assign t[379] = (x[93]);
  assign t[37] = t[195] ^ t[59];
  assign t[380] = (x[102]);
  assign t[381] = (x[102]);
  assign t[38] = t[60] ^ t[23];
  assign t[39] = t[61] & t[62];
  assign t[3] = t[6] ^ t[7];
  assign t[40] = t[36] ? t[63] : t[200];
  assign t[41] = ~(t[64]);
  assign t[42] = t[36] ? t[65] : t[201];
  assign t[43] = t[202] ^ t[66];
  assign t[44] = t[67] ^ t[68];
  assign t[45] = t[69] ^ t[70];
  assign t[46] = t[71] ^ t[72];
  assign t[47] = ~(t[73] ^ t[74]);
  assign t[48] = t[75] ^ t[76];
  assign t[49] = t[77] ^ t[78];
  assign t[4] = t[8] ? t[9] : t[193];
  assign t[50] = ~(t[11] ^ t[79]);
  assign t[51] = ~(t[80] & t[81]);
  assign t[52] = t[82] ^ t[203];
  assign t[53] = ~(t[196]);
  assign t[54] = t[83] & t[82];
  assign t[55] = ~(t[84]);
  assign t[56] = ~(t[202]);
  assign t[57] = ~(t[85] & t[204]);
  assign t[58] = ~(t[8]);
  assign t[59] = t[86] ? x[41] : x[40];
  assign t[5] = ~(t[10]);
  assign t[60] = t[87] & t[88];
  assign t[61] = ~(t[89] ^ t[38]);
  assign t[62] = t[75] ^ t[42];
  assign t[63] = t[200] ^ t[90];
  assign t[64] = t[36] ? t[91] : t[205];
  assign t[65] = t[201] ^ t[92];
  assign t[66] = t[93] ? t[94] : t[206];
  assign t[67] = t[95] ^ t[96];
  assign t[68] = t[97] & t[98];
  assign t[69] = t[99] ^ t[43];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[67] ^ t[100];
  assign t[71] = t[101] ^ t[102];
  assign t[72] = t[103] & t[104];
  assign t[73] = t[105] ^ t[24];
  assign t[74] = t[106] ^ t[107];
  assign t[75] = t[64] ^ t[20];
  assign t[76] = t[38] ^ t[108];
  assign t[77] = t[109] ^ t[110];
  assign t[78] = t[111] ^ t[96];
  assign t[79] = t[112] ^ t[113];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[83] | t[82]);
  assign t[81] = ~(t[114] | t[53]);
  assign t[82] = ~(t[207]);
  assign t[83] = ~(t[203]);
  assign t[84] = ~(t[16]);
  assign t[85] = ~(t[208]);
  assign t[86] = ~(t[55]);
  assign t[87] = ~(t[115]);
  assign t[88] = ~(t[40]);
  assign t[89] = t[40] ^ t[64];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[86] ? x[55] : x[54];
  assign t[91] = t[205] ^ t[116];
  assign t[92] = t[86] ? x[57] : x[56];
  assign t[93] = ~(t[58]);
  assign t[94] = t[206] ^ t[117];
  assign t[95] = t[118] & t[119];
  assign t[96] = t[120] & t[121];
  assign t[97] = ~(t[122] ^ t[67]);
  assign t[98] = t[69] ^ t[121];
  assign t[99] = t[199] ^ t[123];
  assign t[9] = t[193] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [116:0] x;
 output y;

 wire [370:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[31] ? x[71] : x[70];
  assign t[101] = ~(t[112]);
  assign t[102] = t[196] ^ t[131];
  assign t[103] = t[8] ? t[132] : t[204];
  assign t[104] = t[197] ^ t[133];
  assign t[105] = t[198] ^ t[134];
  assign t[106] = t[135] & t[136];
  assign t[107] = ~(t[106] ^ t[137]);
  assign t[108] = t[62] ^ t[138];
  assign t[109] = t[139] & t[140];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[120] ^ t[73]);
  assign t[111] = t[141] ^ t[43];
  assign t[112] = ~(t[8]);
  assign t[113] = t[31] ? x[76] : x[75];
  assign t[114] = t[31] ? x[78] : x[77];
  assign t[115] = t[142] & t[143];
  assign t[116] = t[199] ^ t[144];
  assign t[117] = ~(t[183]);
  assign t[118] = t[201] ^ t[145];
  assign t[119] = ~(t[48]);
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[40] ^ t[68];
  assign t[121] = t[146];
  assign t[122] = t[124] ^ t[147];
  assign t[123] = t[148];
  assign t[124] = t[149] ^ t[150];
  assign t[125] = t[151] & t[152];
  assign t[126] = t[202] ^ t[153];
  assign t[127] = t[203] ^ t[154];
  assign t[128] = t[155] ? x[80] : x[79];
  assign t[129] = ~(t[156] ^ t[71]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[44] ^ t[97];
  assign t[131] = t[157] ? x[82] : x[81];
  assign t[132] = t[204] ^ t[158];
  assign t[133] = t[85] ? x[84] : x[83];
  assign t[134] = t[155] ? x[86] : x[85];
  assign t[135] = ~(t[138]);
  assign t[136] = ~(t[95]);
  assign t[137] = t[44] ^ t[95];
  assign t[138] = t[97] ^ t[70];
  assign t[139] = ~(t[159]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[40]);
  assign t[141] = t[68] ^ t[41];
  assign t[142] = ~(t[160]);
  assign t[143] = ~(t[47]);
  assign t[144] = t[31] ? x[88] : x[87];
  assign t[145] = t[31] ? x[90] : x[89];
  assign t[146] = t[8] ? t[161] : t[205];
  assign t[147] = t[162] & t[163];
  assign t[148] = t[8] ? t[164] : t[206];
  assign t[149] = t[165] & t[166];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[167] & t[168];
  assign t[151] = ~(t[149] ^ t[169]);
  assign t[152] = t[170] ^ t[171];
  assign t[153] = t[155] ? x[98] : x[97];
  assign t[154] = t[155] ? x[100] : x[99];
  assign t[155] = ~(t[55]);
  assign t[156] = t[95] ^ t[70];
  assign t[157] = ~(t[55]);
  assign t[158] = t[31] ? x[102] : x[101];
  assign t[159] = t[43] ^ t[68];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[80] ^ t[48];
  assign t[161] = t[205] ^ t[172];
  assign t[162] = ~(t[173] ^ t[124]);
  assign t[163] = t[93] ^ t[168];
  assign t[164] = t[206] ^ t[174];
  assign t[165] = ~(t[171]);
  assign t[166] = ~(t[175]);
  assign t[167] = ~(t[123]);
  assign t[168] = t[176];
  assign t[169] = t[93] ^ t[175];
  assign t[16] = t[183] | t[30];
  assign t[170] = t[175] ^ t[121];
  assign t[171] = t[168] ^ t[123];
  assign t[172] = t[85] ? x[104] : x[103];
  assign t[173] = t[175] ^ t[123];
  assign t[174] = t[157] ? x[106] : x[105];
  assign t[175] = ~t[177];
  assign t[176] = t[8] ? t[178] : t[207];
  assign t[177] = t[8] ? t[179] : t[208];
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[208] ^ t[181];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[157] ? x[114] : x[113];
  assign t[181] = t[85] ? x[116] : x[115];
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = t[236] ^ x[4];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[7];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[60];
  assign t[228] = t[255] ^ x[63];
  assign t[229] = t[256] ^ x[66];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[69];
  assign t[231] = t[258] ^ x[74];
  assign t[232] = t[259] ^ x[93];
  assign t[233] = t[260] ^ x[96];
  assign t[234] = t[261] ^ x[109];
  assign t[235] = t[262] ^ x[112];
  assign t[236] = (t[263] & ~t[264]);
  assign t[237] = (t[265] & ~t[266]);
  assign t[238] = (t[267] & ~t[268]);
  assign t[239] = (t[269] & ~t[270]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[271] & ~t[272]);
  assign t[241] = (t[273] & ~t[274]);
  assign t[242] = (t[275] & ~t[276]);
  assign t[243] = (t[277] & ~t[278]);
  assign t[244] = (t[279] & ~t[280]);
  assign t[245] = (t[281] & ~t[282]);
  assign t[246] = (t[283] & ~t[284]);
  assign t[247] = (t[285] & ~t[286]);
  assign t[248] = (t[287] & ~t[288]);
  assign t[249] = (t[289] & ~t[290]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[291] & ~t[292]);
  assign t[251] = (t[293] & ~t[294]);
  assign t[252] = (t[295] & ~t[296]);
  assign t[253] = (t[297] & ~t[298]);
  assign t[254] = (t[299] & ~t[300]);
  assign t[255] = (t[301] & ~t[302]);
  assign t[256] = (t[303] & ~t[304]);
  assign t[257] = (t[305] & ~t[306]);
  assign t[258] = (t[307] & ~t[308]);
  assign t[259] = (t[309] & ~t[310]);
  assign t[25] = t[41] ^ t[46];
  assign t[260] = (t[311] & ~t[312]);
  assign t[261] = (t[313] & ~t[314]);
  assign t[262] = (t[315] & ~t[316]);
  assign t[263] = t[317] ^ x[4];
  assign t[264] = t[318] ^ x[3];
  assign t[265] = t[319] ^ x[7];
  assign t[266] = t[320] ^ x[6];
  assign t[267] = t[321] ^ x[12];
  assign t[268] = t[322] ^ x[11];
  assign t[269] = t[323] ^ x[15];
  assign t[26] = t[47] ^ t[48];
  assign t[270] = t[324] ^ x[14];
  assign t[271] = t[325] ^ x[18];
  assign t[272] = t[326] ^ x[17];
  assign t[273] = t[327] ^ x[21];
  assign t[274] = t[328] ^ x[20];
  assign t[275] = t[329] ^ x[24];
  assign t[276] = t[330] ^ x[23];
  assign t[277] = t[331] ^ x[27];
  assign t[278] = t[332] ^ x[26];
  assign t[279] = t[333] ^ x[30];
  assign t[27] = t[49] & t[50];
  assign t[280] = t[334] ^ x[29];
  assign t[281] = t[335] ^ x[33];
  assign t[282] = t[336] ^ x[32];
  assign t[283] = t[337] ^ x[36];
  assign t[284] = t[338] ^ x[35];
  assign t[285] = t[339] ^ x[39];
  assign t[286] = t[340] ^ x[38];
  assign t[287] = t[341] ^ x[42];
  assign t[288] = t[342] ^ x[41];
  assign t[289] = t[343] ^ x[45];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[44];
  assign t[291] = t[345] ^ x[48];
  assign t[292] = t[346] ^ x[47];
  assign t[293] = t[347] ^ x[51];
  assign t[294] = t[348] ^ x[50];
  assign t[295] = t[349] ^ x[54];
  assign t[296] = t[350] ^ x[53];
  assign t[297] = t[351] ^ x[57];
  assign t[298] = t[352] ^ x[56];
  assign t[299] = t[353] ^ x[60];
  assign t[29] = ~(t[184] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[59];
  assign t[301] = t[355] ^ x[63];
  assign t[302] = t[356] ^ x[62];
  assign t[303] = t[357] ^ x[66];
  assign t[304] = t[358] ^ x[65];
  assign t[305] = t[359] ^ x[69];
  assign t[306] = t[360] ^ x[68];
  assign t[307] = t[361] ^ x[74];
  assign t[308] = t[362] ^ x[73];
  assign t[309] = t[363] ^ x[93];
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = t[364] ^ x[92];
  assign t[311] = t[365] ^ x[96];
  assign t[312] = t[366] ^ x[95];
  assign t[313] = t[367] ^ x[109];
  assign t[314] = t[368] ^ x[108];
  assign t[315] = t[369] ^ x[112];
  assign t[316] = t[370] ^ x[111];
  assign t[317] = (x[2]);
  assign t[318] = (x[2]);
  assign t[319] = (x[5]);
  assign t[31] = ~(t[55]);
  assign t[320] = (x[5]);
  assign t[321] = (x[10]);
  assign t[322] = (x[10]);
  assign t[323] = (x[13]);
  assign t[324] = (x[13]);
  assign t[325] = (x[16]);
  assign t[326] = (x[16]);
  assign t[327] = (x[19]);
  assign t[328] = (x[19]);
  assign t[329] = (x[22]);
  assign t[32] = ~(t[185]);
  assign t[330] = (x[22]);
  assign t[331] = (x[25]);
  assign t[332] = (x[25]);
  assign t[333] = (x[28]);
  assign t[334] = (x[28]);
  assign t[335] = (x[31]);
  assign t[336] = (x[31]);
  assign t[337] = (x[34]);
  assign t[338] = (x[34]);
  assign t[339] = (x[37]);
  assign t[33] = ~(t[186]);
  assign t[340] = (x[37]);
  assign t[341] = (x[40]);
  assign t[342] = (x[40]);
  assign t[343] = (x[43]);
  assign t[344] = (x[43]);
  assign t[345] = (x[46]);
  assign t[346] = (x[46]);
  assign t[347] = (x[49]);
  assign t[348] = (x[49]);
  assign t[349] = (x[52]);
  assign t[34] = ~(t[187]);
  assign t[350] = (x[52]);
  assign t[351] = (x[55]);
  assign t[352] = (x[55]);
  assign t[353] = (x[58]);
  assign t[354] = (x[58]);
  assign t[355] = (x[61]);
  assign t[356] = (x[61]);
  assign t[357] = (x[64]);
  assign t[358] = (x[64]);
  assign t[359] = (x[67]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = (x[67]);
  assign t[361] = (x[72]);
  assign t[362] = (x[72]);
  assign t[363] = (x[91]);
  assign t[364] = (x[91]);
  assign t[365] = (x[94]);
  assign t[366] = (x[94]);
  assign t[367] = (x[107]);
  assign t[368] = (x[107]);
  assign t[369] = (x[110]);
  assign t[36] = t[58] ^ t[59];
  assign t[370] = (x[110]);
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[38] = t[62] ^ t[63];
  assign t[39] = t[64] ^ t[65];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[66] : t[188];
  assign t[41] = t[189] ^ t[67];
  assign t[42] = ~(t[68]);
  assign t[43] = t[190] ^ t[69];
  assign t[44] = t[70] ^ t[64];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = t[73] ^ t[74];
  assign t[47] = t[75] ? t[76] : t[191];
  assign t[48] = t[75] ? t[77] : t[192];
  assign t[49] = ~(t[26] ^ t[78]);
  assign t[4] = t[8] ? t[9] : t[182];
  assign t[50] = t[79] ^ t[80];
  assign t[51] = ~(t[81] & t[82]);
  assign t[52] = t[83] ^ t[193];
  assign t[53] = ~(t[184]);
  assign t[54] = t[84] & t[83];
  assign t[55] = ~(t[85]);
  assign t[56] = ~(t[189]);
  assign t[57] = ~(t[86] & t[194]);
  assign t[58] = t[87] ^ t[88];
  assign t[59] = t[89] ^ t[90];
  assign t[5] = ~(t[10]);
  assign t[60] = ~(t[91] ^ t[92]);
  assign t[61] = t[93] ^ t[94];
  assign t[62] = t[95] ^ t[64];
  assign t[63] = t[96] & t[97];
  assign t[64] = t[75] ? t[98] : t[195];
  assign t[65] = t[71] ^ t[99];
  assign t[66] = t[188] ^ t[100];
  assign t[67] = t[101] ? t[102] : t[196];
  assign t[68] = t[187] ^ t[103];
  assign t[69] = t[8] ? t[104] : t[197];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[75] ? t[105] : t[198];
  assign t[71] = t[106] ^ t[63];
  assign t[72] = t[107] & t[108];
  assign t[73] = t[109] ^ t[23];
  assign t[74] = t[110] & t[111];
  assign t[75] = ~(t[112]);
  assign t[76] = t[191] ^ t[113];
  assign t[77] = t[192] ^ t[114];
  assign t[78] = t[115] ^ t[90];
  assign t[79] = t[48] ^ t[87];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[75] ? t[116] : t[199];
  assign t[81] = ~(t[84] | t[83]);
  assign t[82] = ~(t[117] | t[53]);
  assign t[83] = ~(t[200]);
  assign t[84] = ~(t[193]);
  assign t[85] = ~(t[16]);
  assign t[86] = ~(t[190]);
  assign t[87] = t[75] ? t[118] : t[201];
  assign t[88] = t[78] ^ t[27];
  assign t[89] = t[47] ^ t[87];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[119] & t[80];
  assign t[91] = t[120] ^ t[74];
  assign t[92] = t[121] ^ t[122];
  assign t[93] = t[123] ^ t[121];
  assign t[94] = t[124] ^ t[125];
  assign t[95] = t[75] ? t[126] : t[202];
  assign t[96] = ~(t[70]);
  assign t[97] = t[75] ? t[127] : t[203];
  assign t[98] = t[195] ^ t[128];
  assign t[99] = t[129] & t[130];
  assign t[9] = t[182] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind61(x, y);
 input [116:0] x;
 output y;

 wire [370:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[31] ? x[71] : x[70];
  assign t[101] = ~(t[112]);
  assign t[102] = t[196] ^ t[131];
  assign t[103] = t[8] ? t[132] : t[204];
  assign t[104] = t[197] ^ t[133];
  assign t[105] = t[198] ^ t[134];
  assign t[106] = t[135] & t[136];
  assign t[107] = ~(t[106] ^ t[137]);
  assign t[108] = t[62] ^ t[138];
  assign t[109] = t[139] & t[140];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[120] ^ t[73]);
  assign t[111] = t[141] ^ t[43];
  assign t[112] = ~(t[8]);
  assign t[113] = t[31] ? x[76] : x[75];
  assign t[114] = t[31] ? x[78] : x[77];
  assign t[115] = t[142] & t[143];
  assign t[116] = t[199] ^ t[144];
  assign t[117] = ~(t[183]);
  assign t[118] = t[201] ^ t[145];
  assign t[119] = ~(t[48]);
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[40] ^ t[68];
  assign t[121] = t[146];
  assign t[122] = t[124] ^ t[147];
  assign t[123] = t[148];
  assign t[124] = t[149] ^ t[150];
  assign t[125] = t[151] & t[152];
  assign t[126] = t[202] ^ t[153];
  assign t[127] = t[203] ^ t[154];
  assign t[128] = t[155] ? x[80] : x[79];
  assign t[129] = ~(t[156] ^ t[71]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[44] ^ t[97];
  assign t[131] = t[157] ? x[82] : x[81];
  assign t[132] = t[204] ^ t[158];
  assign t[133] = t[85] ? x[84] : x[83];
  assign t[134] = t[155] ? x[86] : x[85];
  assign t[135] = ~(t[138]);
  assign t[136] = ~(t[95]);
  assign t[137] = t[44] ^ t[95];
  assign t[138] = t[97] ^ t[70];
  assign t[139] = ~(t[159]);
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[40]);
  assign t[141] = t[68] ^ t[41];
  assign t[142] = ~(t[160]);
  assign t[143] = ~(t[47]);
  assign t[144] = t[31] ? x[88] : x[87];
  assign t[145] = t[31] ? x[90] : x[89];
  assign t[146] = t[8] ? t[161] : t[205];
  assign t[147] = t[162] & t[163];
  assign t[148] = t[8] ? t[164] : t[206];
  assign t[149] = t[165] & t[166];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[167] & t[168];
  assign t[151] = ~(t[149] ^ t[169]);
  assign t[152] = t[170] ^ t[171];
  assign t[153] = t[155] ? x[98] : x[97];
  assign t[154] = t[155] ? x[100] : x[99];
  assign t[155] = ~(t[55]);
  assign t[156] = t[95] ^ t[70];
  assign t[157] = ~(t[55]);
  assign t[158] = t[31] ? x[102] : x[101];
  assign t[159] = t[43] ^ t[68];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[80] ^ t[48];
  assign t[161] = t[205] ^ t[172];
  assign t[162] = ~(t[173] ^ t[124]);
  assign t[163] = t[93] ^ t[168];
  assign t[164] = t[206] ^ t[174];
  assign t[165] = ~(t[171]);
  assign t[166] = ~(t[175]);
  assign t[167] = ~(t[123]);
  assign t[168] = t[176];
  assign t[169] = t[93] ^ t[175];
  assign t[16] = t[183] | t[30];
  assign t[170] = t[175] ^ t[121];
  assign t[171] = t[168] ^ t[123];
  assign t[172] = t[85] ? x[104] : x[103];
  assign t[173] = t[175] ^ t[123];
  assign t[174] = t[157] ? x[106] : x[105];
  assign t[175] = ~t[177];
  assign t[176] = t[8] ? t[178] : t[207];
  assign t[177] = t[8] ? t[179] : t[208];
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[208] ^ t[181];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[157] ? x[114] : x[113];
  assign t[181] = t[85] ? x[116] : x[115];
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = t[236] ^ x[4];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[7];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[60];
  assign t[228] = t[255] ^ x[63];
  assign t[229] = t[256] ^ x[66];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[69];
  assign t[231] = t[258] ^ x[74];
  assign t[232] = t[259] ^ x[93];
  assign t[233] = t[260] ^ x[96];
  assign t[234] = t[261] ^ x[109];
  assign t[235] = t[262] ^ x[112];
  assign t[236] = (t[263] & ~t[264]);
  assign t[237] = (t[265] & ~t[266]);
  assign t[238] = (t[267] & ~t[268]);
  assign t[239] = (t[269] & ~t[270]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[271] & ~t[272]);
  assign t[241] = (t[273] & ~t[274]);
  assign t[242] = (t[275] & ~t[276]);
  assign t[243] = (t[277] & ~t[278]);
  assign t[244] = (t[279] & ~t[280]);
  assign t[245] = (t[281] & ~t[282]);
  assign t[246] = (t[283] & ~t[284]);
  assign t[247] = (t[285] & ~t[286]);
  assign t[248] = (t[287] & ~t[288]);
  assign t[249] = (t[289] & ~t[290]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[291] & ~t[292]);
  assign t[251] = (t[293] & ~t[294]);
  assign t[252] = (t[295] & ~t[296]);
  assign t[253] = (t[297] & ~t[298]);
  assign t[254] = (t[299] & ~t[300]);
  assign t[255] = (t[301] & ~t[302]);
  assign t[256] = (t[303] & ~t[304]);
  assign t[257] = (t[305] & ~t[306]);
  assign t[258] = (t[307] & ~t[308]);
  assign t[259] = (t[309] & ~t[310]);
  assign t[25] = t[41] ^ t[46];
  assign t[260] = (t[311] & ~t[312]);
  assign t[261] = (t[313] & ~t[314]);
  assign t[262] = (t[315] & ~t[316]);
  assign t[263] = t[317] ^ x[4];
  assign t[264] = t[318] ^ x[3];
  assign t[265] = t[319] ^ x[7];
  assign t[266] = t[320] ^ x[6];
  assign t[267] = t[321] ^ x[12];
  assign t[268] = t[322] ^ x[11];
  assign t[269] = t[323] ^ x[15];
  assign t[26] = t[47] ^ t[48];
  assign t[270] = t[324] ^ x[14];
  assign t[271] = t[325] ^ x[18];
  assign t[272] = t[326] ^ x[17];
  assign t[273] = t[327] ^ x[21];
  assign t[274] = t[328] ^ x[20];
  assign t[275] = t[329] ^ x[24];
  assign t[276] = t[330] ^ x[23];
  assign t[277] = t[331] ^ x[27];
  assign t[278] = t[332] ^ x[26];
  assign t[279] = t[333] ^ x[30];
  assign t[27] = t[49] & t[50];
  assign t[280] = t[334] ^ x[29];
  assign t[281] = t[335] ^ x[33];
  assign t[282] = t[336] ^ x[32];
  assign t[283] = t[337] ^ x[36];
  assign t[284] = t[338] ^ x[35];
  assign t[285] = t[339] ^ x[39];
  assign t[286] = t[340] ^ x[38];
  assign t[287] = t[341] ^ x[42];
  assign t[288] = t[342] ^ x[41];
  assign t[289] = t[343] ^ x[45];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[44];
  assign t[291] = t[345] ^ x[48];
  assign t[292] = t[346] ^ x[47];
  assign t[293] = t[347] ^ x[51];
  assign t[294] = t[348] ^ x[50];
  assign t[295] = t[349] ^ x[54];
  assign t[296] = t[350] ^ x[53];
  assign t[297] = t[351] ^ x[57];
  assign t[298] = t[352] ^ x[56];
  assign t[299] = t[353] ^ x[60];
  assign t[29] = ~(t[184] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[59];
  assign t[301] = t[355] ^ x[63];
  assign t[302] = t[356] ^ x[62];
  assign t[303] = t[357] ^ x[66];
  assign t[304] = t[358] ^ x[65];
  assign t[305] = t[359] ^ x[69];
  assign t[306] = t[360] ^ x[68];
  assign t[307] = t[361] ^ x[74];
  assign t[308] = t[362] ^ x[73];
  assign t[309] = t[363] ^ x[93];
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = t[364] ^ x[92];
  assign t[311] = t[365] ^ x[96];
  assign t[312] = t[366] ^ x[95];
  assign t[313] = t[367] ^ x[109];
  assign t[314] = t[368] ^ x[108];
  assign t[315] = t[369] ^ x[112];
  assign t[316] = t[370] ^ x[111];
  assign t[317] = (x[2]);
  assign t[318] = (x[2]);
  assign t[319] = (x[5]);
  assign t[31] = ~(t[55]);
  assign t[320] = (x[5]);
  assign t[321] = (x[10]);
  assign t[322] = (x[10]);
  assign t[323] = (x[13]);
  assign t[324] = (x[13]);
  assign t[325] = (x[16]);
  assign t[326] = (x[16]);
  assign t[327] = (x[19]);
  assign t[328] = (x[19]);
  assign t[329] = (x[22]);
  assign t[32] = ~(t[185]);
  assign t[330] = (x[22]);
  assign t[331] = (x[25]);
  assign t[332] = (x[25]);
  assign t[333] = (x[28]);
  assign t[334] = (x[28]);
  assign t[335] = (x[31]);
  assign t[336] = (x[31]);
  assign t[337] = (x[34]);
  assign t[338] = (x[34]);
  assign t[339] = (x[37]);
  assign t[33] = ~(t[186]);
  assign t[340] = (x[37]);
  assign t[341] = (x[40]);
  assign t[342] = (x[40]);
  assign t[343] = (x[43]);
  assign t[344] = (x[43]);
  assign t[345] = (x[46]);
  assign t[346] = (x[46]);
  assign t[347] = (x[49]);
  assign t[348] = (x[49]);
  assign t[349] = (x[52]);
  assign t[34] = ~(t[187]);
  assign t[350] = (x[52]);
  assign t[351] = (x[55]);
  assign t[352] = (x[55]);
  assign t[353] = (x[58]);
  assign t[354] = (x[58]);
  assign t[355] = (x[61]);
  assign t[356] = (x[61]);
  assign t[357] = (x[64]);
  assign t[358] = (x[64]);
  assign t[359] = (x[67]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = (x[67]);
  assign t[361] = (x[72]);
  assign t[362] = (x[72]);
  assign t[363] = (x[91]);
  assign t[364] = (x[91]);
  assign t[365] = (x[94]);
  assign t[366] = (x[94]);
  assign t[367] = (x[107]);
  assign t[368] = (x[107]);
  assign t[369] = (x[110]);
  assign t[36] = t[58] ^ t[59];
  assign t[370] = (x[110]);
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[38] = t[62] ^ t[63];
  assign t[39] = t[64] ^ t[65];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[66] : t[188];
  assign t[41] = t[189] ^ t[67];
  assign t[42] = ~(t[68]);
  assign t[43] = t[190] ^ t[69];
  assign t[44] = t[70] ^ t[64];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = t[73] ^ t[74];
  assign t[47] = t[75] ? t[76] : t[191];
  assign t[48] = t[75] ? t[77] : t[192];
  assign t[49] = ~(t[26] ^ t[78]);
  assign t[4] = t[8] ? t[9] : t[182];
  assign t[50] = t[79] ^ t[80];
  assign t[51] = ~(t[81] & t[82]);
  assign t[52] = t[83] ^ t[193];
  assign t[53] = ~(t[184]);
  assign t[54] = t[84] & t[83];
  assign t[55] = ~(t[85]);
  assign t[56] = ~(t[189]);
  assign t[57] = ~(t[86] & t[194]);
  assign t[58] = t[87] ^ t[88];
  assign t[59] = t[89] ^ t[90];
  assign t[5] = ~(t[10]);
  assign t[60] = ~(t[91] ^ t[92]);
  assign t[61] = t[93] ^ t[94];
  assign t[62] = t[95] ^ t[64];
  assign t[63] = t[96] & t[97];
  assign t[64] = t[75] ? t[98] : t[195];
  assign t[65] = t[71] ^ t[99];
  assign t[66] = t[188] ^ t[100];
  assign t[67] = t[101] ? t[102] : t[196];
  assign t[68] = t[187] ^ t[103];
  assign t[69] = t[8] ? t[104] : t[197];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[75] ? t[105] : t[198];
  assign t[71] = t[106] ^ t[63];
  assign t[72] = t[107] & t[108];
  assign t[73] = t[109] ^ t[23];
  assign t[74] = t[110] & t[111];
  assign t[75] = ~(t[112]);
  assign t[76] = t[191] ^ t[113];
  assign t[77] = t[192] ^ t[114];
  assign t[78] = t[115] ^ t[90];
  assign t[79] = t[48] ^ t[87];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[75] ? t[116] : t[199];
  assign t[81] = ~(t[84] | t[83]);
  assign t[82] = ~(t[117] | t[53]);
  assign t[83] = ~(t[200]);
  assign t[84] = ~(t[193]);
  assign t[85] = ~(t[16]);
  assign t[86] = ~(t[190]);
  assign t[87] = t[75] ? t[118] : t[201];
  assign t[88] = t[78] ^ t[27];
  assign t[89] = t[47] ^ t[87];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[119] & t[80];
  assign t[91] = t[120] ^ t[74];
  assign t[92] = t[121] ^ t[122];
  assign t[93] = t[123] ^ t[121];
  assign t[94] = t[124] ^ t[125];
  assign t[95] = t[75] ? t[126] : t[202];
  assign t[96] = ~(t[70]);
  assign t[97] = t[75] ? t[127] : t[203];
  assign t[98] = t[195] ^ t[128];
  assign t[99] = t[129] & t[130];
  assign t[9] = t[182] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind62(x, y);
 input [116:0] x;
 output y;

 wire [361:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[186] ^ t[133];
  assign t[101] = t[134] & t[135];
  assign t[102] = t[136] & t[70];
  assign t[103] = t[184] ^ t[137];
  assign t[104] = t[8] ? t[138] : t[191];
  assign t[105] = t[132] ? x[66] : x[65];
  assign t[106] = t[132] ? x[68] : x[67];
  assign t[107] = ~(t[113]);
  assign t[108] = ~(t[91]);
  assign t[109] = ~(t[44]);
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[48] ? t[139] : t[192];
  assign t[111] = t[24] ^ t[91];
  assign t[112] = t[91] ^ t[45];
  assign t[113] = t[110] ^ t[44];
  assign t[114] = ~(t[140]);
  assign t[115] = ~(t[141]);
  assign t[116] = ~(t[126]);
  assign t[117] = ~(t[127]);
  assign t[118] = t[48] ? t[142] : t[193];
  assign t[119] = t[127] ^ t[26];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = ~(t[174]);
  assign t[121] = t[8] ? t[143] : t[194];
  assign t[122] = t[144];
  assign t[123] = t[8] ? t[145] : t[195];
  assign t[124] = t[189] ^ t[146];
  assign t[125] = t[147] & t[148];
  assign t[126] = t[48] ? t[149] : t[196];
  assign t[127] = t[48] ? t[150] : t[197];
  assign t[128] = t[190] ^ t[151];
  assign t[129] = t[152] & t[153];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = ~(t[154] ^ t[97]);
  assign t[131] = t[155] ^ t[90];
  assign t[132] = ~(t[140]);
  assign t[133] = t[132] ? x[88] : x[87];
  assign t[134] = ~(t[156]);
  assign t[135] = ~(t[40]);
  assign t[136] = ~(t[41]);
  assign t[137] = t[157] ? t[158] : t[198];
  assign t[138] = t[191] ^ t[159];
  assign t[139] = t[192] ^ t[160];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[31]);
  assign t[141] = t[118] ^ t[127];
  assign t[142] = t[193] ^ t[161];
  assign t[143] = t[194] ^ t[162];
  assign t[144] = t[8] ? t[163] : t[199];
  assign t[145] = t[195] ^ t[164];
  assign t[146] = t[132] ? x[96] : x[95];
  assign t[147] = ~(t[101] ^ t[165]);
  assign t[148] = t[166] ^ t[156];
  assign t[149] = t[196] ^ t[167];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[197] ^ t[168];
  assign t[151] = t[31] ? x[98] : x[97];
  assign t[152] = ~(t[169]);
  assign t[153] = ~(t[88]);
  assign t[154] = t[88] ^ t[122];
  assign t[155] = t[122] ^ t[64];
  assign t[156] = t[70] ^ t[41];
  assign t[157] = ~(t[77]);
  assign t[158] = t[198] ^ t[170];
  assign t[159] = t[31] ? x[100] : x[99];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[132] ? x[102] : x[101];
  assign t[161] = t[114] ? x[104] : x[103];
  assign t[162] = t[31] ? x[106] : x[105];
  assign t[163] = t[199] ^ t[171];
  assign t[164] = t[172] ? x[108] : x[107];
  assign t[165] = t[69] ^ t[40];
  assign t[166] = t[40] ^ t[103];
  assign t[167] = t[114] ? x[110] : x[109];
  assign t[168] = t[114] ? x[112] : x[111];
  assign t[169] = t[90] ^ t[122];
  assign t[16] = t[174] | t[30];
  assign t[170] = t[172] ? x[114] : x[113];
  assign t[171] = t[172] ? x[116] : x[115];
  assign t[172] = ~(t[140]);
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[4];
  assign t[201] = t[228] ^ x[7];
  assign t[202] = t[229] ^ x[12];
  assign t[203] = t[230] ^ x[15];
  assign t[204] = t[231] ^ x[18];
  assign t[205] = t[232] ^ x[21];
  assign t[206] = t[233] ^ x[24];
  assign t[207] = t[234] ^ x[27];
  assign t[208] = t[235] ^ x[30];
  assign t[209] = t[236] ^ x[33];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[36];
  assign t[211] = t[238] ^ x[39];
  assign t[212] = t[239] ^ x[42];
  assign t[213] = t[240] ^ x[45];
  assign t[214] = t[241] ^ x[48];
  assign t[215] = t[242] ^ x[53];
  assign t[216] = t[243] ^ x[56];
  assign t[217] = t[244] ^ x[59];
  assign t[218] = t[245] ^ x[64];
  assign t[219] = t[246] ^ x[71];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[74];
  assign t[221] = t[248] ^ x[77];
  assign t[222] = t[249] ^ x[80];
  assign t[223] = t[250] ^ x[83];
  assign t[224] = t[251] ^ x[86];
  assign t[225] = t[252] ^ x[91];
  assign t[226] = t[253] ^ x[94];
  assign t[227] = (t[254] & ~t[255]);
  assign t[228] = (t[256] & ~t[257]);
  assign t[229] = (t[258] & ~t[259]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[260] & ~t[261]);
  assign t[231] = (t[262] & ~t[263]);
  assign t[232] = (t[264] & ~t[265]);
  assign t[233] = (t[266] & ~t[267]);
  assign t[234] = (t[268] & ~t[269]);
  assign t[235] = (t[270] & ~t[271]);
  assign t[236] = (t[272] & ~t[273]);
  assign t[237] = (t[274] & ~t[275]);
  assign t[238] = (t[276] & ~t[277]);
  assign t[239] = (t[278] & ~t[279]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[280] & ~t[281]);
  assign t[241] = (t[282] & ~t[283]);
  assign t[242] = (t[284] & ~t[285]);
  assign t[243] = (t[286] & ~t[287]);
  assign t[244] = (t[288] & ~t[289]);
  assign t[245] = (t[290] & ~t[291]);
  assign t[246] = (t[292] & ~t[293]);
  assign t[247] = (t[294] & ~t[295]);
  assign t[248] = (t[296] & ~t[297]);
  assign t[249] = (t[298] & ~t[299]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[300] & ~t[301]);
  assign t[251] = (t[302] & ~t[303]);
  assign t[252] = (t[304] & ~t[305]);
  assign t[253] = (t[306] & ~t[307]);
  assign t[254] = t[308] ^ x[4];
  assign t[255] = t[309] ^ x[3];
  assign t[256] = t[310] ^ x[7];
  assign t[257] = t[311] ^ x[6];
  assign t[258] = t[312] ^ x[12];
  assign t[259] = t[313] ^ x[11];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[314] ^ x[15];
  assign t[261] = t[315] ^ x[14];
  assign t[262] = t[316] ^ x[18];
  assign t[263] = t[317] ^ x[17];
  assign t[264] = t[318] ^ x[21];
  assign t[265] = t[319] ^ x[20];
  assign t[266] = t[320] ^ x[24];
  assign t[267] = t[321] ^ x[23];
  assign t[268] = t[322] ^ x[27];
  assign t[269] = t[323] ^ x[26];
  assign t[26] = t[48] ? t[49] : t[175];
  assign t[270] = t[324] ^ x[30];
  assign t[271] = t[325] ^ x[29];
  assign t[272] = t[326] ^ x[33];
  assign t[273] = t[327] ^ x[32];
  assign t[274] = t[328] ^ x[36];
  assign t[275] = t[329] ^ x[35];
  assign t[276] = t[330] ^ x[39];
  assign t[277] = t[331] ^ x[38];
  assign t[278] = t[332] ^ x[42];
  assign t[279] = t[333] ^ x[41];
  assign t[27] = t[50] ^ t[51];
  assign t[280] = t[334] ^ x[45];
  assign t[281] = t[335] ^ x[44];
  assign t[282] = t[336] ^ x[48];
  assign t[283] = t[337] ^ x[47];
  assign t[284] = t[338] ^ x[53];
  assign t[285] = t[339] ^ x[52];
  assign t[286] = t[340] ^ x[56];
  assign t[287] = t[341] ^ x[55];
  assign t[288] = t[342] ^ x[59];
  assign t[289] = t[343] ^ x[58];
  assign t[28] = ~(t[30] & t[52]);
  assign t[290] = t[344] ^ x[64];
  assign t[291] = t[345] ^ x[63];
  assign t[292] = t[346] ^ x[71];
  assign t[293] = t[347] ^ x[70];
  assign t[294] = t[348] ^ x[74];
  assign t[295] = t[349] ^ x[73];
  assign t[296] = t[350] ^ x[77];
  assign t[297] = t[351] ^ x[76];
  assign t[298] = t[352] ^ x[80];
  assign t[299] = t[353] ^ x[79];
  assign t[29] = ~(t[176] ^ t[53]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[83];
  assign t[301] = t[355] ^ x[82];
  assign t[302] = t[356] ^ x[86];
  assign t[303] = t[357] ^ x[85];
  assign t[304] = t[358] ^ x[91];
  assign t[305] = t[359] ^ x[90];
  assign t[306] = t[360] ^ x[94];
  assign t[307] = t[361] ^ x[93];
  assign t[308] = (x[2]);
  assign t[309] = (x[2]);
  assign t[30] = ~(t[54] & t[55]);
  assign t[310] = (x[5]);
  assign t[311] = (x[5]);
  assign t[312] = (x[10]);
  assign t[313] = (x[10]);
  assign t[314] = (x[13]);
  assign t[315] = (x[13]);
  assign t[316] = (x[16]);
  assign t[317] = (x[16]);
  assign t[318] = (x[19]);
  assign t[319] = (x[19]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[22]);
  assign t[321] = (x[22]);
  assign t[322] = (x[25]);
  assign t[323] = (x[25]);
  assign t[324] = (x[28]);
  assign t[325] = (x[28]);
  assign t[326] = (x[31]);
  assign t[327] = (x[31]);
  assign t[328] = (x[34]);
  assign t[329] = (x[34]);
  assign t[32] = ~(t[177]);
  assign t[330] = (x[37]);
  assign t[331] = (x[37]);
  assign t[332] = (x[40]);
  assign t[333] = (x[40]);
  assign t[334] = (x[43]);
  assign t[335] = (x[43]);
  assign t[336] = (x[46]);
  assign t[337] = (x[46]);
  assign t[338] = (x[51]);
  assign t[339] = (x[51]);
  assign t[33] = ~(t[178]);
  assign t[340] = (x[54]);
  assign t[341] = (x[54]);
  assign t[342] = (x[57]);
  assign t[343] = (x[57]);
  assign t[344] = (x[62]);
  assign t[345] = (x[62]);
  assign t[346] = (x[69]);
  assign t[347] = (x[69]);
  assign t[348] = (x[72]);
  assign t[349] = (x[72]);
  assign t[34] = ~(t[179]);
  assign t[350] = (x[75]);
  assign t[351] = (x[75]);
  assign t[352] = (x[78]);
  assign t[353] = (x[78]);
  assign t[354] = (x[81]);
  assign t[355] = (x[81]);
  assign t[356] = (x[84]);
  assign t[357] = (x[84]);
  assign t[358] = (x[89]);
  assign t[359] = (x[89]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = (x[92]);
  assign t[361] = (x[92]);
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[62] ^ t[63];
  assign t[39] = t[64] ^ t[65];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[66] : t[180];
  assign t[41] = t[179] ^ t[67];
  assign t[42] = ~(t[22] ^ t[68]);
  assign t[43] = t[69] ^ t[70];
  assign t[44] = t[48] ? t[71] : t[181];
  assign t[45] = t[48] ? t[72] : t[182];
  assign t[46] = t[73] ^ t[74];
  assign t[47] = t[75] & t[76];
  assign t[48] = ~(t[77]);
  assign t[49] = t[175] ^ t[78];
  assign t[4] = t[8] ? t[9] : t[173];
  assign t[50] = t[79] ^ t[80];
  assign t[51] = t[81] & t[82];
  assign t[52] = ~(t[83] & t[84]);
  assign t[53] = t[85] ^ t[183];
  assign t[54] = ~(t[176]);
  assign t[55] = t[86] & t[85];
  assign t[56] = ~(t[184]);
  assign t[57] = ~(t[87] & t[185]);
  assign t[58] = t[88] ^ t[64];
  assign t[59] = t[89] & t[90];
  assign t[5] = ~(t[10]);
  assign t[60] = t[91] ^ t[44];
  assign t[61] = t[92] & t[93];
  assign t[62] = t[69] ^ t[94];
  assign t[63] = t[95] ^ t[51];
  assign t[64] = t[96];
  assign t[65] = t[97] ^ t[98];
  assign t[66] = t[180] ^ t[99];
  assign t[67] = t[8] ? t[100] : t[186];
  assign t[68] = t[101] ^ t[102];
  assign t[69] = t[41] ^ t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[187] ^ t[104];
  assign t[71] = t[181] ^ t[105];
  assign t[72] = t[182] ^ t[106];
  assign t[73] = t[107] & t[108];
  assign t[74] = t[109] & t[110];
  assign t[75] = ~(t[73] ^ t[111]);
  assign t[76] = t[112] ^ t[113];
  assign t[77] = ~(t[8]);
  assign t[78] = t[114] ? x[50] : x[49];
  assign t[79] = t[115] & t[116];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] & t[118];
  assign t[81] = ~(t[95] ^ t[50]);
  assign t[82] = t[119] ^ t[118];
  assign t[83] = ~(t[86] | t[85]);
  assign t[84] = ~(t[120] | t[54]);
  assign t[85] = ~(t[188]);
  assign t[86] = ~(t[183]);
  assign t[87] = ~(t[187]);
  assign t[88] = ~t[121];
  assign t[89] = ~(t[122]);
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[123];
  assign t[91] = t[48] ? t[124] : t[189];
  assign t[92] = ~(t[60] ^ t[46]);
  assign t[93] = t[24] ^ t[110];
  assign t[94] = t[68] ^ t[125];
  assign t[95] = t[126] ^ t[127];
  assign t[96] = t[8] ? t[128] : t[190];
  assign t[97] = t[129] ^ t[59];
  assign t[98] = t[130] & t[131];
  assign t[99] = t[132] ? x[61] : x[60];
  assign t[9] = t[173] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind63(x, y);
 input [116:0] x;
 output y;

 wire [361:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[186] ^ t[133];
  assign t[101] = t[134] & t[135];
  assign t[102] = t[136] & t[70];
  assign t[103] = t[184] ^ t[137];
  assign t[104] = t[8] ? t[138] : t[191];
  assign t[105] = t[132] ? x[66] : x[65];
  assign t[106] = t[132] ? x[68] : x[67];
  assign t[107] = ~(t[113]);
  assign t[108] = ~(t[91]);
  assign t[109] = ~(t[44]);
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[48] ? t[139] : t[192];
  assign t[111] = t[24] ^ t[91];
  assign t[112] = t[91] ^ t[45];
  assign t[113] = t[110] ^ t[44];
  assign t[114] = ~(t[140]);
  assign t[115] = ~(t[141]);
  assign t[116] = ~(t[126]);
  assign t[117] = ~(t[127]);
  assign t[118] = t[48] ? t[142] : t[193];
  assign t[119] = t[127] ^ t[26];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = ~(t[174]);
  assign t[121] = t[8] ? t[143] : t[194];
  assign t[122] = t[144];
  assign t[123] = t[8] ? t[145] : t[195];
  assign t[124] = t[189] ^ t[146];
  assign t[125] = t[147] & t[148];
  assign t[126] = t[48] ? t[149] : t[196];
  assign t[127] = t[48] ? t[150] : t[197];
  assign t[128] = t[190] ^ t[151];
  assign t[129] = t[152] & t[153];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = ~(t[154] ^ t[97]);
  assign t[131] = t[155] ^ t[90];
  assign t[132] = ~(t[140]);
  assign t[133] = t[132] ? x[88] : x[87];
  assign t[134] = ~(t[156]);
  assign t[135] = ~(t[40]);
  assign t[136] = ~(t[41]);
  assign t[137] = t[157] ? t[158] : t[198];
  assign t[138] = t[191] ^ t[159];
  assign t[139] = t[192] ^ t[160];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[31]);
  assign t[141] = t[118] ^ t[127];
  assign t[142] = t[193] ^ t[161];
  assign t[143] = t[194] ^ t[162];
  assign t[144] = t[8] ? t[163] : t[199];
  assign t[145] = t[195] ^ t[164];
  assign t[146] = t[132] ? x[96] : x[95];
  assign t[147] = ~(t[101] ^ t[165]);
  assign t[148] = t[166] ^ t[156];
  assign t[149] = t[196] ^ t[167];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[197] ^ t[168];
  assign t[151] = t[31] ? x[98] : x[97];
  assign t[152] = ~(t[169]);
  assign t[153] = ~(t[88]);
  assign t[154] = t[88] ^ t[122];
  assign t[155] = t[122] ^ t[64];
  assign t[156] = t[70] ^ t[41];
  assign t[157] = ~(t[77]);
  assign t[158] = t[198] ^ t[170];
  assign t[159] = t[31] ? x[100] : x[99];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[132] ? x[102] : x[101];
  assign t[161] = t[114] ? x[104] : x[103];
  assign t[162] = t[31] ? x[106] : x[105];
  assign t[163] = t[199] ^ t[171];
  assign t[164] = t[172] ? x[108] : x[107];
  assign t[165] = t[69] ^ t[40];
  assign t[166] = t[40] ^ t[103];
  assign t[167] = t[114] ? x[110] : x[109];
  assign t[168] = t[114] ? x[112] : x[111];
  assign t[169] = t[90] ^ t[122];
  assign t[16] = t[174] | t[30];
  assign t[170] = t[172] ? x[114] : x[113];
  assign t[171] = t[172] ? x[116] : x[115];
  assign t[172] = ~(t[140]);
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[4];
  assign t[201] = t[228] ^ x[7];
  assign t[202] = t[229] ^ x[12];
  assign t[203] = t[230] ^ x[15];
  assign t[204] = t[231] ^ x[18];
  assign t[205] = t[232] ^ x[21];
  assign t[206] = t[233] ^ x[24];
  assign t[207] = t[234] ^ x[27];
  assign t[208] = t[235] ^ x[30];
  assign t[209] = t[236] ^ x[33];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[36];
  assign t[211] = t[238] ^ x[39];
  assign t[212] = t[239] ^ x[42];
  assign t[213] = t[240] ^ x[45];
  assign t[214] = t[241] ^ x[48];
  assign t[215] = t[242] ^ x[53];
  assign t[216] = t[243] ^ x[56];
  assign t[217] = t[244] ^ x[59];
  assign t[218] = t[245] ^ x[64];
  assign t[219] = t[246] ^ x[71];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[74];
  assign t[221] = t[248] ^ x[77];
  assign t[222] = t[249] ^ x[80];
  assign t[223] = t[250] ^ x[83];
  assign t[224] = t[251] ^ x[86];
  assign t[225] = t[252] ^ x[91];
  assign t[226] = t[253] ^ x[94];
  assign t[227] = (t[254] & ~t[255]);
  assign t[228] = (t[256] & ~t[257]);
  assign t[229] = (t[258] & ~t[259]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[260] & ~t[261]);
  assign t[231] = (t[262] & ~t[263]);
  assign t[232] = (t[264] & ~t[265]);
  assign t[233] = (t[266] & ~t[267]);
  assign t[234] = (t[268] & ~t[269]);
  assign t[235] = (t[270] & ~t[271]);
  assign t[236] = (t[272] & ~t[273]);
  assign t[237] = (t[274] & ~t[275]);
  assign t[238] = (t[276] & ~t[277]);
  assign t[239] = (t[278] & ~t[279]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[280] & ~t[281]);
  assign t[241] = (t[282] & ~t[283]);
  assign t[242] = (t[284] & ~t[285]);
  assign t[243] = (t[286] & ~t[287]);
  assign t[244] = (t[288] & ~t[289]);
  assign t[245] = (t[290] & ~t[291]);
  assign t[246] = (t[292] & ~t[293]);
  assign t[247] = (t[294] & ~t[295]);
  assign t[248] = (t[296] & ~t[297]);
  assign t[249] = (t[298] & ~t[299]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[300] & ~t[301]);
  assign t[251] = (t[302] & ~t[303]);
  assign t[252] = (t[304] & ~t[305]);
  assign t[253] = (t[306] & ~t[307]);
  assign t[254] = t[308] ^ x[4];
  assign t[255] = t[309] ^ x[3];
  assign t[256] = t[310] ^ x[7];
  assign t[257] = t[311] ^ x[6];
  assign t[258] = t[312] ^ x[12];
  assign t[259] = t[313] ^ x[11];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[314] ^ x[15];
  assign t[261] = t[315] ^ x[14];
  assign t[262] = t[316] ^ x[18];
  assign t[263] = t[317] ^ x[17];
  assign t[264] = t[318] ^ x[21];
  assign t[265] = t[319] ^ x[20];
  assign t[266] = t[320] ^ x[24];
  assign t[267] = t[321] ^ x[23];
  assign t[268] = t[322] ^ x[27];
  assign t[269] = t[323] ^ x[26];
  assign t[26] = t[48] ? t[49] : t[175];
  assign t[270] = t[324] ^ x[30];
  assign t[271] = t[325] ^ x[29];
  assign t[272] = t[326] ^ x[33];
  assign t[273] = t[327] ^ x[32];
  assign t[274] = t[328] ^ x[36];
  assign t[275] = t[329] ^ x[35];
  assign t[276] = t[330] ^ x[39];
  assign t[277] = t[331] ^ x[38];
  assign t[278] = t[332] ^ x[42];
  assign t[279] = t[333] ^ x[41];
  assign t[27] = t[50] ^ t[51];
  assign t[280] = t[334] ^ x[45];
  assign t[281] = t[335] ^ x[44];
  assign t[282] = t[336] ^ x[48];
  assign t[283] = t[337] ^ x[47];
  assign t[284] = t[338] ^ x[53];
  assign t[285] = t[339] ^ x[52];
  assign t[286] = t[340] ^ x[56];
  assign t[287] = t[341] ^ x[55];
  assign t[288] = t[342] ^ x[59];
  assign t[289] = t[343] ^ x[58];
  assign t[28] = ~(t[30] & t[52]);
  assign t[290] = t[344] ^ x[64];
  assign t[291] = t[345] ^ x[63];
  assign t[292] = t[346] ^ x[71];
  assign t[293] = t[347] ^ x[70];
  assign t[294] = t[348] ^ x[74];
  assign t[295] = t[349] ^ x[73];
  assign t[296] = t[350] ^ x[77];
  assign t[297] = t[351] ^ x[76];
  assign t[298] = t[352] ^ x[80];
  assign t[299] = t[353] ^ x[79];
  assign t[29] = ~(t[176] ^ t[53]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[83];
  assign t[301] = t[355] ^ x[82];
  assign t[302] = t[356] ^ x[86];
  assign t[303] = t[357] ^ x[85];
  assign t[304] = t[358] ^ x[91];
  assign t[305] = t[359] ^ x[90];
  assign t[306] = t[360] ^ x[94];
  assign t[307] = t[361] ^ x[93];
  assign t[308] = (x[2]);
  assign t[309] = (x[2]);
  assign t[30] = ~(t[54] & t[55]);
  assign t[310] = (x[5]);
  assign t[311] = (x[5]);
  assign t[312] = (x[10]);
  assign t[313] = (x[10]);
  assign t[314] = (x[13]);
  assign t[315] = (x[13]);
  assign t[316] = (x[16]);
  assign t[317] = (x[16]);
  assign t[318] = (x[19]);
  assign t[319] = (x[19]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[22]);
  assign t[321] = (x[22]);
  assign t[322] = (x[25]);
  assign t[323] = (x[25]);
  assign t[324] = (x[28]);
  assign t[325] = (x[28]);
  assign t[326] = (x[31]);
  assign t[327] = (x[31]);
  assign t[328] = (x[34]);
  assign t[329] = (x[34]);
  assign t[32] = ~(t[177]);
  assign t[330] = (x[37]);
  assign t[331] = (x[37]);
  assign t[332] = (x[40]);
  assign t[333] = (x[40]);
  assign t[334] = (x[43]);
  assign t[335] = (x[43]);
  assign t[336] = (x[46]);
  assign t[337] = (x[46]);
  assign t[338] = (x[51]);
  assign t[339] = (x[51]);
  assign t[33] = ~(t[178]);
  assign t[340] = (x[54]);
  assign t[341] = (x[54]);
  assign t[342] = (x[57]);
  assign t[343] = (x[57]);
  assign t[344] = (x[62]);
  assign t[345] = (x[62]);
  assign t[346] = (x[69]);
  assign t[347] = (x[69]);
  assign t[348] = (x[72]);
  assign t[349] = (x[72]);
  assign t[34] = ~(t[179]);
  assign t[350] = (x[75]);
  assign t[351] = (x[75]);
  assign t[352] = (x[78]);
  assign t[353] = (x[78]);
  assign t[354] = (x[81]);
  assign t[355] = (x[81]);
  assign t[356] = (x[84]);
  assign t[357] = (x[84]);
  assign t[358] = (x[89]);
  assign t[359] = (x[89]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = (x[92]);
  assign t[361] = (x[92]);
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[62] ^ t[63];
  assign t[39] = t[64] ^ t[65];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[66] : t[180];
  assign t[41] = t[179] ^ t[67];
  assign t[42] = ~(t[22] ^ t[68]);
  assign t[43] = t[69] ^ t[70];
  assign t[44] = t[48] ? t[71] : t[181];
  assign t[45] = t[48] ? t[72] : t[182];
  assign t[46] = t[73] ^ t[74];
  assign t[47] = t[75] & t[76];
  assign t[48] = ~(t[77]);
  assign t[49] = t[175] ^ t[78];
  assign t[4] = t[8] ? t[9] : t[173];
  assign t[50] = t[79] ^ t[80];
  assign t[51] = t[81] & t[82];
  assign t[52] = ~(t[83] & t[84]);
  assign t[53] = t[85] ^ t[183];
  assign t[54] = ~(t[176]);
  assign t[55] = t[86] & t[85];
  assign t[56] = ~(t[184]);
  assign t[57] = ~(t[87] & t[185]);
  assign t[58] = t[88] ^ t[64];
  assign t[59] = t[89] & t[90];
  assign t[5] = ~(t[10]);
  assign t[60] = t[91] ^ t[44];
  assign t[61] = t[92] & t[93];
  assign t[62] = t[69] ^ t[94];
  assign t[63] = t[95] ^ t[51];
  assign t[64] = t[96];
  assign t[65] = t[97] ^ t[98];
  assign t[66] = t[180] ^ t[99];
  assign t[67] = t[8] ? t[100] : t[186];
  assign t[68] = t[101] ^ t[102];
  assign t[69] = t[41] ^ t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[187] ^ t[104];
  assign t[71] = t[181] ^ t[105];
  assign t[72] = t[182] ^ t[106];
  assign t[73] = t[107] & t[108];
  assign t[74] = t[109] & t[110];
  assign t[75] = ~(t[73] ^ t[111]);
  assign t[76] = t[112] ^ t[113];
  assign t[77] = ~(t[8]);
  assign t[78] = t[114] ? x[50] : x[49];
  assign t[79] = t[115] & t[116];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] & t[118];
  assign t[81] = ~(t[95] ^ t[50]);
  assign t[82] = t[119] ^ t[118];
  assign t[83] = ~(t[86] | t[85]);
  assign t[84] = ~(t[120] | t[54]);
  assign t[85] = ~(t[188]);
  assign t[86] = ~(t[183]);
  assign t[87] = ~(t[187]);
  assign t[88] = ~t[121];
  assign t[89] = ~(t[122]);
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[123];
  assign t[91] = t[48] ? t[124] : t[189];
  assign t[92] = ~(t[60] ^ t[46]);
  assign t[93] = t[24] ^ t[110];
  assign t[94] = t[68] ^ t[125];
  assign t[95] = t[126] ^ t[127];
  assign t[96] = t[8] ? t[128] : t[190];
  assign t[97] = t[129] ^ t[59];
  assign t[98] = t[130] & t[131];
  assign t[99] = t[132] ? x[61] : x[60];
  assign t[9] = t[173] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind64(x, y);
 input [116:0] x;
 output y;

 wire [360:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[53] ? t[126] : t[190];
  assign t[101] = ~(t[71] ^ t[127]);
  assign t[102] = t[128] ^ t[129];
  assign t[103] = t[113] ? x[72] : x[71];
  assign t[104] = ~(t[129]);
  assign t[105] = ~(t[130]);
  assign t[106] = ~(t[68]);
  assign t[107] = t[131];
  assign t[108] = t[130] ^ t[68];
  assign t[109] = ~(t[132] & t[133]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[134] ^ t[191];
  assign t[111] = ~(t[186]);
  assign t[112] = t[135] & t[134];
  assign t[113] = ~(t[50]);
  assign t[114] = t[113] ? x[77] : x[76];
  assign t[115] = ~(t[50]);
  assign t[116] = t[27] ? t[136] : t[192];
  assign t[117] = t[188] ^ t[137];
  assign t[118] = t[138] ^ t[20];
  assign t[119] = t[139] & t[140];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[141] & t[142];
  assign t[121] = t[189] ^ t[143];
  assign t[122] = t[8] ? t[144] : t[193];
  assign t[123] = t[145] ^ t[146];
  assign t[124] = t[97] ^ t[147];
  assign t[125] = t[174] ^ t[148];
  assign t[126] = t[190] ^ t[149];
  assign t[127] = t[43] ^ t[130];
  assign t[128] = t[130] ^ t[25];
  assign t[129] = t[107] ^ t[68];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[150];
  assign t[131] = t[27] ? t[151] : t[194];
  assign t[132] = ~(t[135] | t[134]);
  assign t[133] = ~(t[152] | t[111]);
  assign t[134] = ~(t[195]);
  assign t[135] = ~(t[191]);
  assign t[136] = t[192] ^ t[153];
  assign t[137] = t[78] ? x[91] : x[90];
  assign t[138] = t[154] & t[155];
  assign t[139] = ~(t[138] ^ t[156]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[19] ^ t[157];
  assign t[141] = ~(t[158] ^ t[39]);
  assign t[142] = t[21] ^ t[89];
  assign t[143] = t[28] ? x[93] : x[92];
  assign t[144] = t[193] ^ t[159];
  assign t[145] = t[160] & t[161];
  assign t[146] = t[162] & t[125];
  assign t[147] = t[184] ^ t[163];
  assign t[148] = t[8] ? t[164] : t[196];
  assign t[149] = t[113] ? x[98] : x[97];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[53] ? t[165] : t[197];
  assign t[151] = t[194] ^ t[166];
  assign t[152] = ~(t[182]);
  assign t[153] = t[115] ? x[103] : x[102];
  assign t[154] = ~(t[157]);
  assign t[155] = ~(t[33]);
  assign t[156] = t[93] ^ t[33];
  assign t[157] = t[36] ^ t[56];
  assign t[158] = t[116] ^ t[37];
  assign t[159] = t[28] ? x[105] : x[104];
  assign t[15] = ~(t[27]);
  assign t[160] = ~(t[167]);
  assign t[161] = ~(t[96]);
  assign t[162] = ~(t[97]);
  assign t[163] = t[8] ? t[168] : t[198];
  assign t[164] = t[196] ^ t[169];
  assign t[165] = t[197] ^ t[170];
  assign t[166] = t[113] ? x[110] : x[109];
  assign t[167] = t[125] ^ t[97];
  assign t[168] = t[198] ^ t[171];
  assign t[169] = t[28] ? x[112] : x[111];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[113] ? x[114] : x[113];
  assign t[171] = t[28] ? x[116] : x[115];
  assign t[172] = (t[199]);
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = t[226] ^ x[4];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[9];
  assign t[201] = t[228] ^ x[12];
  assign t[202] = t[229] ^ x[15];
  assign t[203] = t[230] ^ x[18];
  assign t[204] = t[231] ^ x[21];
  assign t[205] = t[232] ^ x[24];
  assign t[206] = t[233] ^ x[27];
  assign t[207] = t[234] ^ x[30];
  assign t[208] = t[235] ^ x[33];
  assign t[209] = t[236] ^ x[36];
  assign t[20] = t[35] & t[36];
  assign t[210] = t[237] ^ x[39];
  assign t[211] = t[238] ^ x[42];
  assign t[212] = t[239] ^ x[45];
  assign t[213] = t[240] ^ x[48];
  assign t[214] = t[241] ^ x[51];
  assign t[215] = t[242] ^ x[64];
  assign t[216] = t[243] ^ x[67];
  assign t[217] = t[244] ^ x[70];
  assign t[218] = t[245] ^ x[75];
  assign t[219] = t[246] ^ x[80];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[83];
  assign t[221] = t[248] ^ x[86];
  assign t[222] = t[249] ^ x[89];
  assign t[223] = t[250] ^ x[96];
  assign t[224] = t[251] ^ x[101];
  assign t[225] = t[252] ^ x[108];
  assign t[226] = (t[253] & ~t[254]);
  assign t[227] = (t[255] & ~t[256]);
  assign t[228] = (t[257] & ~t[258]);
  assign t[229] = (t[259] & ~t[260]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[261] & ~t[262]);
  assign t[231] = (t[263] & ~t[264]);
  assign t[232] = (t[265] & ~t[266]);
  assign t[233] = (t[267] & ~t[268]);
  assign t[234] = (t[269] & ~t[270]);
  assign t[235] = (t[271] & ~t[272]);
  assign t[236] = (t[273] & ~t[274]);
  assign t[237] = (t[275] & ~t[276]);
  assign t[238] = (t[277] & ~t[278]);
  assign t[239] = (t[279] & ~t[280]);
  assign t[23] = ~(t[41] ^ t[42]);
  assign t[240] = (t[281] & ~t[282]);
  assign t[241] = (t[283] & ~t[284]);
  assign t[242] = (t[285] & ~t[286]);
  assign t[243] = (t[287] & ~t[288]);
  assign t[244] = (t[289] & ~t[290]);
  assign t[245] = (t[291] & ~t[292]);
  assign t[246] = (t[293] & ~t[294]);
  assign t[247] = (t[295] & ~t[296]);
  assign t[248] = (t[297] & ~t[298]);
  assign t[249] = (t[299] & ~t[300]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (t[301] & ~t[302]);
  assign t[251] = (t[303] & ~t[304]);
  assign t[252] = (t[305] & ~t[306]);
  assign t[253] = t[307] ^ x[4];
  assign t[254] = t[308] ^ x[3];
  assign t[255] = t[309] ^ x[9];
  assign t[256] = t[310] ^ x[8];
  assign t[257] = t[311] ^ x[12];
  assign t[258] = t[312] ^ x[11];
  assign t[259] = t[313] ^ x[15];
  assign t[25] = ~t[45];
  assign t[260] = t[314] ^ x[14];
  assign t[261] = t[315] ^ x[18];
  assign t[262] = t[316] ^ x[17];
  assign t[263] = t[317] ^ x[21];
  assign t[264] = t[318] ^ x[20];
  assign t[265] = t[319] ^ x[24];
  assign t[266] = t[320] ^ x[23];
  assign t[267] = t[321] ^ x[27];
  assign t[268] = t[322] ^ x[26];
  assign t[269] = t[323] ^ x[30];
  assign t[26] = t[46] ^ t[47];
  assign t[270] = t[324] ^ x[29];
  assign t[271] = t[325] ^ x[33];
  assign t[272] = t[326] ^ x[32];
  assign t[273] = t[327] ^ x[36];
  assign t[274] = t[328] ^ x[35];
  assign t[275] = t[329] ^ x[39];
  assign t[276] = t[330] ^ x[38];
  assign t[277] = t[331] ^ x[42];
  assign t[278] = t[332] ^ x[41];
  assign t[279] = t[333] ^ x[45];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[44];
  assign t[281] = t[335] ^ x[48];
  assign t[282] = t[336] ^ x[47];
  assign t[283] = t[337] ^ x[51];
  assign t[284] = t[338] ^ x[50];
  assign t[285] = t[339] ^ x[64];
  assign t[286] = t[340] ^ x[63];
  assign t[287] = t[341] ^ x[67];
  assign t[288] = t[342] ^ x[66];
  assign t[289] = t[343] ^ x[70];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[69];
  assign t[291] = t[345] ^ x[75];
  assign t[292] = t[346] ^ x[74];
  assign t[293] = t[347] ^ x[80];
  assign t[294] = t[348] ^ x[79];
  assign t[295] = t[349] ^ x[83];
  assign t[296] = t[350] ^ x[82];
  assign t[297] = t[351] ^ x[86];
  assign t[298] = t[352] ^ x[85];
  assign t[299] = t[353] ^ x[89];
  assign t[29] = ~(t[173]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[88];
  assign t[301] = t[355] ^ x[96];
  assign t[302] = t[356] ^ x[95];
  assign t[303] = t[357] ^ x[101];
  assign t[304] = t[358] ^ x[100];
  assign t[305] = t[359] ^ x[108];
  assign t[306] = t[360] ^ x[107];
  assign t[307] = (x[2]);
  assign t[308] = (x[2]);
  assign t[309] = (x[7]);
  assign t[30] = ~(t[174]);
  assign t[310] = (x[7]);
  assign t[311] = (x[10]);
  assign t[312] = (x[10]);
  assign t[313] = (x[13]);
  assign t[314] = (x[13]);
  assign t[315] = (x[16]);
  assign t[316] = (x[16]);
  assign t[317] = (x[19]);
  assign t[318] = (x[19]);
  assign t[319] = (x[22]);
  assign t[31] = ~(t[175]);
  assign t[320] = (x[22]);
  assign t[321] = (x[25]);
  assign t[322] = (x[25]);
  assign t[323] = (x[28]);
  assign t[324] = (x[28]);
  assign t[325] = (x[31]);
  assign t[326] = (x[31]);
  assign t[327] = (x[34]);
  assign t[328] = (x[34]);
  assign t[329] = (x[37]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[37]);
  assign t[331] = (x[40]);
  assign t[332] = (x[40]);
  assign t[333] = (x[43]);
  assign t[334] = (x[43]);
  assign t[335] = (x[46]);
  assign t[336] = (x[46]);
  assign t[337] = (x[49]);
  assign t[338] = (x[49]);
  assign t[339] = (x[62]);
  assign t[33] = t[53] ? t[54] : t[176];
  assign t[340] = (x[62]);
  assign t[341] = (x[65]);
  assign t[342] = (x[65]);
  assign t[343] = (x[68]);
  assign t[344] = (x[68]);
  assign t[345] = (x[73]);
  assign t[346] = (x[73]);
  assign t[347] = (x[78]);
  assign t[348] = (x[78]);
  assign t[349] = (x[81]);
  assign t[34] = t[53] ? t[55] : t[177];
  assign t[350] = (x[81]);
  assign t[351] = (x[84]);
  assign t[352] = (x[84]);
  assign t[353] = (x[87]);
  assign t[354] = (x[87]);
  assign t[355] = (x[94]);
  assign t[356] = (x[94]);
  assign t[357] = (x[99]);
  assign t[358] = (x[99]);
  assign t[359] = (x[106]);
  assign t[35] = ~(t[56]);
  assign t[360] = (x[106]);
  assign t[36] = t[53] ? t[57] : t[178];
  assign t[37] = t[27] ? t[58] : t[179];
  assign t[38] = t[27] ? t[59] : t[180];
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[62] & t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[25];
  assign t[44] = t[46] ^ t[69];
  assign t[45] = t[53] ? t[70] : t[181];
  assign t[46] = t[71] ^ t[72];
  assign t[47] = t[73] & t[74];
  assign t[48] = ~(t[75] & t[76]);
  assign t[49] = t[182] | t[77];
  assign t[4] = t[8] ? t[9] : t[172];
  assign t[50] = ~(t[78]);
  assign t[51] = ~(t[183]);
  assign t[52] = ~(t[79] & t[184]);
  assign t[53] = ~(t[15]);
  assign t[54] = t[176] ^ t[80];
  assign t[55] = t[177] ^ t[81];
  assign t[56] = t[53] ? t[82] : t[185];
  assign t[57] = t[178] ^ t[83];
  assign t[58] = t[179] ^ t[84];
  assign t[59] = t[180] ^ t[85];
  assign t[5] = ~(t[10]);
  assign t[60] = t[86] & t[87];
  assign t[61] = t[88] & t[89];
  assign t[62] = ~(t[60] ^ t[90]);
  assign t[63] = t[91] ^ t[92];
  assign t[64] = t[93] ^ t[94];
  assign t[65] = t[38] ^ t[95];
  assign t[66] = t[96] ^ t[97];
  assign t[67] = t[98] & t[99];
  assign t[68] = ~t[100];
  assign t[69] = t[101] & t[102];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[181] ^ t[103];
  assign t[71] = t[104] & t[105];
  assign t[72] = t[106] & t[107];
  assign t[73] = ~(t[108] ^ t[46]);
  assign t[74] = t[43] ^ t[107];
  assign t[75] = ~(t[77] & t[109]);
  assign t[76] = ~(t[186] ^ t[110]);
  assign t[77] = ~(t[111] & t[112]);
  assign t[78] = ~(t[49]);
  assign t[79] = ~(t[187]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[113] ? x[53] : x[52];
  assign t[81] = t[113] ? x[55] : x[54];
  assign t[82] = t[185] ^ t[114];
  assign t[83] = t[113] ? x[57] : x[56];
  assign t[84] = t[115] ? x[59] : x[58];
  assign t[85] = t[78] ? x[61] : x[60];
  assign t[86] = ~(t[92]);
  assign t[87] = ~(t[116]);
  assign t[88] = ~(t[37]);
  assign t[89] = t[27] ? t[117] : t[188];
  assign t[8] = ~(t[15]);
  assign t[90] = t[21] ^ t[116];
  assign t[91] = t[116] ^ t[38];
  assign t[92] = t[89] ^ t[37];
  assign t[93] = t[56] ^ t[34];
  assign t[94] = t[118] ^ t[119];
  assign t[95] = t[39] ^ t[120];
  assign t[96] = t[8] ? t[121] : t[189];
  assign t[97] = t[173] ^ t[122];
  assign t[98] = ~(t[66] ^ t[123]);
  assign t[99] = t[124] ^ t[125];
  assign t[9] = t[172] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [116:0] x;
 output y;

 wire [360:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[53] ? t[126] : t[190];
  assign t[101] = ~(t[71] ^ t[127]);
  assign t[102] = t[128] ^ t[129];
  assign t[103] = t[113] ? x[72] : x[71];
  assign t[104] = ~(t[129]);
  assign t[105] = ~(t[130]);
  assign t[106] = ~(t[68]);
  assign t[107] = t[131];
  assign t[108] = t[130] ^ t[68];
  assign t[109] = ~(t[132] & t[133]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[134] ^ t[191];
  assign t[111] = ~(t[186]);
  assign t[112] = t[135] & t[134];
  assign t[113] = ~(t[50]);
  assign t[114] = t[113] ? x[77] : x[76];
  assign t[115] = ~(t[50]);
  assign t[116] = t[27] ? t[136] : t[192];
  assign t[117] = t[188] ^ t[137];
  assign t[118] = t[138] ^ t[20];
  assign t[119] = t[139] & t[140];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[141] & t[142];
  assign t[121] = t[189] ^ t[143];
  assign t[122] = t[8] ? t[144] : t[193];
  assign t[123] = t[145] ^ t[146];
  assign t[124] = t[97] ^ t[147];
  assign t[125] = t[174] ^ t[148];
  assign t[126] = t[190] ^ t[149];
  assign t[127] = t[43] ^ t[130];
  assign t[128] = t[130] ^ t[25];
  assign t[129] = t[107] ^ t[68];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[150];
  assign t[131] = t[27] ? t[151] : t[194];
  assign t[132] = ~(t[135] | t[134]);
  assign t[133] = ~(t[152] | t[111]);
  assign t[134] = ~(t[195]);
  assign t[135] = ~(t[191]);
  assign t[136] = t[192] ^ t[153];
  assign t[137] = t[78] ? x[91] : x[90];
  assign t[138] = t[154] & t[155];
  assign t[139] = ~(t[138] ^ t[156]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[19] ^ t[157];
  assign t[141] = ~(t[158] ^ t[39]);
  assign t[142] = t[21] ^ t[89];
  assign t[143] = t[28] ? x[93] : x[92];
  assign t[144] = t[193] ^ t[159];
  assign t[145] = t[160] & t[161];
  assign t[146] = t[162] & t[125];
  assign t[147] = t[184] ^ t[163];
  assign t[148] = t[8] ? t[164] : t[196];
  assign t[149] = t[113] ? x[98] : x[97];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[53] ? t[165] : t[197];
  assign t[151] = t[194] ^ t[166];
  assign t[152] = ~(t[182]);
  assign t[153] = t[115] ? x[103] : x[102];
  assign t[154] = ~(t[157]);
  assign t[155] = ~(t[33]);
  assign t[156] = t[93] ^ t[33];
  assign t[157] = t[36] ^ t[56];
  assign t[158] = t[116] ^ t[37];
  assign t[159] = t[28] ? x[105] : x[104];
  assign t[15] = ~(t[27]);
  assign t[160] = ~(t[167]);
  assign t[161] = ~(t[96]);
  assign t[162] = ~(t[97]);
  assign t[163] = t[8] ? t[168] : t[198];
  assign t[164] = t[196] ^ t[169];
  assign t[165] = t[197] ^ t[170];
  assign t[166] = t[113] ? x[110] : x[109];
  assign t[167] = t[125] ^ t[97];
  assign t[168] = t[198] ^ t[171];
  assign t[169] = t[28] ? x[112] : x[111];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[113] ? x[114] : x[113];
  assign t[171] = t[28] ? x[116] : x[115];
  assign t[172] = (t[199]);
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = t[226] ^ x[4];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[9];
  assign t[201] = t[228] ^ x[12];
  assign t[202] = t[229] ^ x[15];
  assign t[203] = t[230] ^ x[18];
  assign t[204] = t[231] ^ x[21];
  assign t[205] = t[232] ^ x[24];
  assign t[206] = t[233] ^ x[27];
  assign t[207] = t[234] ^ x[30];
  assign t[208] = t[235] ^ x[33];
  assign t[209] = t[236] ^ x[36];
  assign t[20] = t[35] & t[36];
  assign t[210] = t[237] ^ x[39];
  assign t[211] = t[238] ^ x[42];
  assign t[212] = t[239] ^ x[45];
  assign t[213] = t[240] ^ x[48];
  assign t[214] = t[241] ^ x[51];
  assign t[215] = t[242] ^ x[64];
  assign t[216] = t[243] ^ x[67];
  assign t[217] = t[244] ^ x[70];
  assign t[218] = t[245] ^ x[75];
  assign t[219] = t[246] ^ x[80];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[83];
  assign t[221] = t[248] ^ x[86];
  assign t[222] = t[249] ^ x[89];
  assign t[223] = t[250] ^ x[96];
  assign t[224] = t[251] ^ x[101];
  assign t[225] = t[252] ^ x[108];
  assign t[226] = (t[253] & ~t[254]);
  assign t[227] = (t[255] & ~t[256]);
  assign t[228] = (t[257] & ~t[258]);
  assign t[229] = (t[259] & ~t[260]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[261] & ~t[262]);
  assign t[231] = (t[263] & ~t[264]);
  assign t[232] = (t[265] & ~t[266]);
  assign t[233] = (t[267] & ~t[268]);
  assign t[234] = (t[269] & ~t[270]);
  assign t[235] = (t[271] & ~t[272]);
  assign t[236] = (t[273] & ~t[274]);
  assign t[237] = (t[275] & ~t[276]);
  assign t[238] = (t[277] & ~t[278]);
  assign t[239] = (t[279] & ~t[280]);
  assign t[23] = ~(t[41] ^ t[42]);
  assign t[240] = (t[281] & ~t[282]);
  assign t[241] = (t[283] & ~t[284]);
  assign t[242] = (t[285] & ~t[286]);
  assign t[243] = (t[287] & ~t[288]);
  assign t[244] = (t[289] & ~t[290]);
  assign t[245] = (t[291] & ~t[292]);
  assign t[246] = (t[293] & ~t[294]);
  assign t[247] = (t[295] & ~t[296]);
  assign t[248] = (t[297] & ~t[298]);
  assign t[249] = (t[299] & ~t[300]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (t[301] & ~t[302]);
  assign t[251] = (t[303] & ~t[304]);
  assign t[252] = (t[305] & ~t[306]);
  assign t[253] = t[307] ^ x[4];
  assign t[254] = t[308] ^ x[3];
  assign t[255] = t[309] ^ x[9];
  assign t[256] = t[310] ^ x[8];
  assign t[257] = t[311] ^ x[12];
  assign t[258] = t[312] ^ x[11];
  assign t[259] = t[313] ^ x[15];
  assign t[25] = ~t[45];
  assign t[260] = t[314] ^ x[14];
  assign t[261] = t[315] ^ x[18];
  assign t[262] = t[316] ^ x[17];
  assign t[263] = t[317] ^ x[21];
  assign t[264] = t[318] ^ x[20];
  assign t[265] = t[319] ^ x[24];
  assign t[266] = t[320] ^ x[23];
  assign t[267] = t[321] ^ x[27];
  assign t[268] = t[322] ^ x[26];
  assign t[269] = t[323] ^ x[30];
  assign t[26] = t[46] ^ t[47];
  assign t[270] = t[324] ^ x[29];
  assign t[271] = t[325] ^ x[33];
  assign t[272] = t[326] ^ x[32];
  assign t[273] = t[327] ^ x[36];
  assign t[274] = t[328] ^ x[35];
  assign t[275] = t[329] ^ x[39];
  assign t[276] = t[330] ^ x[38];
  assign t[277] = t[331] ^ x[42];
  assign t[278] = t[332] ^ x[41];
  assign t[279] = t[333] ^ x[45];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[44];
  assign t[281] = t[335] ^ x[48];
  assign t[282] = t[336] ^ x[47];
  assign t[283] = t[337] ^ x[51];
  assign t[284] = t[338] ^ x[50];
  assign t[285] = t[339] ^ x[64];
  assign t[286] = t[340] ^ x[63];
  assign t[287] = t[341] ^ x[67];
  assign t[288] = t[342] ^ x[66];
  assign t[289] = t[343] ^ x[70];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[69];
  assign t[291] = t[345] ^ x[75];
  assign t[292] = t[346] ^ x[74];
  assign t[293] = t[347] ^ x[80];
  assign t[294] = t[348] ^ x[79];
  assign t[295] = t[349] ^ x[83];
  assign t[296] = t[350] ^ x[82];
  assign t[297] = t[351] ^ x[86];
  assign t[298] = t[352] ^ x[85];
  assign t[299] = t[353] ^ x[89];
  assign t[29] = ~(t[173]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[88];
  assign t[301] = t[355] ^ x[96];
  assign t[302] = t[356] ^ x[95];
  assign t[303] = t[357] ^ x[101];
  assign t[304] = t[358] ^ x[100];
  assign t[305] = t[359] ^ x[108];
  assign t[306] = t[360] ^ x[107];
  assign t[307] = (x[2]);
  assign t[308] = (x[2]);
  assign t[309] = (x[7]);
  assign t[30] = ~(t[174]);
  assign t[310] = (x[7]);
  assign t[311] = (x[10]);
  assign t[312] = (x[10]);
  assign t[313] = (x[13]);
  assign t[314] = (x[13]);
  assign t[315] = (x[16]);
  assign t[316] = (x[16]);
  assign t[317] = (x[19]);
  assign t[318] = (x[19]);
  assign t[319] = (x[22]);
  assign t[31] = ~(t[175]);
  assign t[320] = (x[22]);
  assign t[321] = (x[25]);
  assign t[322] = (x[25]);
  assign t[323] = (x[28]);
  assign t[324] = (x[28]);
  assign t[325] = (x[31]);
  assign t[326] = (x[31]);
  assign t[327] = (x[34]);
  assign t[328] = (x[34]);
  assign t[329] = (x[37]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[37]);
  assign t[331] = (x[40]);
  assign t[332] = (x[40]);
  assign t[333] = (x[43]);
  assign t[334] = (x[43]);
  assign t[335] = (x[46]);
  assign t[336] = (x[46]);
  assign t[337] = (x[49]);
  assign t[338] = (x[49]);
  assign t[339] = (x[62]);
  assign t[33] = t[53] ? t[54] : t[176];
  assign t[340] = (x[62]);
  assign t[341] = (x[65]);
  assign t[342] = (x[65]);
  assign t[343] = (x[68]);
  assign t[344] = (x[68]);
  assign t[345] = (x[73]);
  assign t[346] = (x[73]);
  assign t[347] = (x[78]);
  assign t[348] = (x[78]);
  assign t[349] = (x[81]);
  assign t[34] = t[53] ? t[55] : t[177];
  assign t[350] = (x[81]);
  assign t[351] = (x[84]);
  assign t[352] = (x[84]);
  assign t[353] = (x[87]);
  assign t[354] = (x[87]);
  assign t[355] = (x[94]);
  assign t[356] = (x[94]);
  assign t[357] = (x[99]);
  assign t[358] = (x[99]);
  assign t[359] = (x[106]);
  assign t[35] = ~(t[56]);
  assign t[360] = (x[106]);
  assign t[36] = t[53] ? t[57] : t[178];
  assign t[37] = t[27] ? t[58] : t[179];
  assign t[38] = t[27] ? t[59] : t[180];
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[62] & t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[25];
  assign t[44] = t[46] ^ t[69];
  assign t[45] = t[53] ? t[70] : t[181];
  assign t[46] = t[71] ^ t[72];
  assign t[47] = t[73] & t[74];
  assign t[48] = ~(t[75] & t[76]);
  assign t[49] = t[182] | t[77];
  assign t[4] = t[8] ? t[9] : t[172];
  assign t[50] = ~(t[78]);
  assign t[51] = ~(t[183]);
  assign t[52] = ~(t[79] & t[184]);
  assign t[53] = ~(t[15]);
  assign t[54] = t[176] ^ t[80];
  assign t[55] = t[177] ^ t[81];
  assign t[56] = t[53] ? t[82] : t[185];
  assign t[57] = t[178] ^ t[83];
  assign t[58] = t[179] ^ t[84];
  assign t[59] = t[180] ^ t[85];
  assign t[5] = ~(t[10]);
  assign t[60] = t[86] & t[87];
  assign t[61] = t[88] & t[89];
  assign t[62] = ~(t[60] ^ t[90]);
  assign t[63] = t[91] ^ t[92];
  assign t[64] = t[93] ^ t[94];
  assign t[65] = t[38] ^ t[95];
  assign t[66] = t[96] ^ t[97];
  assign t[67] = t[98] & t[99];
  assign t[68] = ~t[100];
  assign t[69] = t[101] & t[102];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[181] ^ t[103];
  assign t[71] = t[104] & t[105];
  assign t[72] = t[106] & t[107];
  assign t[73] = ~(t[108] ^ t[46]);
  assign t[74] = t[43] ^ t[107];
  assign t[75] = ~(t[77] & t[109]);
  assign t[76] = ~(t[186] ^ t[110]);
  assign t[77] = ~(t[111] & t[112]);
  assign t[78] = ~(t[49]);
  assign t[79] = ~(t[187]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[113] ? x[53] : x[52];
  assign t[81] = t[113] ? x[55] : x[54];
  assign t[82] = t[185] ^ t[114];
  assign t[83] = t[113] ? x[57] : x[56];
  assign t[84] = t[115] ? x[59] : x[58];
  assign t[85] = t[78] ? x[61] : x[60];
  assign t[86] = ~(t[92]);
  assign t[87] = ~(t[116]);
  assign t[88] = ~(t[37]);
  assign t[89] = t[27] ? t[117] : t[188];
  assign t[8] = ~(t[15]);
  assign t[90] = t[21] ^ t[116];
  assign t[91] = t[116] ^ t[38];
  assign t[92] = t[89] ^ t[37];
  assign t[93] = t[56] ^ t[34];
  assign t[94] = t[118] ^ t[119];
  assign t[95] = t[39] ^ t[120];
  assign t[96] = t[8] ? t[121] : t[189];
  assign t[97] = t[173] ^ t[122];
  assign t[98] = ~(t[66] ^ t[123]);
  assign t[99] = t[124] ^ t[125];
  assign t[9] = t[172] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind66(x, y);
 input [116:0] x;
 output y;

 wire [381:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[57] ? t[127] : t[210];
  assign t[101] = t[57] ? t[128] : t[211];
  assign t[102] = ~(t[70] ^ t[129]);
  assign t[103] = t[130] ^ t[131];
  assign t[104] = t[130] ^ t[132];
  assign t[105] = t[133] ^ t[134];
  assign t[106] = t[135] & t[136];
  assign t[107] = t[137] & t[138];
  assign t[108] = t[134] ^ t[139];
  assign t[109] = t[140] ^ t[141];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[142] ^ t[42];
  assign t[111] = t[57] ? t[143] : t[212];
  assign t[112] = t[129] ^ t[71];
  assign t[113] = ~(t[194]);
  assign t[114] = ~(t[54]);
  assign t[115] = t[41] ^ t[63];
  assign t[116] = t[114] ? x[69] : x[68];
  assign t[117] = t[208] ^ t[144];
  assign t[118] = t[114] ? x[71] : x[70];
  assign t[119] = ~(t[145]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = ~(t[142]);
  assign t[121] = ~(t[98]);
  assign t[122] = t[8] ? t[146] : t[213];
  assign t[123] = t[142] ^ t[98];
  assign t[124] = t[209] ^ t[147];
  assign t[125] = ~(t[94] ^ t[148]);
  assign t[126] = t[110] ^ t[145];
  assign t[127] = t[210] ^ t[149];
  assign t[128] = t[211] ^ t[150];
  assign t[129] = t[151] ^ t[152];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[101] ^ t[111];
  assign t[131] = t[57] ? t[153] : t[214];
  assign t[132] = t[129] ^ t[154];
  assign t[133] = t[155] ? t[156] : t[215];
  assign t[134] = t[196] ^ t[157];
  assign t[135] = ~(t[105] ^ t[140]);
  assign t[136] = t[108] ^ t[158];
  assign t[137] = ~(t[59] ^ t[159]);
  assign t[138] = t[22] ^ t[115];
  assign t[139] = t[203] ^ t[160];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[161] ^ t[162];
  assign t[141] = t[163] & t[164];
  assign t[142] = t[8] ? t[165] : t[216];
  assign t[143] = t[212] ^ t[166];
  assign t[144] = t[114] ? x[85] : x[84];
  assign t[145] = t[122] ^ t[98];
  assign t[146] = t[213] ^ t[167];
  assign t[147] = t[31] ? x[87] : x[86];
  assign t[148] = t[68] ^ t[142];
  assign t[149] = t[114] ? x[89] : x[88];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[114] ? x[91] : x[90];
  assign t[151] = t[168] & t[169];
  assign t[152] = t[170] & t[131];
  assign t[153] = t[214] ^ t[171];
  assign t[154] = t[172] & t[173];
  assign t[155] = ~(t[85]);
  assign t[156] = t[215] ^ t[174];
  assign t[157] = t[155] ? t[175] : t[217];
  assign t[158] = t[197] ^ t[176];
  assign t[159] = t[74] ^ t[39];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[155] ? t[177] : t[218];
  assign t[161] = t[178] & t[179];
  assign t[162] = t[180] & t[158];
  assign t[163] = ~(t[161] ^ t[181]);
  assign t[164] = t[182] ^ t[183];
  assign t[165] = t[216] ^ t[184];
  assign t[166] = t[114] ? x[99] : x[98];
  assign t[167] = t[83] ? x[101] : x[100];
  assign t[168] = ~(t[185]);
  assign t[169] = ~(t[100]);
  assign t[16] = t[194] | t[30];
  assign t[170] = ~(t[101]);
  assign t[171] = t[114] ? x[103] : x[102];
  assign t[172] = ~(t[151] ^ t[186]);
  assign t[173] = t[187] ^ t[185];
  assign t[174] = t[188] ? x[105] : x[104];
  assign t[175] = t[217] ^ t[189];
  assign t[176] = t[155] ? t[190] : t[219];
  assign t[177] = t[218] ^ t[191];
  assign t[178] = ~(t[183]);
  assign t[179] = ~(t[133]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = ~(t[134]);
  assign t[181] = t[108] ^ t[133];
  assign t[182] = t[133] ^ t[139];
  assign t[183] = t[158] ^ t[134];
  assign t[184] = t[31] ? x[110] : x[109];
  assign t[185] = t[131] ^ t[101];
  assign t[186] = t[130] ^ t[100];
  assign t[187] = t[100] ^ t[111];
  assign t[188] = ~(t[54]);
  assign t[189] = t[188] ? x[112] : x[111];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[219] ^ t[192];
  assign t[191] = t[188] ? x[114] : x[113];
  assign t[192] = t[188] ? x[116] : x[115];
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = ~t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[4];
  assign t[221] = t[248] ^ x[7];
  assign t[222] = t[249] ^ x[12];
  assign t[223] = t[250] ^ x[15];
  assign t[224] = t[251] ^ x[18];
  assign t[225] = t[252] ^ x[21];
  assign t[226] = t[253] ^ x[24];
  assign t[227] = t[254] ^ x[27];
  assign t[228] = t[255] ^ x[30];
  assign t[229] = t[256] ^ x[33];
  assign t[22] = t[39] ^ t[20];
  assign t[230] = t[257] ^ x[36];
  assign t[231] = t[258] ^ x[39];
  assign t[232] = t[259] ^ x[42];
  assign t[233] = t[260] ^ x[45];
  assign t[234] = t[261] ^ x[48];
  assign t[235] = t[262] ^ x[53];
  assign t[236] = t[263] ^ x[58];
  assign t[237] = t[264] ^ x[61];
  assign t[238] = t[265] ^ x[64];
  assign t[239] = t[266] ^ x[67];
  assign t[23] = t[40] & t[41];
  assign t[240] = t[267] ^ x[74];
  assign t[241] = t[268] ^ x[77];
  assign t[242] = t[269] ^ x[80];
  assign t[243] = t[270] ^ x[83];
  assign t[244] = t[271] ^ x[94];
  assign t[245] = t[272] ^ x[97];
  assign t[246] = t[273] ^ x[108];
  assign t[247] = (t[274] & ~t[275]);
  assign t[248] = (t[276] & ~t[277]);
  assign t[249] = (t[278] & ~t[279]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[280] & ~t[281]);
  assign t[251] = (t[282] & ~t[283]);
  assign t[252] = (t[284] & ~t[285]);
  assign t[253] = (t[286] & ~t[287]);
  assign t[254] = (t[288] & ~t[289]);
  assign t[255] = (t[290] & ~t[291]);
  assign t[256] = (t[292] & ~t[293]);
  assign t[257] = (t[294] & ~t[295]);
  assign t[258] = (t[296] & ~t[297]);
  assign t[259] = (t[298] & ~t[299]);
  assign t[25] = t[44] ^ t[45];
  assign t[260] = (t[300] & ~t[301]);
  assign t[261] = (t[302] & ~t[303]);
  assign t[262] = (t[304] & ~t[305]);
  assign t[263] = (t[306] & ~t[307]);
  assign t[264] = (t[308] & ~t[309]);
  assign t[265] = (t[310] & ~t[311]);
  assign t[266] = (t[312] & ~t[313]);
  assign t[267] = (t[314] & ~t[315]);
  assign t[268] = (t[316] & ~t[317]);
  assign t[269] = (t[318] & ~t[319]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[320] & ~t[321]);
  assign t[271] = (t[322] & ~t[323]);
  assign t[272] = (t[324] & ~t[325]);
  assign t[273] = (t[326] & ~t[327]);
  assign t[274] = t[328] ^ x[4];
  assign t[275] = t[329] ^ x[3];
  assign t[276] = t[330] ^ x[7];
  assign t[277] = t[331] ^ x[6];
  assign t[278] = t[332] ^ x[12];
  assign t[279] = t[333] ^ x[11];
  assign t[27] = ~(t[48] ^ t[49]);
  assign t[280] = t[334] ^ x[15];
  assign t[281] = t[335] ^ x[14];
  assign t[282] = t[336] ^ x[18];
  assign t[283] = t[337] ^ x[17];
  assign t[284] = t[338] ^ x[21];
  assign t[285] = t[339] ^ x[20];
  assign t[286] = t[340] ^ x[24];
  assign t[287] = t[341] ^ x[23];
  assign t[288] = t[342] ^ x[27];
  assign t[289] = t[343] ^ x[26];
  assign t[28] = ~(t[30] & t[50]);
  assign t[290] = t[344] ^ x[30];
  assign t[291] = t[345] ^ x[29];
  assign t[292] = t[346] ^ x[33];
  assign t[293] = t[347] ^ x[32];
  assign t[294] = t[348] ^ x[36];
  assign t[295] = t[349] ^ x[35];
  assign t[296] = t[350] ^ x[39];
  assign t[297] = t[351] ^ x[38];
  assign t[298] = t[352] ^ x[42];
  assign t[299] = t[353] ^ x[41];
  assign t[29] = ~(t[195] ^ t[51]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[45];
  assign t[301] = t[355] ^ x[44];
  assign t[302] = t[356] ^ x[48];
  assign t[303] = t[357] ^ x[47];
  assign t[304] = t[358] ^ x[53];
  assign t[305] = t[359] ^ x[52];
  assign t[306] = t[360] ^ x[58];
  assign t[307] = t[361] ^ x[57];
  assign t[308] = t[362] ^ x[61];
  assign t[309] = t[363] ^ x[60];
  assign t[30] = ~(t[52] & t[53]);
  assign t[310] = t[364] ^ x[64];
  assign t[311] = t[365] ^ x[63];
  assign t[312] = t[366] ^ x[67];
  assign t[313] = t[367] ^ x[66];
  assign t[314] = t[368] ^ x[74];
  assign t[315] = t[369] ^ x[73];
  assign t[316] = t[370] ^ x[77];
  assign t[317] = t[371] ^ x[76];
  assign t[318] = t[372] ^ x[80];
  assign t[319] = t[373] ^ x[79];
  assign t[31] = ~(t[54]);
  assign t[320] = t[374] ^ x[83];
  assign t[321] = t[375] ^ x[82];
  assign t[322] = t[376] ^ x[94];
  assign t[323] = t[377] ^ x[93];
  assign t[324] = t[378] ^ x[97];
  assign t[325] = t[379] ^ x[96];
  assign t[326] = t[380] ^ x[108];
  assign t[327] = t[381] ^ x[107];
  assign t[328] = (x[2]);
  assign t[329] = (x[2]);
  assign t[32] = ~(t[196]);
  assign t[330] = (x[5]);
  assign t[331] = (x[5]);
  assign t[332] = (x[10]);
  assign t[333] = (x[10]);
  assign t[334] = (x[13]);
  assign t[335] = (x[13]);
  assign t[336] = (x[16]);
  assign t[337] = (x[16]);
  assign t[338] = (x[19]);
  assign t[339] = (x[19]);
  assign t[33] = ~(t[197]);
  assign t[340] = (x[22]);
  assign t[341] = (x[22]);
  assign t[342] = (x[25]);
  assign t[343] = (x[25]);
  assign t[344] = (x[28]);
  assign t[345] = (x[28]);
  assign t[346] = (x[31]);
  assign t[347] = (x[31]);
  assign t[348] = (x[34]);
  assign t[349] = (x[34]);
  assign t[34] = ~(t[198]);
  assign t[350] = (x[37]);
  assign t[351] = (x[37]);
  assign t[352] = (x[40]);
  assign t[353] = (x[40]);
  assign t[354] = (x[43]);
  assign t[355] = (x[43]);
  assign t[356] = (x[46]);
  assign t[357] = (x[46]);
  assign t[358] = (x[51]);
  assign t[359] = (x[51]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[56]);
  assign t[361] = (x[56]);
  assign t[362] = (x[59]);
  assign t[363] = (x[59]);
  assign t[364] = (x[62]);
  assign t[365] = (x[62]);
  assign t[366] = (x[65]);
  assign t[367] = (x[65]);
  assign t[368] = (x[72]);
  assign t[369] = (x[72]);
  assign t[36] = t[57] ? t[58] : t[199];
  assign t[370] = (x[75]);
  assign t[371] = (x[75]);
  assign t[372] = (x[78]);
  assign t[373] = (x[78]);
  assign t[374] = (x[81]);
  assign t[375] = (x[81]);
  assign t[376] = (x[92]);
  assign t[377] = (x[92]);
  assign t[378] = (x[95]);
  assign t[379] = (x[95]);
  assign t[37] = t[59] ^ t[23];
  assign t[380] = (x[106]);
  assign t[381] = (x[106]);
  assign t[38] = t[60] & t[61];
  assign t[39] = t[62];
  assign t[3] = t[6] ^ t[7];
  assign t[40] = ~(t[63]);
  assign t[41] = t[64];
  assign t[42] = t[8] ? t[65] : t[200];
  assign t[43] = t[66] ^ t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] ^ t[73]);
  assign t[47] = t[74] ^ t[75];
  assign t[48] = t[76] ^ t[77];
  assign t[49] = ~(t[11] ^ t[78]);
  assign t[4] = t[8] ? t[9] : t[193];
  assign t[50] = ~(t[79] & t[80]);
  assign t[51] = t[81] ^ t[201];
  assign t[52] = ~(t[195]);
  assign t[53] = t[82] & t[81];
  assign t[54] = ~(t[83]);
  assign t[55] = ~(t[202]);
  assign t[56] = ~(t[84] & t[203]);
  assign t[57] = ~(t[85]);
  assign t[58] = t[199] ^ t[86];
  assign t[59] = t[87] & t[88];
  assign t[5] = ~(t[10]);
  assign t[60] = ~(t[89] ^ t[37]);
  assign t[61] = t[74] ^ t[41];
  assign t[62] = t[57] ? t[90] : t[204];
  assign t[63] = ~t[91];
  assign t[64] = t[8] ? t[92] : t[205];
  assign t[65] = t[200] ^ t[93];
  assign t[66] = t[94] ^ t[95];
  assign t[67] = t[96] & t[97];
  assign t[68] = t[98] ^ t[42];
  assign t[69] = t[66] ^ t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[100] ^ t[101];
  assign t[71] = t[102] & t[103];
  assign t[72] = t[104] ^ t[24];
  assign t[73] = t[105] ^ t[106];
  assign t[74] = t[63] ^ t[20];
  assign t[75] = t[37] ^ t[107];
  assign t[76] = t[108] ^ t[109];
  assign t[77] = t[110] ^ t[95];
  assign t[78] = t[111] ^ t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[113] | t[52]);
  assign t[81] = ~(t[206]);
  assign t[82] = ~(t[201]);
  assign t[83] = ~(t[16]);
  assign t[84] = ~(t[207]);
  assign t[85] = ~(t[8]);
  assign t[86] = t[114] ? x[50] : x[49];
  assign t[87] = ~(t[115]);
  assign t[88] = ~(t[39]);
  assign t[89] = t[39] ^ t[63];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[204] ^ t[116];
  assign t[91] = t[57] ? t[117] : t[208];
  assign t[92] = t[205] ^ t[118];
  assign t[93] = t[83] ? x[55] : x[54];
  assign t[94] = t[119] & t[120];
  assign t[95] = t[121] & t[122];
  assign t[96] = ~(t[123] ^ t[66]);
  assign t[97] = t[68] ^ t[122];
  assign t[98] = t[8] ? t[124] : t[209];
  assign t[99] = t[125] & t[126];
  assign t[9] = t[193] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind67(x, y);
 input [116:0] x;
 output y;

 wire [381:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[57] ? t[127] : t[210];
  assign t[101] = t[57] ? t[128] : t[211];
  assign t[102] = ~(t[70] ^ t[129]);
  assign t[103] = t[130] ^ t[131];
  assign t[104] = t[130] ^ t[132];
  assign t[105] = t[133] ^ t[134];
  assign t[106] = t[135] & t[136];
  assign t[107] = t[137] & t[138];
  assign t[108] = t[134] ^ t[139];
  assign t[109] = t[140] ^ t[141];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[142] ^ t[42];
  assign t[111] = t[57] ? t[143] : t[212];
  assign t[112] = t[129] ^ t[71];
  assign t[113] = ~(t[194]);
  assign t[114] = ~(t[54]);
  assign t[115] = t[41] ^ t[63];
  assign t[116] = t[114] ? x[69] : x[68];
  assign t[117] = t[208] ^ t[144];
  assign t[118] = t[114] ? x[71] : x[70];
  assign t[119] = ~(t[145]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = ~(t[142]);
  assign t[121] = ~(t[98]);
  assign t[122] = t[8] ? t[146] : t[213];
  assign t[123] = t[142] ^ t[98];
  assign t[124] = t[209] ^ t[147];
  assign t[125] = ~(t[94] ^ t[148]);
  assign t[126] = t[110] ^ t[145];
  assign t[127] = t[210] ^ t[149];
  assign t[128] = t[211] ^ t[150];
  assign t[129] = t[151] ^ t[152];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[101] ^ t[111];
  assign t[131] = t[57] ? t[153] : t[214];
  assign t[132] = t[129] ^ t[154];
  assign t[133] = t[155] ? t[156] : t[215];
  assign t[134] = t[196] ^ t[157];
  assign t[135] = ~(t[105] ^ t[140]);
  assign t[136] = t[108] ^ t[158];
  assign t[137] = ~(t[59] ^ t[159]);
  assign t[138] = t[22] ^ t[115];
  assign t[139] = t[203] ^ t[160];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[161] ^ t[162];
  assign t[141] = t[163] & t[164];
  assign t[142] = t[8] ? t[165] : t[216];
  assign t[143] = t[212] ^ t[166];
  assign t[144] = t[114] ? x[85] : x[84];
  assign t[145] = t[122] ^ t[98];
  assign t[146] = t[213] ^ t[167];
  assign t[147] = t[31] ? x[87] : x[86];
  assign t[148] = t[68] ^ t[142];
  assign t[149] = t[114] ? x[89] : x[88];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[114] ? x[91] : x[90];
  assign t[151] = t[168] & t[169];
  assign t[152] = t[170] & t[131];
  assign t[153] = t[214] ^ t[171];
  assign t[154] = t[172] & t[173];
  assign t[155] = ~(t[85]);
  assign t[156] = t[215] ^ t[174];
  assign t[157] = t[155] ? t[175] : t[217];
  assign t[158] = t[197] ^ t[176];
  assign t[159] = t[74] ^ t[39];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[155] ? t[177] : t[218];
  assign t[161] = t[178] & t[179];
  assign t[162] = t[180] & t[158];
  assign t[163] = ~(t[161] ^ t[181]);
  assign t[164] = t[182] ^ t[183];
  assign t[165] = t[216] ^ t[184];
  assign t[166] = t[114] ? x[99] : x[98];
  assign t[167] = t[83] ? x[101] : x[100];
  assign t[168] = ~(t[185]);
  assign t[169] = ~(t[100]);
  assign t[16] = t[194] | t[30];
  assign t[170] = ~(t[101]);
  assign t[171] = t[114] ? x[103] : x[102];
  assign t[172] = ~(t[151] ^ t[186]);
  assign t[173] = t[187] ^ t[185];
  assign t[174] = t[188] ? x[105] : x[104];
  assign t[175] = t[217] ^ t[189];
  assign t[176] = t[155] ? t[190] : t[219];
  assign t[177] = t[218] ^ t[191];
  assign t[178] = ~(t[183]);
  assign t[179] = ~(t[133]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = ~(t[134]);
  assign t[181] = t[108] ^ t[133];
  assign t[182] = t[133] ^ t[139];
  assign t[183] = t[158] ^ t[134];
  assign t[184] = t[31] ? x[110] : x[109];
  assign t[185] = t[131] ^ t[101];
  assign t[186] = t[130] ^ t[100];
  assign t[187] = t[100] ^ t[111];
  assign t[188] = ~(t[54]);
  assign t[189] = t[188] ? x[112] : x[111];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[219] ^ t[192];
  assign t[191] = t[188] ? x[114] : x[113];
  assign t[192] = t[188] ? x[116] : x[115];
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = ~t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[4];
  assign t[221] = t[248] ^ x[7];
  assign t[222] = t[249] ^ x[12];
  assign t[223] = t[250] ^ x[15];
  assign t[224] = t[251] ^ x[18];
  assign t[225] = t[252] ^ x[21];
  assign t[226] = t[253] ^ x[24];
  assign t[227] = t[254] ^ x[27];
  assign t[228] = t[255] ^ x[30];
  assign t[229] = t[256] ^ x[33];
  assign t[22] = t[39] ^ t[20];
  assign t[230] = t[257] ^ x[36];
  assign t[231] = t[258] ^ x[39];
  assign t[232] = t[259] ^ x[42];
  assign t[233] = t[260] ^ x[45];
  assign t[234] = t[261] ^ x[48];
  assign t[235] = t[262] ^ x[53];
  assign t[236] = t[263] ^ x[58];
  assign t[237] = t[264] ^ x[61];
  assign t[238] = t[265] ^ x[64];
  assign t[239] = t[266] ^ x[67];
  assign t[23] = t[40] & t[41];
  assign t[240] = t[267] ^ x[74];
  assign t[241] = t[268] ^ x[77];
  assign t[242] = t[269] ^ x[80];
  assign t[243] = t[270] ^ x[83];
  assign t[244] = t[271] ^ x[94];
  assign t[245] = t[272] ^ x[97];
  assign t[246] = t[273] ^ x[108];
  assign t[247] = (t[274] & ~t[275]);
  assign t[248] = (t[276] & ~t[277]);
  assign t[249] = (t[278] & ~t[279]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[280] & ~t[281]);
  assign t[251] = (t[282] & ~t[283]);
  assign t[252] = (t[284] & ~t[285]);
  assign t[253] = (t[286] & ~t[287]);
  assign t[254] = (t[288] & ~t[289]);
  assign t[255] = (t[290] & ~t[291]);
  assign t[256] = (t[292] & ~t[293]);
  assign t[257] = (t[294] & ~t[295]);
  assign t[258] = (t[296] & ~t[297]);
  assign t[259] = (t[298] & ~t[299]);
  assign t[25] = t[44] ^ t[45];
  assign t[260] = (t[300] & ~t[301]);
  assign t[261] = (t[302] & ~t[303]);
  assign t[262] = (t[304] & ~t[305]);
  assign t[263] = (t[306] & ~t[307]);
  assign t[264] = (t[308] & ~t[309]);
  assign t[265] = (t[310] & ~t[311]);
  assign t[266] = (t[312] & ~t[313]);
  assign t[267] = (t[314] & ~t[315]);
  assign t[268] = (t[316] & ~t[317]);
  assign t[269] = (t[318] & ~t[319]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[320] & ~t[321]);
  assign t[271] = (t[322] & ~t[323]);
  assign t[272] = (t[324] & ~t[325]);
  assign t[273] = (t[326] & ~t[327]);
  assign t[274] = t[328] ^ x[4];
  assign t[275] = t[329] ^ x[3];
  assign t[276] = t[330] ^ x[7];
  assign t[277] = t[331] ^ x[6];
  assign t[278] = t[332] ^ x[12];
  assign t[279] = t[333] ^ x[11];
  assign t[27] = ~(t[48] ^ t[49]);
  assign t[280] = t[334] ^ x[15];
  assign t[281] = t[335] ^ x[14];
  assign t[282] = t[336] ^ x[18];
  assign t[283] = t[337] ^ x[17];
  assign t[284] = t[338] ^ x[21];
  assign t[285] = t[339] ^ x[20];
  assign t[286] = t[340] ^ x[24];
  assign t[287] = t[341] ^ x[23];
  assign t[288] = t[342] ^ x[27];
  assign t[289] = t[343] ^ x[26];
  assign t[28] = ~(t[30] & t[50]);
  assign t[290] = t[344] ^ x[30];
  assign t[291] = t[345] ^ x[29];
  assign t[292] = t[346] ^ x[33];
  assign t[293] = t[347] ^ x[32];
  assign t[294] = t[348] ^ x[36];
  assign t[295] = t[349] ^ x[35];
  assign t[296] = t[350] ^ x[39];
  assign t[297] = t[351] ^ x[38];
  assign t[298] = t[352] ^ x[42];
  assign t[299] = t[353] ^ x[41];
  assign t[29] = ~(t[195] ^ t[51]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[45];
  assign t[301] = t[355] ^ x[44];
  assign t[302] = t[356] ^ x[48];
  assign t[303] = t[357] ^ x[47];
  assign t[304] = t[358] ^ x[53];
  assign t[305] = t[359] ^ x[52];
  assign t[306] = t[360] ^ x[58];
  assign t[307] = t[361] ^ x[57];
  assign t[308] = t[362] ^ x[61];
  assign t[309] = t[363] ^ x[60];
  assign t[30] = ~(t[52] & t[53]);
  assign t[310] = t[364] ^ x[64];
  assign t[311] = t[365] ^ x[63];
  assign t[312] = t[366] ^ x[67];
  assign t[313] = t[367] ^ x[66];
  assign t[314] = t[368] ^ x[74];
  assign t[315] = t[369] ^ x[73];
  assign t[316] = t[370] ^ x[77];
  assign t[317] = t[371] ^ x[76];
  assign t[318] = t[372] ^ x[80];
  assign t[319] = t[373] ^ x[79];
  assign t[31] = ~(t[54]);
  assign t[320] = t[374] ^ x[83];
  assign t[321] = t[375] ^ x[82];
  assign t[322] = t[376] ^ x[94];
  assign t[323] = t[377] ^ x[93];
  assign t[324] = t[378] ^ x[97];
  assign t[325] = t[379] ^ x[96];
  assign t[326] = t[380] ^ x[108];
  assign t[327] = t[381] ^ x[107];
  assign t[328] = (x[2]);
  assign t[329] = (x[2]);
  assign t[32] = ~(t[196]);
  assign t[330] = (x[5]);
  assign t[331] = (x[5]);
  assign t[332] = (x[10]);
  assign t[333] = (x[10]);
  assign t[334] = (x[13]);
  assign t[335] = (x[13]);
  assign t[336] = (x[16]);
  assign t[337] = (x[16]);
  assign t[338] = (x[19]);
  assign t[339] = (x[19]);
  assign t[33] = ~(t[197]);
  assign t[340] = (x[22]);
  assign t[341] = (x[22]);
  assign t[342] = (x[25]);
  assign t[343] = (x[25]);
  assign t[344] = (x[28]);
  assign t[345] = (x[28]);
  assign t[346] = (x[31]);
  assign t[347] = (x[31]);
  assign t[348] = (x[34]);
  assign t[349] = (x[34]);
  assign t[34] = ~(t[198]);
  assign t[350] = (x[37]);
  assign t[351] = (x[37]);
  assign t[352] = (x[40]);
  assign t[353] = (x[40]);
  assign t[354] = (x[43]);
  assign t[355] = (x[43]);
  assign t[356] = (x[46]);
  assign t[357] = (x[46]);
  assign t[358] = (x[51]);
  assign t[359] = (x[51]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[56]);
  assign t[361] = (x[56]);
  assign t[362] = (x[59]);
  assign t[363] = (x[59]);
  assign t[364] = (x[62]);
  assign t[365] = (x[62]);
  assign t[366] = (x[65]);
  assign t[367] = (x[65]);
  assign t[368] = (x[72]);
  assign t[369] = (x[72]);
  assign t[36] = t[57] ? t[58] : t[199];
  assign t[370] = (x[75]);
  assign t[371] = (x[75]);
  assign t[372] = (x[78]);
  assign t[373] = (x[78]);
  assign t[374] = (x[81]);
  assign t[375] = (x[81]);
  assign t[376] = (x[92]);
  assign t[377] = (x[92]);
  assign t[378] = (x[95]);
  assign t[379] = (x[95]);
  assign t[37] = t[59] ^ t[23];
  assign t[380] = (x[106]);
  assign t[381] = (x[106]);
  assign t[38] = t[60] & t[61];
  assign t[39] = t[62];
  assign t[3] = t[6] ^ t[7];
  assign t[40] = ~(t[63]);
  assign t[41] = t[64];
  assign t[42] = t[8] ? t[65] : t[200];
  assign t[43] = t[66] ^ t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] ^ t[73]);
  assign t[47] = t[74] ^ t[75];
  assign t[48] = t[76] ^ t[77];
  assign t[49] = ~(t[11] ^ t[78]);
  assign t[4] = t[8] ? t[9] : t[193];
  assign t[50] = ~(t[79] & t[80]);
  assign t[51] = t[81] ^ t[201];
  assign t[52] = ~(t[195]);
  assign t[53] = t[82] & t[81];
  assign t[54] = ~(t[83]);
  assign t[55] = ~(t[202]);
  assign t[56] = ~(t[84] & t[203]);
  assign t[57] = ~(t[85]);
  assign t[58] = t[199] ^ t[86];
  assign t[59] = t[87] & t[88];
  assign t[5] = ~(t[10]);
  assign t[60] = ~(t[89] ^ t[37]);
  assign t[61] = t[74] ^ t[41];
  assign t[62] = t[57] ? t[90] : t[204];
  assign t[63] = ~t[91];
  assign t[64] = t[8] ? t[92] : t[205];
  assign t[65] = t[200] ^ t[93];
  assign t[66] = t[94] ^ t[95];
  assign t[67] = t[96] & t[97];
  assign t[68] = t[98] ^ t[42];
  assign t[69] = t[66] ^ t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[100] ^ t[101];
  assign t[71] = t[102] & t[103];
  assign t[72] = t[104] ^ t[24];
  assign t[73] = t[105] ^ t[106];
  assign t[74] = t[63] ^ t[20];
  assign t[75] = t[37] ^ t[107];
  assign t[76] = t[108] ^ t[109];
  assign t[77] = t[110] ^ t[95];
  assign t[78] = t[111] ^ t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[113] | t[52]);
  assign t[81] = ~(t[206]);
  assign t[82] = ~(t[201]);
  assign t[83] = ~(t[16]);
  assign t[84] = ~(t[207]);
  assign t[85] = ~(t[8]);
  assign t[86] = t[114] ? x[50] : x[49];
  assign t[87] = ~(t[115]);
  assign t[88] = ~(t[39]);
  assign t[89] = t[39] ^ t[63];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[204] ^ t[116];
  assign t[91] = t[57] ? t[117] : t[208];
  assign t[92] = t[205] ^ t[118];
  assign t[93] = t[83] ? x[55] : x[54];
  assign t[94] = t[119] & t[120];
  assign t[95] = t[121] & t[122];
  assign t[96] = ~(t[123] ^ t[66]);
  assign t[97] = t[68] ^ t[122];
  assign t[98] = t[8] ? t[124] : t[209];
  assign t[99] = t[125] & t[126];
  assign t[9] = t[193] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind68(x, y);
 input [116:0] x;
 output y;

 wire [370:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[195] ^ t[129];
  assign t[101] = t[31] ? x[72] : x[71];
  assign t[102] = t[196] ^ t[130];
  assign t[103] = t[131] & t[132];
  assign t[104] = ~(t[103] ^ t[133]);
  assign t[105] = t[61] ^ t[134];
  assign t[106] = t[135] & t[136];
  assign t[107] = ~(t[116] ^ t[72]);
  assign t[108] = t[137] ^ t[43];
  assign t[109] = t[197] ^ t[138];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[198] ^ t[139];
  assign t[111] = t[140] & t[141];
  assign t[112] = t[8] ? t[142] : t[203];
  assign t[113] = ~(t[183]);
  assign t[114] = t[95] ? t[143] : t[204];
  assign t[115] = ~(t[48]);
  assign t[116] = t[40] ^ t[67];
  assign t[117] = t[193] ^ t[144];
  assign t[118] = t[120] ^ t[145];
  assign t[119] = t[185] ^ t[146];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[147] ^ t[148];
  assign t[121] = t[149] & t[150];
  assign t[122] = t[201] ^ t[151];
  assign t[123] = t[202] ^ t[152];
  assign t[124] = ~(t[8]);
  assign t[125] = t[153] ? x[80] : x[79];
  assign t[126] = ~(t[154] ^ t[70]);
  assign t[127] = t[44] ^ t[94];
  assign t[128] = ~(t[155]);
  assign t[129] = t[128] ? x[82] : x[81];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[153] ? x[84] : x[83];
  assign t[131] = ~(t[134]);
  assign t[132] = ~(t[92]);
  assign t[133] = t[44] ^ t[92];
  assign t[134] = t[94] ^ t[69];
  assign t[135] = ~(t[156]);
  assign t[136] = ~(t[40]);
  assign t[137] = t[67] ^ t[41];
  assign t[138] = t[153] ? x[86] : x[85];
  assign t[139] = t[153] ? x[88] : x[87];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[157]);
  assign t[141] = ~(t[47]);
  assign t[142] = t[203] ^ t[158];
  assign t[143] = t[204] ^ t[159];
  assign t[144] = t[160] ? t[161] : t[205];
  assign t[145] = t[162] & t[163];
  assign t[146] = t[160] ? t[164] : t[206];
  assign t[147] = t[165] & t[166];
  assign t[148] = t[167] & t[168];
  assign t[149] = ~(t[147] ^ t[169]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[170] ^ t[171];
  assign t[151] = t[153] ? x[96] : x[95];
  assign t[152] = t[153] ? x[98] : x[97];
  assign t[153] = ~(t[155]);
  assign t[154] = t[92] ^ t[69];
  assign t[155] = ~(t[31]);
  assign t[156] = t[43] ^ t[67];
  assign t[157] = t[78] ^ t[48];
  assign t[158] = t[153] ? x[100] : x[99];
  assign t[159] = t[153] ? x[102] : x[101];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = ~(t[124]);
  assign t[161] = t[205] ^ t[172];
  assign t[162] = ~(t[173] ^ t[120]);
  assign t[163] = t[90] ^ t[168];
  assign t[164] = t[206] ^ t[174];
  assign t[165] = ~(t[171]);
  assign t[166] = ~(t[175]);
  assign t[167] = ~(t[119]);
  assign t[168] = t[186] ^ t[176];
  assign t[169] = t[90] ^ t[175];
  assign t[16] = t[183] | t[30];
  assign t[170] = t[175] ^ t[117];
  assign t[171] = t[168] ^ t[119];
  assign t[172] = t[177] ? x[104] : x[103];
  assign t[173] = t[175] ^ t[119];
  assign t[174] = t[177] ? x[106] : x[105];
  assign t[175] = t[160] ? t[178] : t[207];
  assign t[176] = t[160] ? t[179] : t[208];
  assign t[177] = ~(t[155]);
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[208] ^ t[181];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[177] ? x[114] : x[113];
  assign t[181] = t[177] ? x[116] : x[115];
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = t[236] ^ x[4];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[7];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[60];
  assign t[228] = t[255] ^ x[63];
  assign t[229] = t[256] ^ x[66];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[75];
  assign t[231] = t[258] ^ x[78];
  assign t[232] = t[259] ^ x[91];
  assign t[233] = t[260] ^ x[94];
  assign t[234] = t[261] ^ x[109];
  assign t[235] = t[262] ^ x[112];
  assign t[236] = (t[263] & ~t[264]);
  assign t[237] = (t[265] & ~t[266]);
  assign t[238] = (t[267] & ~t[268]);
  assign t[239] = (t[269] & ~t[270]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[271] & ~t[272]);
  assign t[241] = (t[273] & ~t[274]);
  assign t[242] = (t[275] & ~t[276]);
  assign t[243] = (t[277] & ~t[278]);
  assign t[244] = (t[279] & ~t[280]);
  assign t[245] = (t[281] & ~t[282]);
  assign t[246] = (t[283] & ~t[284]);
  assign t[247] = (t[285] & ~t[286]);
  assign t[248] = (t[287] & ~t[288]);
  assign t[249] = (t[289] & ~t[290]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[291] & ~t[292]);
  assign t[251] = (t[293] & ~t[294]);
  assign t[252] = (t[295] & ~t[296]);
  assign t[253] = (t[297] & ~t[298]);
  assign t[254] = (t[299] & ~t[300]);
  assign t[255] = (t[301] & ~t[302]);
  assign t[256] = (t[303] & ~t[304]);
  assign t[257] = (t[305] & ~t[306]);
  assign t[258] = (t[307] & ~t[308]);
  assign t[259] = (t[309] & ~t[310]);
  assign t[25] = t[41] ^ t[46];
  assign t[260] = (t[311] & ~t[312]);
  assign t[261] = (t[313] & ~t[314]);
  assign t[262] = (t[315] & ~t[316]);
  assign t[263] = t[317] ^ x[4];
  assign t[264] = t[318] ^ x[3];
  assign t[265] = t[319] ^ x[7];
  assign t[266] = t[320] ^ x[6];
  assign t[267] = t[321] ^ x[12];
  assign t[268] = t[322] ^ x[11];
  assign t[269] = t[323] ^ x[15];
  assign t[26] = t[47] ^ t[48];
  assign t[270] = t[324] ^ x[14];
  assign t[271] = t[325] ^ x[18];
  assign t[272] = t[326] ^ x[17];
  assign t[273] = t[327] ^ x[21];
  assign t[274] = t[328] ^ x[20];
  assign t[275] = t[329] ^ x[24];
  assign t[276] = t[330] ^ x[23];
  assign t[277] = t[331] ^ x[27];
  assign t[278] = t[332] ^ x[26];
  assign t[279] = t[333] ^ x[30];
  assign t[27] = t[49] & t[50];
  assign t[280] = t[334] ^ x[29];
  assign t[281] = t[335] ^ x[33];
  assign t[282] = t[336] ^ x[32];
  assign t[283] = t[337] ^ x[36];
  assign t[284] = t[338] ^ x[35];
  assign t[285] = t[339] ^ x[39];
  assign t[286] = t[340] ^ x[38];
  assign t[287] = t[341] ^ x[42];
  assign t[288] = t[342] ^ x[41];
  assign t[289] = t[343] ^ x[45];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[44];
  assign t[291] = t[345] ^ x[48];
  assign t[292] = t[346] ^ x[47];
  assign t[293] = t[347] ^ x[51];
  assign t[294] = t[348] ^ x[50];
  assign t[295] = t[349] ^ x[54];
  assign t[296] = t[350] ^ x[53];
  assign t[297] = t[351] ^ x[57];
  assign t[298] = t[352] ^ x[56];
  assign t[299] = t[353] ^ x[60];
  assign t[29] = ~(t[184] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[59];
  assign t[301] = t[355] ^ x[63];
  assign t[302] = t[356] ^ x[62];
  assign t[303] = t[357] ^ x[66];
  assign t[304] = t[358] ^ x[65];
  assign t[305] = t[359] ^ x[75];
  assign t[306] = t[360] ^ x[74];
  assign t[307] = t[361] ^ x[78];
  assign t[308] = t[362] ^ x[77];
  assign t[309] = t[363] ^ x[91];
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = t[364] ^ x[90];
  assign t[311] = t[365] ^ x[94];
  assign t[312] = t[366] ^ x[93];
  assign t[313] = t[367] ^ x[109];
  assign t[314] = t[368] ^ x[108];
  assign t[315] = t[369] ^ x[112];
  assign t[316] = t[370] ^ x[111];
  assign t[317] = (x[2]);
  assign t[318] = (x[2]);
  assign t[319] = (x[5]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[5]);
  assign t[321] = (x[10]);
  assign t[322] = (x[10]);
  assign t[323] = (x[13]);
  assign t[324] = (x[13]);
  assign t[325] = (x[16]);
  assign t[326] = (x[16]);
  assign t[327] = (x[19]);
  assign t[328] = (x[19]);
  assign t[329] = (x[22]);
  assign t[32] = ~(t[185]);
  assign t[330] = (x[22]);
  assign t[331] = (x[25]);
  assign t[332] = (x[25]);
  assign t[333] = (x[28]);
  assign t[334] = (x[28]);
  assign t[335] = (x[31]);
  assign t[336] = (x[31]);
  assign t[337] = (x[34]);
  assign t[338] = (x[34]);
  assign t[339] = (x[37]);
  assign t[33] = ~(t[186]);
  assign t[340] = (x[37]);
  assign t[341] = (x[40]);
  assign t[342] = (x[40]);
  assign t[343] = (x[43]);
  assign t[344] = (x[43]);
  assign t[345] = (x[46]);
  assign t[346] = (x[46]);
  assign t[347] = (x[49]);
  assign t[348] = (x[49]);
  assign t[349] = (x[52]);
  assign t[34] = ~(t[187]);
  assign t[350] = (x[52]);
  assign t[351] = (x[55]);
  assign t[352] = (x[55]);
  assign t[353] = (x[58]);
  assign t[354] = (x[58]);
  assign t[355] = (x[61]);
  assign t[356] = (x[61]);
  assign t[357] = (x[64]);
  assign t[358] = (x[64]);
  assign t[359] = (x[73]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[73]);
  assign t[361] = (x[76]);
  assign t[362] = (x[76]);
  assign t[363] = (x[89]);
  assign t[364] = (x[89]);
  assign t[365] = (x[92]);
  assign t[366] = (x[92]);
  assign t[367] = (x[107]);
  assign t[368] = (x[107]);
  assign t[369] = (x[110]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[110]);
  assign t[37] = ~(t[59] ^ t[60]);
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[64];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[65] : t[188];
  assign t[41] = t[8] ? t[66] : t[189];
  assign t[42] = ~(t[67]);
  assign t[43] = t[8] ? t[68] : t[190];
  assign t[44] = t[69] ^ t[63];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] ^ t[73];
  assign t[47] = t[74];
  assign t[48] = ~t[75];
  assign t[49] = ~(t[26] ^ t[76]);
  assign t[4] = t[8] ? t[9] : t[182];
  assign t[50] = t[77] ^ t[78];
  assign t[51] = ~(t[79] & t[80]);
  assign t[52] = t[81] ^ t[191];
  assign t[53] = ~(t[184]);
  assign t[54] = t[82] & t[81];
  assign t[55] = ~(t[192]);
  assign t[56] = ~(t[83] & t[193]);
  assign t[57] = t[84] ^ t[85];
  assign t[58] = t[86] ^ t[87];
  assign t[59] = ~(t[88] ^ t[89]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92] ^ t[63];
  assign t[62] = t[93] & t[94];
  assign t[63] = t[95] ? t[96] : t[194];
  assign t[64] = t[70] ^ t[97];
  assign t[65] = t[188] ^ t[98];
  assign t[66] = t[189] ^ t[99];
  assign t[67] = t[8] ? t[100] : t[195];
  assign t[68] = t[190] ^ t[101];
  assign t[69] = t[95] ? t[102] : t[196];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[103] ^ t[62];
  assign t[71] = t[104] & t[105];
  assign t[72] = t[106] ^ t[23];
  assign t[73] = t[107] & t[108];
  assign t[74] = t[95] ? t[109] : t[197];
  assign t[75] = t[95] ? t[110] : t[198];
  assign t[76] = t[111] ^ t[87];
  assign t[77] = t[48] ^ t[84];
  assign t[78] = t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[113] | t[53]);
  assign t[81] = ~(t[199]);
  assign t[82] = ~(t[191]);
  assign t[83] = ~(t[200]);
  assign t[84] = ~t[114];
  assign t[85] = t[76] ^ t[27];
  assign t[86] = t[47] ^ t[84];
  assign t[87] = t[115] & t[78];
  assign t[88] = t[116] ^ t[73];
  assign t[89] = t[117] ^ t[118];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[119] ^ t[117];
  assign t[91] = t[120] ^ t[121];
  assign t[92] = t[95] ? t[122] : t[201];
  assign t[93] = ~(t[69]);
  assign t[94] = t[95] ? t[123] : t[202];
  assign t[95] = ~(t[124]);
  assign t[96] = t[194] ^ t[125];
  assign t[97] = t[126] & t[127];
  assign t[98] = t[128] ? x[68] : x[67];
  assign t[99] = t[31] ? x[70] : x[69];
  assign t[9] = t[182] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind69(x, y);
 input [116:0] x;
 output y;

 wire [370:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[195] ^ t[129];
  assign t[101] = t[31] ? x[72] : x[71];
  assign t[102] = t[196] ^ t[130];
  assign t[103] = t[131] & t[132];
  assign t[104] = ~(t[103] ^ t[133]);
  assign t[105] = t[61] ^ t[134];
  assign t[106] = t[135] & t[136];
  assign t[107] = ~(t[116] ^ t[72]);
  assign t[108] = t[137] ^ t[43];
  assign t[109] = t[197] ^ t[138];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[198] ^ t[139];
  assign t[111] = t[140] & t[141];
  assign t[112] = t[8] ? t[142] : t[203];
  assign t[113] = ~(t[183]);
  assign t[114] = t[95] ? t[143] : t[204];
  assign t[115] = ~(t[48]);
  assign t[116] = t[40] ^ t[67];
  assign t[117] = t[193] ^ t[144];
  assign t[118] = t[120] ^ t[145];
  assign t[119] = t[185] ^ t[146];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[147] ^ t[148];
  assign t[121] = t[149] & t[150];
  assign t[122] = t[201] ^ t[151];
  assign t[123] = t[202] ^ t[152];
  assign t[124] = ~(t[8]);
  assign t[125] = t[153] ? x[80] : x[79];
  assign t[126] = ~(t[154] ^ t[70]);
  assign t[127] = t[44] ^ t[94];
  assign t[128] = ~(t[155]);
  assign t[129] = t[128] ? x[82] : x[81];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[153] ? x[84] : x[83];
  assign t[131] = ~(t[134]);
  assign t[132] = ~(t[92]);
  assign t[133] = t[44] ^ t[92];
  assign t[134] = t[94] ^ t[69];
  assign t[135] = ~(t[156]);
  assign t[136] = ~(t[40]);
  assign t[137] = t[67] ^ t[41];
  assign t[138] = t[153] ? x[86] : x[85];
  assign t[139] = t[153] ? x[88] : x[87];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[157]);
  assign t[141] = ~(t[47]);
  assign t[142] = t[203] ^ t[158];
  assign t[143] = t[204] ^ t[159];
  assign t[144] = t[160] ? t[161] : t[205];
  assign t[145] = t[162] & t[163];
  assign t[146] = t[160] ? t[164] : t[206];
  assign t[147] = t[165] & t[166];
  assign t[148] = t[167] & t[168];
  assign t[149] = ~(t[147] ^ t[169]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[170] ^ t[171];
  assign t[151] = t[153] ? x[96] : x[95];
  assign t[152] = t[153] ? x[98] : x[97];
  assign t[153] = ~(t[155]);
  assign t[154] = t[92] ^ t[69];
  assign t[155] = ~(t[31]);
  assign t[156] = t[43] ^ t[67];
  assign t[157] = t[78] ^ t[48];
  assign t[158] = t[153] ? x[100] : x[99];
  assign t[159] = t[153] ? x[102] : x[101];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = ~(t[124]);
  assign t[161] = t[205] ^ t[172];
  assign t[162] = ~(t[173] ^ t[120]);
  assign t[163] = t[90] ^ t[168];
  assign t[164] = t[206] ^ t[174];
  assign t[165] = ~(t[171]);
  assign t[166] = ~(t[175]);
  assign t[167] = ~(t[119]);
  assign t[168] = t[186] ^ t[176];
  assign t[169] = t[90] ^ t[175];
  assign t[16] = t[183] | t[30];
  assign t[170] = t[175] ^ t[117];
  assign t[171] = t[168] ^ t[119];
  assign t[172] = t[177] ? x[104] : x[103];
  assign t[173] = t[175] ^ t[119];
  assign t[174] = t[177] ? x[106] : x[105];
  assign t[175] = t[160] ? t[178] : t[207];
  assign t[176] = t[160] ? t[179] : t[208];
  assign t[177] = ~(t[155]);
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[208] ^ t[181];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[177] ? x[114] : x[113];
  assign t[181] = t[177] ? x[116] : x[115];
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = t[236] ^ x[4];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[7];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[60];
  assign t[228] = t[255] ^ x[63];
  assign t[229] = t[256] ^ x[66];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[75];
  assign t[231] = t[258] ^ x[78];
  assign t[232] = t[259] ^ x[91];
  assign t[233] = t[260] ^ x[94];
  assign t[234] = t[261] ^ x[109];
  assign t[235] = t[262] ^ x[112];
  assign t[236] = (t[263] & ~t[264]);
  assign t[237] = (t[265] & ~t[266]);
  assign t[238] = (t[267] & ~t[268]);
  assign t[239] = (t[269] & ~t[270]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[271] & ~t[272]);
  assign t[241] = (t[273] & ~t[274]);
  assign t[242] = (t[275] & ~t[276]);
  assign t[243] = (t[277] & ~t[278]);
  assign t[244] = (t[279] & ~t[280]);
  assign t[245] = (t[281] & ~t[282]);
  assign t[246] = (t[283] & ~t[284]);
  assign t[247] = (t[285] & ~t[286]);
  assign t[248] = (t[287] & ~t[288]);
  assign t[249] = (t[289] & ~t[290]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[291] & ~t[292]);
  assign t[251] = (t[293] & ~t[294]);
  assign t[252] = (t[295] & ~t[296]);
  assign t[253] = (t[297] & ~t[298]);
  assign t[254] = (t[299] & ~t[300]);
  assign t[255] = (t[301] & ~t[302]);
  assign t[256] = (t[303] & ~t[304]);
  assign t[257] = (t[305] & ~t[306]);
  assign t[258] = (t[307] & ~t[308]);
  assign t[259] = (t[309] & ~t[310]);
  assign t[25] = t[41] ^ t[46];
  assign t[260] = (t[311] & ~t[312]);
  assign t[261] = (t[313] & ~t[314]);
  assign t[262] = (t[315] & ~t[316]);
  assign t[263] = t[317] ^ x[4];
  assign t[264] = t[318] ^ x[3];
  assign t[265] = t[319] ^ x[7];
  assign t[266] = t[320] ^ x[6];
  assign t[267] = t[321] ^ x[12];
  assign t[268] = t[322] ^ x[11];
  assign t[269] = t[323] ^ x[15];
  assign t[26] = t[47] ^ t[48];
  assign t[270] = t[324] ^ x[14];
  assign t[271] = t[325] ^ x[18];
  assign t[272] = t[326] ^ x[17];
  assign t[273] = t[327] ^ x[21];
  assign t[274] = t[328] ^ x[20];
  assign t[275] = t[329] ^ x[24];
  assign t[276] = t[330] ^ x[23];
  assign t[277] = t[331] ^ x[27];
  assign t[278] = t[332] ^ x[26];
  assign t[279] = t[333] ^ x[30];
  assign t[27] = t[49] & t[50];
  assign t[280] = t[334] ^ x[29];
  assign t[281] = t[335] ^ x[33];
  assign t[282] = t[336] ^ x[32];
  assign t[283] = t[337] ^ x[36];
  assign t[284] = t[338] ^ x[35];
  assign t[285] = t[339] ^ x[39];
  assign t[286] = t[340] ^ x[38];
  assign t[287] = t[341] ^ x[42];
  assign t[288] = t[342] ^ x[41];
  assign t[289] = t[343] ^ x[45];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[44];
  assign t[291] = t[345] ^ x[48];
  assign t[292] = t[346] ^ x[47];
  assign t[293] = t[347] ^ x[51];
  assign t[294] = t[348] ^ x[50];
  assign t[295] = t[349] ^ x[54];
  assign t[296] = t[350] ^ x[53];
  assign t[297] = t[351] ^ x[57];
  assign t[298] = t[352] ^ x[56];
  assign t[299] = t[353] ^ x[60];
  assign t[29] = ~(t[184] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[59];
  assign t[301] = t[355] ^ x[63];
  assign t[302] = t[356] ^ x[62];
  assign t[303] = t[357] ^ x[66];
  assign t[304] = t[358] ^ x[65];
  assign t[305] = t[359] ^ x[75];
  assign t[306] = t[360] ^ x[74];
  assign t[307] = t[361] ^ x[78];
  assign t[308] = t[362] ^ x[77];
  assign t[309] = t[363] ^ x[91];
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = t[364] ^ x[90];
  assign t[311] = t[365] ^ x[94];
  assign t[312] = t[366] ^ x[93];
  assign t[313] = t[367] ^ x[109];
  assign t[314] = t[368] ^ x[108];
  assign t[315] = t[369] ^ x[112];
  assign t[316] = t[370] ^ x[111];
  assign t[317] = (x[2]);
  assign t[318] = (x[2]);
  assign t[319] = (x[5]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[5]);
  assign t[321] = (x[10]);
  assign t[322] = (x[10]);
  assign t[323] = (x[13]);
  assign t[324] = (x[13]);
  assign t[325] = (x[16]);
  assign t[326] = (x[16]);
  assign t[327] = (x[19]);
  assign t[328] = (x[19]);
  assign t[329] = (x[22]);
  assign t[32] = ~(t[185]);
  assign t[330] = (x[22]);
  assign t[331] = (x[25]);
  assign t[332] = (x[25]);
  assign t[333] = (x[28]);
  assign t[334] = (x[28]);
  assign t[335] = (x[31]);
  assign t[336] = (x[31]);
  assign t[337] = (x[34]);
  assign t[338] = (x[34]);
  assign t[339] = (x[37]);
  assign t[33] = ~(t[186]);
  assign t[340] = (x[37]);
  assign t[341] = (x[40]);
  assign t[342] = (x[40]);
  assign t[343] = (x[43]);
  assign t[344] = (x[43]);
  assign t[345] = (x[46]);
  assign t[346] = (x[46]);
  assign t[347] = (x[49]);
  assign t[348] = (x[49]);
  assign t[349] = (x[52]);
  assign t[34] = ~(t[187]);
  assign t[350] = (x[52]);
  assign t[351] = (x[55]);
  assign t[352] = (x[55]);
  assign t[353] = (x[58]);
  assign t[354] = (x[58]);
  assign t[355] = (x[61]);
  assign t[356] = (x[61]);
  assign t[357] = (x[64]);
  assign t[358] = (x[64]);
  assign t[359] = (x[73]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[73]);
  assign t[361] = (x[76]);
  assign t[362] = (x[76]);
  assign t[363] = (x[89]);
  assign t[364] = (x[89]);
  assign t[365] = (x[92]);
  assign t[366] = (x[92]);
  assign t[367] = (x[107]);
  assign t[368] = (x[107]);
  assign t[369] = (x[110]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[110]);
  assign t[37] = ~(t[59] ^ t[60]);
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[64];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[65] : t[188];
  assign t[41] = t[8] ? t[66] : t[189];
  assign t[42] = ~(t[67]);
  assign t[43] = t[8] ? t[68] : t[190];
  assign t[44] = t[69] ^ t[63];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] ^ t[73];
  assign t[47] = t[74];
  assign t[48] = ~t[75];
  assign t[49] = ~(t[26] ^ t[76]);
  assign t[4] = t[8] ? t[9] : t[182];
  assign t[50] = t[77] ^ t[78];
  assign t[51] = ~(t[79] & t[80]);
  assign t[52] = t[81] ^ t[191];
  assign t[53] = ~(t[184]);
  assign t[54] = t[82] & t[81];
  assign t[55] = ~(t[192]);
  assign t[56] = ~(t[83] & t[193]);
  assign t[57] = t[84] ^ t[85];
  assign t[58] = t[86] ^ t[87];
  assign t[59] = ~(t[88] ^ t[89]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92] ^ t[63];
  assign t[62] = t[93] & t[94];
  assign t[63] = t[95] ? t[96] : t[194];
  assign t[64] = t[70] ^ t[97];
  assign t[65] = t[188] ^ t[98];
  assign t[66] = t[189] ^ t[99];
  assign t[67] = t[8] ? t[100] : t[195];
  assign t[68] = t[190] ^ t[101];
  assign t[69] = t[95] ? t[102] : t[196];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[103] ^ t[62];
  assign t[71] = t[104] & t[105];
  assign t[72] = t[106] ^ t[23];
  assign t[73] = t[107] & t[108];
  assign t[74] = t[95] ? t[109] : t[197];
  assign t[75] = t[95] ? t[110] : t[198];
  assign t[76] = t[111] ^ t[87];
  assign t[77] = t[48] ^ t[84];
  assign t[78] = t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[113] | t[53]);
  assign t[81] = ~(t[199]);
  assign t[82] = ~(t[191]);
  assign t[83] = ~(t[200]);
  assign t[84] = ~t[114];
  assign t[85] = t[76] ^ t[27];
  assign t[86] = t[47] ^ t[84];
  assign t[87] = t[115] & t[78];
  assign t[88] = t[116] ^ t[73];
  assign t[89] = t[117] ^ t[118];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[119] ^ t[117];
  assign t[91] = t[120] ^ t[121];
  assign t[92] = t[95] ? t[122] : t[201];
  assign t[93] = ~(t[69]);
  assign t[94] = t[95] ? t[123] : t[202];
  assign t[95] = ~(t[124]);
  assign t[96] = t[194] ^ t[125];
  assign t[97] = t[126] & t[127];
  assign t[98] = t[128] ? x[68] : x[67];
  assign t[99] = t[31] ? x[70] : x[69];
  assign t[9] = t[182] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [116:0] x;
 output y;

 wire [361:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[133] & t[134];
  assign t[101] = t[31] ? x[64] : x[63];
  assign t[102] = t[31] ? x[66] : x[65];
  assign t[103] = t[135] & t[136];
  assign t[104] = t[137] & t[71];
  assign t[105] = t[8] ? t[138] : t[192];
  assign t[106] = t[185] ^ t[139];
  assign t[107] = t[186] ^ t[140];
  assign t[108] = t[187] ^ t[141];
  assign t[109] = ~(t[115]);
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[93]);
  assign t[111] = ~(t[44]);
  assign t[112] = t[142];
  assign t[113] = t[24] ^ t[93];
  assign t[114] = t[93] ^ t[45];
  assign t[115] = t[112] ^ t[44];
  assign t[116] = ~(t[56]);
  assign t[117] = ~(t[143]);
  assign t[118] = ~(t[129]);
  assign t[119] = ~(t[130]);
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[48] ? t[144] : t[193];
  assign t[121] = t[130] ^ t[26];
  assign t[122] = ~(t[174]);
  assign t[123] = ~(t[78]);
  assign t[124] = t[190] ^ t[145];
  assign t[125] = t[177] ^ t[146];
  assign t[126] = t[123] ? t[147] : t[194];
  assign t[127] = t[48] ? t[148] : t[195];
  assign t[128] = t[149] & t[150];
  assign t[129] = t[48] ? t[151] : t[196];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[48] ? t[152] : t[197];
  assign t[131] = t[191] ^ t[153];
  assign t[132] = t[154] & t[155];
  assign t[133] = ~(t[156] ^ t[99]);
  assign t[134] = t[157] ^ t[92];
  assign t[135] = ~(t[158]);
  assign t[136] = ~(t[40]);
  assign t[137] = ~(t[41]);
  assign t[138] = t[192] ^ t[159];
  assign t[139] = t[88] ? x[86] : x[85];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[116] ? x[88] : x[87];
  assign t[141] = t[116] ? x[90] : x[89];
  assign t[142] = t[8] ? t[160] : t[198];
  assign t[143] = t[120] ^ t[130];
  assign t[144] = t[193] ^ t[161];
  assign t[145] = t[162] ? x[95] : x[94];
  assign t[146] = t[123] ? t[163] : t[199];
  assign t[147] = t[194] ^ t[164];
  assign t[148] = t[195] ^ t[165];
  assign t[149] = ~(t[103] ^ t[166]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[167] ^ t[158];
  assign t[151] = t[196] ^ t[168];
  assign t[152] = t[197] ^ t[169];
  assign t[153] = t[162] ? x[100] : x[99];
  assign t[154] = ~(t[170]);
  assign t[155] = ~(t[90]);
  assign t[156] = t[90] ^ t[125];
  assign t[157] = t[125] ^ t[65];
  assign t[158] = t[71] ^ t[41];
  assign t[159] = t[88] ? x[102] : x[101];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[198] ^ t[171];
  assign t[161] = t[116] ? x[104] : x[103];
  assign t[162] = ~(t[56]);
  assign t[163] = t[199] ^ t[172];
  assign t[164] = t[162] ? x[106] : x[105];
  assign t[165] = t[116] ? x[108] : x[107];
  assign t[166] = t[70] ^ t[40];
  assign t[167] = t[40] ^ t[105];
  assign t[168] = t[116] ? x[110] : x[109];
  assign t[169] = t[116] ? x[112] : x[111];
  assign t[16] = t[174] | t[30];
  assign t[170] = t[92] ^ t[125];
  assign t[171] = t[116] ? x[114] : x[113];
  assign t[172] = t[162] ? x[116] : x[115];
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[4];
  assign t[201] = t[228] ^ x[7];
  assign t[202] = t[229] ^ x[12];
  assign t[203] = t[230] ^ x[15];
  assign t[204] = t[231] ^ x[18];
  assign t[205] = t[232] ^ x[21];
  assign t[206] = t[233] ^ x[24];
  assign t[207] = t[234] ^ x[27];
  assign t[208] = t[235] ^ x[30];
  assign t[209] = t[236] ^ x[33];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[36];
  assign t[211] = t[238] ^ x[39];
  assign t[212] = t[239] ^ x[42];
  assign t[213] = t[240] ^ x[45];
  assign t[214] = t[241] ^ x[48];
  assign t[215] = t[242] ^ x[53];
  assign t[216] = t[243] ^ x[56];
  assign t[217] = t[244] ^ x[59];
  assign t[218] = t[245] ^ x[62];
  assign t[219] = t[246] ^ x[69];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[72];
  assign t[221] = t[248] ^ x[75];
  assign t[222] = t[249] ^ x[78];
  assign t[223] = t[250] ^ x[81];
  assign t[224] = t[251] ^ x[84];
  assign t[225] = t[252] ^ x[93];
  assign t[226] = t[253] ^ x[98];
  assign t[227] = (t[254] & ~t[255]);
  assign t[228] = (t[256] & ~t[257]);
  assign t[229] = (t[258] & ~t[259]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[260] & ~t[261]);
  assign t[231] = (t[262] & ~t[263]);
  assign t[232] = (t[264] & ~t[265]);
  assign t[233] = (t[266] & ~t[267]);
  assign t[234] = (t[268] & ~t[269]);
  assign t[235] = (t[270] & ~t[271]);
  assign t[236] = (t[272] & ~t[273]);
  assign t[237] = (t[274] & ~t[275]);
  assign t[238] = (t[276] & ~t[277]);
  assign t[239] = (t[278] & ~t[279]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[280] & ~t[281]);
  assign t[241] = (t[282] & ~t[283]);
  assign t[242] = (t[284] & ~t[285]);
  assign t[243] = (t[286] & ~t[287]);
  assign t[244] = (t[288] & ~t[289]);
  assign t[245] = (t[290] & ~t[291]);
  assign t[246] = (t[292] & ~t[293]);
  assign t[247] = (t[294] & ~t[295]);
  assign t[248] = (t[296] & ~t[297]);
  assign t[249] = (t[298] & ~t[299]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[300] & ~t[301]);
  assign t[251] = (t[302] & ~t[303]);
  assign t[252] = (t[304] & ~t[305]);
  assign t[253] = (t[306] & ~t[307]);
  assign t[254] = t[308] ^ x[4];
  assign t[255] = t[309] ^ x[3];
  assign t[256] = t[310] ^ x[7];
  assign t[257] = t[311] ^ x[6];
  assign t[258] = t[312] ^ x[12];
  assign t[259] = t[313] ^ x[11];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[314] ^ x[15];
  assign t[261] = t[315] ^ x[14];
  assign t[262] = t[316] ^ x[18];
  assign t[263] = t[317] ^ x[17];
  assign t[264] = t[318] ^ x[21];
  assign t[265] = t[319] ^ x[20];
  assign t[266] = t[320] ^ x[24];
  assign t[267] = t[321] ^ x[23];
  assign t[268] = t[322] ^ x[27];
  assign t[269] = t[323] ^ x[26];
  assign t[26] = t[48] ? t[49] : t[175];
  assign t[270] = t[324] ^ x[30];
  assign t[271] = t[325] ^ x[29];
  assign t[272] = t[326] ^ x[33];
  assign t[273] = t[327] ^ x[32];
  assign t[274] = t[328] ^ x[36];
  assign t[275] = t[329] ^ x[35];
  assign t[276] = t[330] ^ x[39];
  assign t[277] = t[331] ^ x[38];
  assign t[278] = t[332] ^ x[42];
  assign t[279] = t[333] ^ x[41];
  assign t[27] = t[50] ^ t[51];
  assign t[280] = t[334] ^ x[45];
  assign t[281] = t[335] ^ x[44];
  assign t[282] = t[336] ^ x[48];
  assign t[283] = t[337] ^ x[47];
  assign t[284] = t[338] ^ x[53];
  assign t[285] = t[339] ^ x[52];
  assign t[286] = t[340] ^ x[56];
  assign t[287] = t[341] ^ x[55];
  assign t[288] = t[342] ^ x[59];
  assign t[289] = t[343] ^ x[58];
  assign t[28] = ~(t[30] & t[52]);
  assign t[290] = t[344] ^ x[62];
  assign t[291] = t[345] ^ x[61];
  assign t[292] = t[346] ^ x[69];
  assign t[293] = t[347] ^ x[68];
  assign t[294] = t[348] ^ x[72];
  assign t[295] = t[349] ^ x[71];
  assign t[296] = t[350] ^ x[75];
  assign t[297] = t[351] ^ x[74];
  assign t[298] = t[352] ^ x[78];
  assign t[299] = t[353] ^ x[77];
  assign t[29] = ~(t[176] ^ t[53]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[81];
  assign t[301] = t[355] ^ x[80];
  assign t[302] = t[356] ^ x[84];
  assign t[303] = t[357] ^ x[83];
  assign t[304] = t[358] ^ x[93];
  assign t[305] = t[359] ^ x[92];
  assign t[306] = t[360] ^ x[98];
  assign t[307] = t[361] ^ x[97];
  assign t[308] = (x[2]);
  assign t[309] = (x[2]);
  assign t[30] = ~(t[54] & t[55]);
  assign t[310] = (x[5]);
  assign t[311] = (x[5]);
  assign t[312] = (x[10]);
  assign t[313] = (x[10]);
  assign t[314] = (x[13]);
  assign t[315] = (x[13]);
  assign t[316] = (x[16]);
  assign t[317] = (x[16]);
  assign t[318] = (x[19]);
  assign t[319] = (x[19]);
  assign t[31] = ~(t[56]);
  assign t[320] = (x[22]);
  assign t[321] = (x[22]);
  assign t[322] = (x[25]);
  assign t[323] = (x[25]);
  assign t[324] = (x[28]);
  assign t[325] = (x[28]);
  assign t[326] = (x[31]);
  assign t[327] = (x[31]);
  assign t[328] = (x[34]);
  assign t[329] = (x[34]);
  assign t[32] = ~(t[177]);
  assign t[330] = (x[37]);
  assign t[331] = (x[37]);
  assign t[332] = (x[40]);
  assign t[333] = (x[40]);
  assign t[334] = (x[43]);
  assign t[335] = (x[43]);
  assign t[336] = (x[46]);
  assign t[337] = (x[46]);
  assign t[338] = (x[51]);
  assign t[339] = (x[51]);
  assign t[33] = ~(t[178]);
  assign t[340] = (x[54]);
  assign t[341] = (x[54]);
  assign t[342] = (x[57]);
  assign t[343] = (x[57]);
  assign t[344] = (x[60]);
  assign t[345] = (x[60]);
  assign t[346] = (x[67]);
  assign t[347] = (x[67]);
  assign t[348] = (x[70]);
  assign t[349] = (x[70]);
  assign t[34] = ~(t[179]);
  assign t[350] = (x[73]);
  assign t[351] = (x[73]);
  assign t[352] = (x[76]);
  assign t[353] = (x[76]);
  assign t[354] = (x[79]);
  assign t[355] = (x[79]);
  assign t[356] = (x[82]);
  assign t[357] = (x[82]);
  assign t[358] = (x[91]);
  assign t[359] = (x[91]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = (x[96]);
  assign t[361] = (x[96]);
  assign t[36] = t[59] ^ t[60];
  assign t[37] = t[61] ^ t[62];
  assign t[38] = t[63] ^ t[64];
  assign t[39] = t[65] ^ t[66];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[67] : t[180];
  assign t[41] = t[8] ? t[68] : t[181];
  assign t[42] = ~(t[22] ^ t[69]);
  assign t[43] = t[70] ^ t[71];
  assign t[44] = ~t[72];
  assign t[45] = ~t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = t[76] & t[77];
  assign t[48] = ~(t[78]);
  assign t[49] = t[175] ^ t[79];
  assign t[4] = t[8] ? t[9] : t[173];
  assign t[50] = t[80] ^ t[81];
  assign t[51] = t[82] & t[83];
  assign t[52] = ~(t[84] & t[85]);
  assign t[53] = t[86] ^ t[182];
  assign t[54] = ~(t[176]);
  assign t[55] = t[87] & t[86];
  assign t[56] = ~(t[88]);
  assign t[57] = ~(t[183]);
  assign t[58] = ~(t[89] & t[184]);
  assign t[59] = t[90] ^ t[65];
  assign t[5] = ~(t[10]);
  assign t[60] = t[91] & t[92];
  assign t[61] = t[93] ^ t[44];
  assign t[62] = t[94] & t[95];
  assign t[63] = t[70] ^ t[96];
  assign t[64] = t[97] ^ t[51];
  assign t[65] = t[184] ^ t[98];
  assign t[66] = t[99] ^ t[100];
  assign t[67] = t[180] ^ t[101];
  assign t[68] = t[181] ^ t[102];
  assign t[69] = t[103] ^ t[104];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[41] ^ t[105];
  assign t[71] = t[8] ? t[106] : t[185];
  assign t[72] = t[48] ? t[107] : t[186];
  assign t[73] = t[48] ? t[108] : t[187];
  assign t[74] = t[109] & t[110];
  assign t[75] = t[111] & t[112];
  assign t[76] = ~(t[74] ^ t[113]);
  assign t[77] = t[114] ^ t[115];
  assign t[78] = ~(t[8]);
  assign t[79] = t[116] ? x[50] : x[49];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] & t[118];
  assign t[81] = t[119] & t[120];
  assign t[82] = ~(t[97] ^ t[50]);
  assign t[83] = t[121] ^ t[120];
  assign t[84] = ~(t[87] | t[86]);
  assign t[85] = ~(t[122] | t[54]);
  assign t[86] = ~(t[188]);
  assign t[87] = ~(t[182]);
  assign t[88] = ~(t[16]);
  assign t[89] = ~(t[189]);
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[123] ? t[124] : t[190];
  assign t[91] = ~(t[125]);
  assign t[92] = t[178] ^ t[126];
  assign t[93] = t[127];
  assign t[94] = ~(t[61] ^ t[46]);
  assign t[95] = t[24] ^ t[112];
  assign t[96] = t[69] ^ t[128];
  assign t[97] = t[129] ^ t[130];
  assign t[98] = t[123] ? t[131] : t[191];
  assign t[99] = t[132] ^ t[60];
  assign t[9] = t[173] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind71(x, y);
 input [116:0] x;
 output y;

 wire [361:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[133] & t[134];
  assign t[101] = t[31] ? x[64] : x[63];
  assign t[102] = t[31] ? x[66] : x[65];
  assign t[103] = t[135] & t[136];
  assign t[104] = t[137] & t[71];
  assign t[105] = t[8] ? t[138] : t[192];
  assign t[106] = t[185] ^ t[139];
  assign t[107] = t[186] ^ t[140];
  assign t[108] = t[187] ^ t[141];
  assign t[109] = ~(t[115]);
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[93]);
  assign t[111] = ~(t[44]);
  assign t[112] = t[142];
  assign t[113] = t[24] ^ t[93];
  assign t[114] = t[93] ^ t[45];
  assign t[115] = t[112] ^ t[44];
  assign t[116] = ~(t[56]);
  assign t[117] = ~(t[143]);
  assign t[118] = ~(t[129]);
  assign t[119] = ~(t[130]);
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[48] ? t[144] : t[193];
  assign t[121] = t[130] ^ t[26];
  assign t[122] = ~(t[174]);
  assign t[123] = ~(t[78]);
  assign t[124] = t[190] ^ t[145];
  assign t[125] = t[177] ^ t[146];
  assign t[126] = t[123] ? t[147] : t[194];
  assign t[127] = t[48] ? t[148] : t[195];
  assign t[128] = t[149] & t[150];
  assign t[129] = t[48] ? t[151] : t[196];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[48] ? t[152] : t[197];
  assign t[131] = t[191] ^ t[153];
  assign t[132] = t[154] & t[155];
  assign t[133] = ~(t[156] ^ t[99]);
  assign t[134] = t[157] ^ t[92];
  assign t[135] = ~(t[158]);
  assign t[136] = ~(t[40]);
  assign t[137] = ~(t[41]);
  assign t[138] = t[192] ^ t[159];
  assign t[139] = t[88] ? x[86] : x[85];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[116] ? x[88] : x[87];
  assign t[141] = t[116] ? x[90] : x[89];
  assign t[142] = t[8] ? t[160] : t[198];
  assign t[143] = t[120] ^ t[130];
  assign t[144] = t[193] ^ t[161];
  assign t[145] = t[162] ? x[95] : x[94];
  assign t[146] = t[123] ? t[163] : t[199];
  assign t[147] = t[194] ^ t[164];
  assign t[148] = t[195] ^ t[165];
  assign t[149] = ~(t[103] ^ t[166]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[167] ^ t[158];
  assign t[151] = t[196] ^ t[168];
  assign t[152] = t[197] ^ t[169];
  assign t[153] = t[162] ? x[100] : x[99];
  assign t[154] = ~(t[170]);
  assign t[155] = ~(t[90]);
  assign t[156] = t[90] ^ t[125];
  assign t[157] = t[125] ^ t[65];
  assign t[158] = t[71] ^ t[41];
  assign t[159] = t[88] ? x[102] : x[101];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[198] ^ t[171];
  assign t[161] = t[116] ? x[104] : x[103];
  assign t[162] = ~(t[56]);
  assign t[163] = t[199] ^ t[172];
  assign t[164] = t[162] ? x[106] : x[105];
  assign t[165] = t[116] ? x[108] : x[107];
  assign t[166] = t[70] ^ t[40];
  assign t[167] = t[40] ^ t[105];
  assign t[168] = t[116] ? x[110] : x[109];
  assign t[169] = t[116] ? x[112] : x[111];
  assign t[16] = t[174] | t[30];
  assign t[170] = t[92] ^ t[125];
  assign t[171] = t[116] ? x[114] : x[113];
  assign t[172] = t[162] ? x[116] : x[115];
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[4];
  assign t[201] = t[228] ^ x[7];
  assign t[202] = t[229] ^ x[12];
  assign t[203] = t[230] ^ x[15];
  assign t[204] = t[231] ^ x[18];
  assign t[205] = t[232] ^ x[21];
  assign t[206] = t[233] ^ x[24];
  assign t[207] = t[234] ^ x[27];
  assign t[208] = t[235] ^ x[30];
  assign t[209] = t[236] ^ x[33];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[36];
  assign t[211] = t[238] ^ x[39];
  assign t[212] = t[239] ^ x[42];
  assign t[213] = t[240] ^ x[45];
  assign t[214] = t[241] ^ x[48];
  assign t[215] = t[242] ^ x[53];
  assign t[216] = t[243] ^ x[56];
  assign t[217] = t[244] ^ x[59];
  assign t[218] = t[245] ^ x[62];
  assign t[219] = t[246] ^ x[69];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[72];
  assign t[221] = t[248] ^ x[75];
  assign t[222] = t[249] ^ x[78];
  assign t[223] = t[250] ^ x[81];
  assign t[224] = t[251] ^ x[84];
  assign t[225] = t[252] ^ x[93];
  assign t[226] = t[253] ^ x[98];
  assign t[227] = (t[254] & ~t[255]);
  assign t[228] = (t[256] & ~t[257]);
  assign t[229] = (t[258] & ~t[259]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[260] & ~t[261]);
  assign t[231] = (t[262] & ~t[263]);
  assign t[232] = (t[264] & ~t[265]);
  assign t[233] = (t[266] & ~t[267]);
  assign t[234] = (t[268] & ~t[269]);
  assign t[235] = (t[270] & ~t[271]);
  assign t[236] = (t[272] & ~t[273]);
  assign t[237] = (t[274] & ~t[275]);
  assign t[238] = (t[276] & ~t[277]);
  assign t[239] = (t[278] & ~t[279]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[280] & ~t[281]);
  assign t[241] = (t[282] & ~t[283]);
  assign t[242] = (t[284] & ~t[285]);
  assign t[243] = (t[286] & ~t[287]);
  assign t[244] = (t[288] & ~t[289]);
  assign t[245] = (t[290] & ~t[291]);
  assign t[246] = (t[292] & ~t[293]);
  assign t[247] = (t[294] & ~t[295]);
  assign t[248] = (t[296] & ~t[297]);
  assign t[249] = (t[298] & ~t[299]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[300] & ~t[301]);
  assign t[251] = (t[302] & ~t[303]);
  assign t[252] = (t[304] & ~t[305]);
  assign t[253] = (t[306] & ~t[307]);
  assign t[254] = t[308] ^ x[4];
  assign t[255] = t[309] ^ x[3];
  assign t[256] = t[310] ^ x[7];
  assign t[257] = t[311] ^ x[6];
  assign t[258] = t[312] ^ x[12];
  assign t[259] = t[313] ^ x[11];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[314] ^ x[15];
  assign t[261] = t[315] ^ x[14];
  assign t[262] = t[316] ^ x[18];
  assign t[263] = t[317] ^ x[17];
  assign t[264] = t[318] ^ x[21];
  assign t[265] = t[319] ^ x[20];
  assign t[266] = t[320] ^ x[24];
  assign t[267] = t[321] ^ x[23];
  assign t[268] = t[322] ^ x[27];
  assign t[269] = t[323] ^ x[26];
  assign t[26] = t[48] ? t[49] : t[175];
  assign t[270] = t[324] ^ x[30];
  assign t[271] = t[325] ^ x[29];
  assign t[272] = t[326] ^ x[33];
  assign t[273] = t[327] ^ x[32];
  assign t[274] = t[328] ^ x[36];
  assign t[275] = t[329] ^ x[35];
  assign t[276] = t[330] ^ x[39];
  assign t[277] = t[331] ^ x[38];
  assign t[278] = t[332] ^ x[42];
  assign t[279] = t[333] ^ x[41];
  assign t[27] = t[50] ^ t[51];
  assign t[280] = t[334] ^ x[45];
  assign t[281] = t[335] ^ x[44];
  assign t[282] = t[336] ^ x[48];
  assign t[283] = t[337] ^ x[47];
  assign t[284] = t[338] ^ x[53];
  assign t[285] = t[339] ^ x[52];
  assign t[286] = t[340] ^ x[56];
  assign t[287] = t[341] ^ x[55];
  assign t[288] = t[342] ^ x[59];
  assign t[289] = t[343] ^ x[58];
  assign t[28] = ~(t[30] & t[52]);
  assign t[290] = t[344] ^ x[62];
  assign t[291] = t[345] ^ x[61];
  assign t[292] = t[346] ^ x[69];
  assign t[293] = t[347] ^ x[68];
  assign t[294] = t[348] ^ x[72];
  assign t[295] = t[349] ^ x[71];
  assign t[296] = t[350] ^ x[75];
  assign t[297] = t[351] ^ x[74];
  assign t[298] = t[352] ^ x[78];
  assign t[299] = t[353] ^ x[77];
  assign t[29] = ~(t[176] ^ t[53]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[81];
  assign t[301] = t[355] ^ x[80];
  assign t[302] = t[356] ^ x[84];
  assign t[303] = t[357] ^ x[83];
  assign t[304] = t[358] ^ x[93];
  assign t[305] = t[359] ^ x[92];
  assign t[306] = t[360] ^ x[98];
  assign t[307] = t[361] ^ x[97];
  assign t[308] = (x[2]);
  assign t[309] = (x[2]);
  assign t[30] = ~(t[54] & t[55]);
  assign t[310] = (x[5]);
  assign t[311] = (x[5]);
  assign t[312] = (x[10]);
  assign t[313] = (x[10]);
  assign t[314] = (x[13]);
  assign t[315] = (x[13]);
  assign t[316] = (x[16]);
  assign t[317] = (x[16]);
  assign t[318] = (x[19]);
  assign t[319] = (x[19]);
  assign t[31] = ~(t[56]);
  assign t[320] = (x[22]);
  assign t[321] = (x[22]);
  assign t[322] = (x[25]);
  assign t[323] = (x[25]);
  assign t[324] = (x[28]);
  assign t[325] = (x[28]);
  assign t[326] = (x[31]);
  assign t[327] = (x[31]);
  assign t[328] = (x[34]);
  assign t[329] = (x[34]);
  assign t[32] = ~(t[177]);
  assign t[330] = (x[37]);
  assign t[331] = (x[37]);
  assign t[332] = (x[40]);
  assign t[333] = (x[40]);
  assign t[334] = (x[43]);
  assign t[335] = (x[43]);
  assign t[336] = (x[46]);
  assign t[337] = (x[46]);
  assign t[338] = (x[51]);
  assign t[339] = (x[51]);
  assign t[33] = ~(t[178]);
  assign t[340] = (x[54]);
  assign t[341] = (x[54]);
  assign t[342] = (x[57]);
  assign t[343] = (x[57]);
  assign t[344] = (x[60]);
  assign t[345] = (x[60]);
  assign t[346] = (x[67]);
  assign t[347] = (x[67]);
  assign t[348] = (x[70]);
  assign t[349] = (x[70]);
  assign t[34] = ~(t[179]);
  assign t[350] = (x[73]);
  assign t[351] = (x[73]);
  assign t[352] = (x[76]);
  assign t[353] = (x[76]);
  assign t[354] = (x[79]);
  assign t[355] = (x[79]);
  assign t[356] = (x[82]);
  assign t[357] = (x[82]);
  assign t[358] = (x[91]);
  assign t[359] = (x[91]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = (x[96]);
  assign t[361] = (x[96]);
  assign t[36] = t[59] ^ t[60];
  assign t[37] = t[61] ^ t[62];
  assign t[38] = t[63] ^ t[64];
  assign t[39] = t[65] ^ t[66];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[67] : t[180];
  assign t[41] = t[8] ? t[68] : t[181];
  assign t[42] = ~(t[22] ^ t[69]);
  assign t[43] = t[70] ^ t[71];
  assign t[44] = ~t[72];
  assign t[45] = ~t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = t[76] & t[77];
  assign t[48] = ~(t[78]);
  assign t[49] = t[175] ^ t[79];
  assign t[4] = t[8] ? t[9] : t[173];
  assign t[50] = t[80] ^ t[81];
  assign t[51] = t[82] & t[83];
  assign t[52] = ~(t[84] & t[85]);
  assign t[53] = t[86] ^ t[182];
  assign t[54] = ~(t[176]);
  assign t[55] = t[87] & t[86];
  assign t[56] = ~(t[88]);
  assign t[57] = ~(t[183]);
  assign t[58] = ~(t[89] & t[184]);
  assign t[59] = t[90] ^ t[65];
  assign t[5] = ~(t[10]);
  assign t[60] = t[91] & t[92];
  assign t[61] = t[93] ^ t[44];
  assign t[62] = t[94] & t[95];
  assign t[63] = t[70] ^ t[96];
  assign t[64] = t[97] ^ t[51];
  assign t[65] = t[184] ^ t[98];
  assign t[66] = t[99] ^ t[100];
  assign t[67] = t[180] ^ t[101];
  assign t[68] = t[181] ^ t[102];
  assign t[69] = t[103] ^ t[104];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[41] ^ t[105];
  assign t[71] = t[8] ? t[106] : t[185];
  assign t[72] = t[48] ? t[107] : t[186];
  assign t[73] = t[48] ? t[108] : t[187];
  assign t[74] = t[109] & t[110];
  assign t[75] = t[111] & t[112];
  assign t[76] = ~(t[74] ^ t[113]);
  assign t[77] = t[114] ^ t[115];
  assign t[78] = ~(t[8]);
  assign t[79] = t[116] ? x[50] : x[49];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] & t[118];
  assign t[81] = t[119] & t[120];
  assign t[82] = ~(t[97] ^ t[50]);
  assign t[83] = t[121] ^ t[120];
  assign t[84] = ~(t[87] | t[86]);
  assign t[85] = ~(t[122] | t[54]);
  assign t[86] = ~(t[188]);
  assign t[87] = ~(t[182]);
  assign t[88] = ~(t[16]);
  assign t[89] = ~(t[189]);
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[123] ? t[124] : t[190];
  assign t[91] = ~(t[125]);
  assign t[92] = t[178] ^ t[126];
  assign t[93] = t[127];
  assign t[94] = ~(t[61] ^ t[46]);
  assign t[95] = t[24] ^ t[112];
  assign t[96] = t[69] ^ t[128];
  assign t[97] = t[129] ^ t[130];
  assign t[98] = t[123] ? t[131] : t[191];
  assign t[99] = t[132] ^ t[60];
  assign t[9] = t[173] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind72(x, y);
 input [116:0] x;
 output y;

 wire [360:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[42] ^ t[124];
  assign t[101] = t[125] ? t[126] : t[191];
  assign t[102] = t[125] ? t[127] : t[192];
  assign t[103] = ~(t[70] ^ t[128]);
  assign t[104] = t[129] ^ t[130];
  assign t[105] = t[61] ? t[131] : t[193];
  assign t[106] = ~(t[75] ^ t[132]);
  assign t[107] = t[133] ^ t[134];
  assign t[108] = t[135] ? x[75] : x[74];
  assign t[109] = ~(t[134]);
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[136]);
  assign t[111] = ~(t[72]);
  assign t[112] = t[188] ^ t[137];
  assign t[113] = t[136] ^ t[72];
  assign t[114] = ~(t[173]);
  assign t[115] = t[31] ? x[77] : x[76];
  assign t[116] = t[31] ? x[79] : x[78];
  assign t[117] = t[189] ^ t[138];
  assign t[118] = t[31] ? x[81] : x[80];
  assign t[119] = ~(t[139]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[61] ? t[140] : t[194];
  assign t[121] = t[190] ^ t[141];
  assign t[122] = t[142] ^ t[21];
  assign t[123] = t[143] & t[144];
  assign t[124] = t[145] & t[146];
  assign t[125] = ~(t[88]);
  assign t[126] = t[191] ^ t[147];
  assign t[127] = t[192] ^ t[148];
  assign t[128] = t[149] ^ t[150];
  assign t[129] = t[102] ^ t[151];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[125] ? t[152] : t[195];
  assign t[131] = t[193] ^ t[153];
  assign t[132] = t[46] ^ t[136];
  assign t[133] = t[136] ^ t[26];
  assign t[134] = t[112] ^ t[72];
  assign t[135] = ~(t[139]);
  assign t[136] = t[61] ? t[154] : t[196];
  assign t[137] = t[61] ? t[155] : t[197];
  assign t[138] = t[135] ? x[95] : x[94];
  assign t[139] = ~(t[31]);
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[194] ^ t[156];
  assign t[141] = t[119] ? x[97] : x[96];
  assign t[142] = t[157] & t[158];
  assign t[143] = ~(t[142] ^ t[159]);
  assign t[144] = t[20] ^ t[160];
  assign t[145] = ~(t[161] ^ t[42]);
  assign t[146] = t[22] ^ t[94];
  assign t[147] = t[162] ? x[99] : x[98];
  assign t[148] = t[162] ? x[101] : x[100];
  assign t[149] = t[163] & t[164];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[165] & t[130];
  assign t[151] = t[125] ? t[166] : t[198];
  assign t[152] = t[195] ^ t[167];
  assign t[153] = t[135] ? x[106] : x[105];
  assign t[154] = t[196] ^ t[168];
  assign t[155] = t[197] ^ t[169];
  assign t[156] = t[119] ? x[108] : x[107];
  assign t[157] = ~(t[160]);
  assign t[158] = ~(t[36]);
  assign t[159] = t[98] ^ t[36];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[39] ^ t[59];
  assign t[161] = t[120] ^ t[40];
  assign t[162] = ~(t[139]);
  assign t[163] = ~(t[170]);
  assign t[164] = ~(t[101]);
  assign t[165] = ~(t[102]);
  assign t[166] = t[198] ^ t[171];
  assign t[167] = t[162] ? x[110] : x[109];
  assign t[168] = t[135] ? x[112] : x[111];
  assign t[169] = t[135] ? x[114] : x[113];
  assign t[16] = t[173] | t[30];
  assign t[170] = t[130] ^ t[102];
  assign t[171] = t[162] ? x[116] : x[115];
  assign t[172] = (t[199]);
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = t[226] ^ x[4];
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[7];
  assign t[201] = t[228] ^ x[12];
  assign t[202] = t[229] ^ x[15];
  assign t[203] = t[230] ^ x[18];
  assign t[204] = t[231] ^ x[21];
  assign t[205] = t[232] ^ x[24];
  assign t[206] = t[233] ^ x[27];
  assign t[207] = t[234] ^ x[30];
  assign t[208] = t[235] ^ x[33];
  assign t[209] = t[236] ^ x[36];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[39];
  assign t[211] = t[238] ^ x[42];
  assign t[212] = t[239] ^ x[45];
  assign t[213] = t[240] ^ x[48];
  assign t[214] = t[241] ^ x[51];
  assign t[215] = t[242] ^ x[54];
  assign t[216] = t[243] ^ x[57];
  assign t[217] = t[244] ^ x[64];
  assign t[218] = t[245] ^ x[67];
  assign t[219] = t[246] ^ x[70];
  assign t[21] = t[38] & t[39];
  assign t[220] = t[247] ^ x[73];
  assign t[221] = t[248] ^ x[84];
  assign t[222] = t[249] ^ x[87];
  assign t[223] = t[250] ^ x[90];
  assign t[224] = t[251] ^ x[93];
  assign t[225] = t[252] ^ x[104];
  assign t[226] = (t[253] & ~t[254]);
  assign t[227] = (t[255] & ~t[256]);
  assign t[228] = (t[257] & ~t[258]);
  assign t[229] = (t[259] & ~t[260]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[261] & ~t[262]);
  assign t[231] = (t[263] & ~t[264]);
  assign t[232] = (t[265] & ~t[266]);
  assign t[233] = (t[267] & ~t[268]);
  assign t[234] = (t[269] & ~t[270]);
  assign t[235] = (t[271] & ~t[272]);
  assign t[236] = (t[273] & ~t[274]);
  assign t[237] = (t[275] & ~t[276]);
  assign t[238] = (t[277] & ~t[278]);
  assign t[239] = (t[279] & ~t[280]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (t[281] & ~t[282]);
  assign t[241] = (t[283] & ~t[284]);
  assign t[242] = (t[285] & ~t[286]);
  assign t[243] = (t[287] & ~t[288]);
  assign t[244] = (t[289] & ~t[290]);
  assign t[245] = (t[291] & ~t[292]);
  assign t[246] = (t[293] & ~t[294]);
  assign t[247] = (t[295] & ~t[296]);
  assign t[248] = (t[297] & ~t[298]);
  assign t[249] = (t[299] & ~t[300]);
  assign t[24] = ~(t[44] ^ t[45]);
  assign t[250] = (t[301] & ~t[302]);
  assign t[251] = (t[303] & ~t[304]);
  assign t[252] = (t[305] & ~t[306]);
  assign t[253] = t[307] ^ x[4];
  assign t[254] = t[308] ^ x[3];
  assign t[255] = t[309] ^ x[7];
  assign t[256] = t[310] ^ x[6];
  assign t[257] = t[311] ^ x[12];
  assign t[258] = t[312] ^ x[11];
  assign t[259] = t[313] ^ x[15];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[314] ^ x[14];
  assign t[261] = t[315] ^ x[18];
  assign t[262] = t[316] ^ x[17];
  assign t[263] = t[317] ^ x[21];
  assign t[264] = t[318] ^ x[20];
  assign t[265] = t[319] ^ x[24];
  assign t[266] = t[320] ^ x[23];
  assign t[267] = t[321] ^ x[27];
  assign t[268] = t[322] ^ x[26];
  assign t[269] = t[323] ^ x[30];
  assign t[26] = t[174] ^ t[48];
  assign t[270] = t[324] ^ x[29];
  assign t[271] = t[325] ^ x[33];
  assign t[272] = t[326] ^ x[32];
  assign t[273] = t[327] ^ x[36];
  assign t[274] = t[328] ^ x[35];
  assign t[275] = t[329] ^ x[39];
  assign t[276] = t[330] ^ x[38];
  assign t[277] = t[331] ^ x[42];
  assign t[278] = t[332] ^ x[41];
  assign t[279] = t[333] ^ x[45];
  assign t[27] = t[49] ^ t[50];
  assign t[280] = t[334] ^ x[44];
  assign t[281] = t[335] ^ x[48];
  assign t[282] = t[336] ^ x[47];
  assign t[283] = t[337] ^ x[51];
  assign t[284] = t[338] ^ x[50];
  assign t[285] = t[339] ^ x[54];
  assign t[286] = t[340] ^ x[53];
  assign t[287] = t[341] ^ x[57];
  assign t[288] = t[342] ^ x[56];
  assign t[289] = t[343] ^ x[64];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[63];
  assign t[291] = t[345] ^ x[67];
  assign t[292] = t[346] ^ x[66];
  assign t[293] = t[347] ^ x[70];
  assign t[294] = t[348] ^ x[69];
  assign t[295] = t[349] ^ x[73];
  assign t[296] = t[350] ^ x[72];
  assign t[297] = t[351] ^ x[84];
  assign t[298] = t[352] ^ x[83];
  assign t[299] = t[353] ^ x[87];
  assign t[29] = ~(t[175] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[86];
  assign t[301] = t[355] ^ x[90];
  assign t[302] = t[356] ^ x[89];
  assign t[303] = t[357] ^ x[93];
  assign t[304] = t[358] ^ x[92];
  assign t[305] = t[359] ^ x[104];
  assign t[306] = t[360] ^ x[103];
  assign t[307] = (x[2]);
  assign t[308] = (x[2]);
  assign t[309] = (x[5]);
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = (x[5]);
  assign t[311] = (x[10]);
  assign t[312] = (x[10]);
  assign t[313] = (x[13]);
  assign t[314] = (x[13]);
  assign t[315] = (x[16]);
  assign t[316] = (x[16]);
  assign t[317] = (x[19]);
  assign t[318] = (x[19]);
  assign t[319] = (x[22]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[22]);
  assign t[321] = (x[25]);
  assign t[322] = (x[25]);
  assign t[323] = (x[28]);
  assign t[324] = (x[28]);
  assign t[325] = (x[31]);
  assign t[326] = (x[31]);
  assign t[327] = (x[34]);
  assign t[328] = (x[34]);
  assign t[329] = (x[37]);
  assign t[32] = ~(t[176]);
  assign t[330] = (x[37]);
  assign t[331] = (x[40]);
  assign t[332] = (x[40]);
  assign t[333] = (x[43]);
  assign t[334] = (x[43]);
  assign t[335] = (x[46]);
  assign t[336] = (x[46]);
  assign t[337] = (x[49]);
  assign t[338] = (x[49]);
  assign t[339] = (x[52]);
  assign t[33] = ~(t[177]);
  assign t[340] = (x[52]);
  assign t[341] = (x[55]);
  assign t[342] = (x[55]);
  assign t[343] = (x[62]);
  assign t[344] = (x[62]);
  assign t[345] = (x[65]);
  assign t[346] = (x[65]);
  assign t[347] = (x[68]);
  assign t[348] = (x[68]);
  assign t[349] = (x[71]);
  assign t[34] = ~(t[178]);
  assign t[350] = (x[71]);
  assign t[351] = (x[82]);
  assign t[352] = (x[82]);
  assign t[353] = (x[85]);
  assign t[354] = (x[85]);
  assign t[355] = (x[88]);
  assign t[356] = (x[88]);
  assign t[357] = (x[91]);
  assign t[358] = (x[91]);
  assign t[359] = (x[102]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[102]);
  assign t[36] = t[57];
  assign t[37] = t[58];
  assign t[38] = ~(t[59]);
  assign t[39] = t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[61] ? t[62] : t[179];
  assign t[41] = t[61] ? t[63] : t[180];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] ^ t[26];
  assign t[47] = t[49] ^ t[73];
  assign t[48] = t[61] ? t[74] : t[181];
  assign t[49] = t[75] ^ t[76];
  assign t[4] = t[8] ? t[9] : t[172];
  assign t[50] = t[77] & t[78];
  assign t[51] = ~(t[79] & t[80]);
  assign t[52] = t[81] ^ t[182];
  assign t[53] = ~(t[175]);
  assign t[54] = t[82] & t[81];
  assign t[55] = ~(t[174]);
  assign t[56] = ~(t[83] & t[183]);
  assign t[57] = t[61] ? t[84] : t[184];
  assign t[58] = t[61] ? t[85] : t[185];
  assign t[59] = ~t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[61] ? t[87] : t[186];
  assign t[61] = ~(t[88]);
  assign t[62] = t[179] ^ t[89];
  assign t[63] = t[180] ^ t[90];
  assign t[64] = t[91] & t[92];
  assign t[65] = t[93] & t[94];
  assign t[66] = ~(t[64] ^ t[95]);
  assign t[67] = t[96] ^ t[97];
  assign t[68] = t[98] ^ t[99];
  assign t[69] = t[41] ^ t[100];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[101] ^ t[102];
  assign t[71] = t[103] & t[104];
  assign t[72] = t[178] ^ t[105];
  assign t[73] = t[106] & t[107];
  assign t[74] = t[181] ^ t[108];
  assign t[75] = t[109] & t[110];
  assign t[76] = t[111] & t[112];
  assign t[77] = ~(t[113] ^ t[49]);
  assign t[78] = t[46] ^ t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[114] | t[53]);
  assign t[81] = ~(t[187]);
  assign t[82] = ~(t[182]);
  assign t[83] = ~(t[188]);
  assign t[84] = t[184] ^ t[115];
  assign t[85] = t[185] ^ t[116];
  assign t[86] = t[61] ? t[117] : t[189];
  assign t[87] = t[186] ^ t[118];
  assign t[88] = ~(t[8]);
  assign t[89] = t[119] ? x[59] : x[58];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[31] ? x[61] : x[60];
  assign t[91] = ~(t[97]);
  assign t[92] = ~(t[120]);
  assign t[93] = ~(t[40]);
  assign t[94] = t[61] ? t[121] : t[190];
  assign t[95] = t[22] ^ t[120];
  assign t[96] = t[120] ^ t[41];
  assign t[97] = t[94] ^ t[40];
  assign t[98] = t[59] ^ t[37];
  assign t[99] = t[122] ^ t[123];
  assign t[9] = t[172] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind73(x, y);
 input [116:0] x;
 output y;

 wire [360:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[42] ^ t[124];
  assign t[101] = t[125] ? t[126] : t[191];
  assign t[102] = t[125] ? t[127] : t[192];
  assign t[103] = ~(t[70] ^ t[128]);
  assign t[104] = t[129] ^ t[130];
  assign t[105] = t[61] ? t[131] : t[193];
  assign t[106] = ~(t[75] ^ t[132]);
  assign t[107] = t[133] ^ t[134];
  assign t[108] = t[135] ? x[75] : x[74];
  assign t[109] = ~(t[134]);
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[136]);
  assign t[111] = ~(t[72]);
  assign t[112] = t[188] ^ t[137];
  assign t[113] = t[136] ^ t[72];
  assign t[114] = ~(t[173]);
  assign t[115] = t[31] ? x[77] : x[76];
  assign t[116] = t[31] ? x[79] : x[78];
  assign t[117] = t[189] ^ t[138];
  assign t[118] = t[31] ? x[81] : x[80];
  assign t[119] = ~(t[139]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[61] ? t[140] : t[194];
  assign t[121] = t[190] ^ t[141];
  assign t[122] = t[142] ^ t[21];
  assign t[123] = t[143] & t[144];
  assign t[124] = t[145] & t[146];
  assign t[125] = ~(t[88]);
  assign t[126] = t[191] ^ t[147];
  assign t[127] = t[192] ^ t[148];
  assign t[128] = t[149] ^ t[150];
  assign t[129] = t[102] ^ t[151];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[125] ? t[152] : t[195];
  assign t[131] = t[193] ^ t[153];
  assign t[132] = t[46] ^ t[136];
  assign t[133] = t[136] ^ t[26];
  assign t[134] = t[112] ^ t[72];
  assign t[135] = ~(t[139]);
  assign t[136] = t[61] ? t[154] : t[196];
  assign t[137] = t[61] ? t[155] : t[197];
  assign t[138] = t[135] ? x[95] : x[94];
  assign t[139] = ~(t[31]);
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[194] ^ t[156];
  assign t[141] = t[119] ? x[97] : x[96];
  assign t[142] = t[157] & t[158];
  assign t[143] = ~(t[142] ^ t[159]);
  assign t[144] = t[20] ^ t[160];
  assign t[145] = ~(t[161] ^ t[42]);
  assign t[146] = t[22] ^ t[94];
  assign t[147] = t[162] ? x[99] : x[98];
  assign t[148] = t[162] ? x[101] : x[100];
  assign t[149] = t[163] & t[164];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[165] & t[130];
  assign t[151] = t[125] ? t[166] : t[198];
  assign t[152] = t[195] ^ t[167];
  assign t[153] = t[135] ? x[106] : x[105];
  assign t[154] = t[196] ^ t[168];
  assign t[155] = t[197] ^ t[169];
  assign t[156] = t[119] ? x[108] : x[107];
  assign t[157] = ~(t[160]);
  assign t[158] = ~(t[36]);
  assign t[159] = t[98] ^ t[36];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[39] ^ t[59];
  assign t[161] = t[120] ^ t[40];
  assign t[162] = ~(t[139]);
  assign t[163] = ~(t[170]);
  assign t[164] = ~(t[101]);
  assign t[165] = ~(t[102]);
  assign t[166] = t[198] ^ t[171];
  assign t[167] = t[162] ? x[110] : x[109];
  assign t[168] = t[135] ? x[112] : x[111];
  assign t[169] = t[135] ? x[114] : x[113];
  assign t[16] = t[173] | t[30];
  assign t[170] = t[130] ^ t[102];
  assign t[171] = t[162] ? x[116] : x[115];
  assign t[172] = (t[199]);
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = t[226] ^ x[4];
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[7];
  assign t[201] = t[228] ^ x[12];
  assign t[202] = t[229] ^ x[15];
  assign t[203] = t[230] ^ x[18];
  assign t[204] = t[231] ^ x[21];
  assign t[205] = t[232] ^ x[24];
  assign t[206] = t[233] ^ x[27];
  assign t[207] = t[234] ^ x[30];
  assign t[208] = t[235] ^ x[33];
  assign t[209] = t[236] ^ x[36];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[39];
  assign t[211] = t[238] ^ x[42];
  assign t[212] = t[239] ^ x[45];
  assign t[213] = t[240] ^ x[48];
  assign t[214] = t[241] ^ x[51];
  assign t[215] = t[242] ^ x[54];
  assign t[216] = t[243] ^ x[57];
  assign t[217] = t[244] ^ x[64];
  assign t[218] = t[245] ^ x[67];
  assign t[219] = t[246] ^ x[70];
  assign t[21] = t[38] & t[39];
  assign t[220] = t[247] ^ x[73];
  assign t[221] = t[248] ^ x[84];
  assign t[222] = t[249] ^ x[87];
  assign t[223] = t[250] ^ x[90];
  assign t[224] = t[251] ^ x[93];
  assign t[225] = t[252] ^ x[104];
  assign t[226] = (t[253] & ~t[254]);
  assign t[227] = (t[255] & ~t[256]);
  assign t[228] = (t[257] & ~t[258]);
  assign t[229] = (t[259] & ~t[260]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[261] & ~t[262]);
  assign t[231] = (t[263] & ~t[264]);
  assign t[232] = (t[265] & ~t[266]);
  assign t[233] = (t[267] & ~t[268]);
  assign t[234] = (t[269] & ~t[270]);
  assign t[235] = (t[271] & ~t[272]);
  assign t[236] = (t[273] & ~t[274]);
  assign t[237] = (t[275] & ~t[276]);
  assign t[238] = (t[277] & ~t[278]);
  assign t[239] = (t[279] & ~t[280]);
  assign t[23] = t[42] ^ t[43];
  assign t[240] = (t[281] & ~t[282]);
  assign t[241] = (t[283] & ~t[284]);
  assign t[242] = (t[285] & ~t[286]);
  assign t[243] = (t[287] & ~t[288]);
  assign t[244] = (t[289] & ~t[290]);
  assign t[245] = (t[291] & ~t[292]);
  assign t[246] = (t[293] & ~t[294]);
  assign t[247] = (t[295] & ~t[296]);
  assign t[248] = (t[297] & ~t[298]);
  assign t[249] = (t[299] & ~t[300]);
  assign t[24] = ~(t[44] ^ t[45]);
  assign t[250] = (t[301] & ~t[302]);
  assign t[251] = (t[303] & ~t[304]);
  assign t[252] = (t[305] & ~t[306]);
  assign t[253] = t[307] ^ x[4];
  assign t[254] = t[308] ^ x[3];
  assign t[255] = t[309] ^ x[7];
  assign t[256] = t[310] ^ x[6];
  assign t[257] = t[311] ^ x[12];
  assign t[258] = t[312] ^ x[11];
  assign t[259] = t[313] ^ x[15];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[314] ^ x[14];
  assign t[261] = t[315] ^ x[18];
  assign t[262] = t[316] ^ x[17];
  assign t[263] = t[317] ^ x[21];
  assign t[264] = t[318] ^ x[20];
  assign t[265] = t[319] ^ x[24];
  assign t[266] = t[320] ^ x[23];
  assign t[267] = t[321] ^ x[27];
  assign t[268] = t[322] ^ x[26];
  assign t[269] = t[323] ^ x[30];
  assign t[26] = t[174] ^ t[48];
  assign t[270] = t[324] ^ x[29];
  assign t[271] = t[325] ^ x[33];
  assign t[272] = t[326] ^ x[32];
  assign t[273] = t[327] ^ x[36];
  assign t[274] = t[328] ^ x[35];
  assign t[275] = t[329] ^ x[39];
  assign t[276] = t[330] ^ x[38];
  assign t[277] = t[331] ^ x[42];
  assign t[278] = t[332] ^ x[41];
  assign t[279] = t[333] ^ x[45];
  assign t[27] = t[49] ^ t[50];
  assign t[280] = t[334] ^ x[44];
  assign t[281] = t[335] ^ x[48];
  assign t[282] = t[336] ^ x[47];
  assign t[283] = t[337] ^ x[51];
  assign t[284] = t[338] ^ x[50];
  assign t[285] = t[339] ^ x[54];
  assign t[286] = t[340] ^ x[53];
  assign t[287] = t[341] ^ x[57];
  assign t[288] = t[342] ^ x[56];
  assign t[289] = t[343] ^ x[64];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[63];
  assign t[291] = t[345] ^ x[67];
  assign t[292] = t[346] ^ x[66];
  assign t[293] = t[347] ^ x[70];
  assign t[294] = t[348] ^ x[69];
  assign t[295] = t[349] ^ x[73];
  assign t[296] = t[350] ^ x[72];
  assign t[297] = t[351] ^ x[84];
  assign t[298] = t[352] ^ x[83];
  assign t[299] = t[353] ^ x[87];
  assign t[29] = ~(t[175] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[86];
  assign t[301] = t[355] ^ x[90];
  assign t[302] = t[356] ^ x[89];
  assign t[303] = t[357] ^ x[93];
  assign t[304] = t[358] ^ x[92];
  assign t[305] = t[359] ^ x[104];
  assign t[306] = t[360] ^ x[103];
  assign t[307] = (x[2]);
  assign t[308] = (x[2]);
  assign t[309] = (x[5]);
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = (x[5]);
  assign t[311] = (x[10]);
  assign t[312] = (x[10]);
  assign t[313] = (x[13]);
  assign t[314] = (x[13]);
  assign t[315] = (x[16]);
  assign t[316] = (x[16]);
  assign t[317] = (x[19]);
  assign t[318] = (x[19]);
  assign t[319] = (x[22]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[22]);
  assign t[321] = (x[25]);
  assign t[322] = (x[25]);
  assign t[323] = (x[28]);
  assign t[324] = (x[28]);
  assign t[325] = (x[31]);
  assign t[326] = (x[31]);
  assign t[327] = (x[34]);
  assign t[328] = (x[34]);
  assign t[329] = (x[37]);
  assign t[32] = ~(t[176]);
  assign t[330] = (x[37]);
  assign t[331] = (x[40]);
  assign t[332] = (x[40]);
  assign t[333] = (x[43]);
  assign t[334] = (x[43]);
  assign t[335] = (x[46]);
  assign t[336] = (x[46]);
  assign t[337] = (x[49]);
  assign t[338] = (x[49]);
  assign t[339] = (x[52]);
  assign t[33] = ~(t[177]);
  assign t[340] = (x[52]);
  assign t[341] = (x[55]);
  assign t[342] = (x[55]);
  assign t[343] = (x[62]);
  assign t[344] = (x[62]);
  assign t[345] = (x[65]);
  assign t[346] = (x[65]);
  assign t[347] = (x[68]);
  assign t[348] = (x[68]);
  assign t[349] = (x[71]);
  assign t[34] = ~(t[178]);
  assign t[350] = (x[71]);
  assign t[351] = (x[82]);
  assign t[352] = (x[82]);
  assign t[353] = (x[85]);
  assign t[354] = (x[85]);
  assign t[355] = (x[88]);
  assign t[356] = (x[88]);
  assign t[357] = (x[91]);
  assign t[358] = (x[91]);
  assign t[359] = (x[102]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[102]);
  assign t[36] = t[57];
  assign t[37] = t[58];
  assign t[38] = ~(t[59]);
  assign t[39] = t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[61] ? t[62] : t[179];
  assign t[41] = t[61] ? t[63] : t[180];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] ^ t[26];
  assign t[47] = t[49] ^ t[73];
  assign t[48] = t[61] ? t[74] : t[181];
  assign t[49] = t[75] ^ t[76];
  assign t[4] = t[8] ? t[9] : t[172];
  assign t[50] = t[77] & t[78];
  assign t[51] = ~(t[79] & t[80]);
  assign t[52] = t[81] ^ t[182];
  assign t[53] = ~(t[175]);
  assign t[54] = t[82] & t[81];
  assign t[55] = ~(t[174]);
  assign t[56] = ~(t[83] & t[183]);
  assign t[57] = t[61] ? t[84] : t[184];
  assign t[58] = t[61] ? t[85] : t[185];
  assign t[59] = ~t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = t[61] ? t[87] : t[186];
  assign t[61] = ~(t[88]);
  assign t[62] = t[179] ^ t[89];
  assign t[63] = t[180] ^ t[90];
  assign t[64] = t[91] & t[92];
  assign t[65] = t[93] & t[94];
  assign t[66] = ~(t[64] ^ t[95]);
  assign t[67] = t[96] ^ t[97];
  assign t[68] = t[98] ^ t[99];
  assign t[69] = t[41] ^ t[100];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[101] ^ t[102];
  assign t[71] = t[103] & t[104];
  assign t[72] = t[178] ^ t[105];
  assign t[73] = t[106] & t[107];
  assign t[74] = t[181] ^ t[108];
  assign t[75] = t[109] & t[110];
  assign t[76] = t[111] & t[112];
  assign t[77] = ~(t[113] ^ t[49]);
  assign t[78] = t[46] ^ t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[114] | t[53]);
  assign t[81] = ~(t[187]);
  assign t[82] = ~(t[182]);
  assign t[83] = ~(t[188]);
  assign t[84] = t[184] ^ t[115];
  assign t[85] = t[185] ^ t[116];
  assign t[86] = t[61] ? t[117] : t[189];
  assign t[87] = t[186] ^ t[118];
  assign t[88] = ~(t[8]);
  assign t[89] = t[119] ? x[59] : x[58];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[31] ? x[61] : x[60];
  assign t[91] = ~(t[97]);
  assign t[92] = ~(t[120]);
  assign t[93] = ~(t[40]);
  assign t[94] = t[61] ? t[121] : t[190];
  assign t[95] = t[22] ^ t[120];
  assign t[96] = t[120] ^ t[41];
  assign t[97] = t[94] ^ t[40];
  assign t[98] = t[59] ^ t[37];
  assign t[99] = t[122] ^ t[123];
  assign t[9] = t[172] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind74(x, y);
 input [116:0] x;
 output y;

 wire [381:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[125];
  assign t[101] = ~t[126];
  assign t[102] = ~(t[70] ^ t[127]);
  assign t[103] = t[128] ^ t[129];
  assign t[104] = t[128] ^ t[130];
  assign t[105] = t[131] ^ t[132];
  assign t[106] = t[133] & t[134];
  assign t[107] = t[135] & t[136];
  assign t[108] = t[132] ^ t[137];
  assign t[109] = t[138] ^ t[139];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[140] ^ t[42];
  assign t[111] = t[141];
  assign t[112] = t[127] ^ t[71];
  assign t[113] = ~(t[194]);
  assign t[114] = t[41] ^ t[63];
  assign t[115] = t[208] ^ t[142];
  assign t[116] = t[31] ? x[62] : x[61];
  assign t[117] = ~(t[143]);
  assign t[118] = ~(t[140]);
  assign t[119] = ~(t[98]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[57] ? t[144] : t[210];
  assign t[121] = t[140] ^ t[98];
  assign t[122] = t[209] ^ t[145];
  assign t[123] = ~(t[94] ^ t[146]);
  assign t[124] = t[110] ^ t[143];
  assign t[125] = t[57] ? t[147] : t[211];
  assign t[126] = t[57] ? t[148] : t[212];
  assign t[127] = t[149] ^ t[150];
  assign t[128] = t[101] ^ t[111];
  assign t[129] = t[151];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[127] ^ t[152];
  assign t[131] = t[153] ? t[154] : t[213];
  assign t[132] = t[153] ? t[155] : t[214];
  assign t[133] = ~(t[105] ^ t[138]);
  assign t[134] = t[108] ^ t[156];
  assign t[135] = ~(t[59] ^ t[157]);
  assign t[136] = t[22] ^ t[114];
  assign t[137] = t[153] ? t[158] : t[215];
  assign t[138] = t[159] ^ t[160];
  assign t[139] = t[161] & t[162];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[57] ? t[163] : t[216];
  assign t[141] = t[57] ? t[164] : t[217];
  assign t[142] = t[31] ? x[88] : x[87];
  assign t[143] = t[120] ^ t[98];
  assign t[144] = t[210] ^ t[165];
  assign t[145] = t[166] ? x[90] : x[89];
  assign t[146] = t[68] ^ t[140];
  assign t[147] = t[211] ^ t[167];
  assign t[148] = t[212] ^ t[168];
  assign t[149] = t[169] & t[170];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[171] & t[129];
  assign t[151] = t[57] ? t[172] : t[218];
  assign t[152] = t[173] & t[174];
  assign t[153] = ~(t[85]);
  assign t[154] = t[213] ^ t[175];
  assign t[155] = t[214] ^ t[176];
  assign t[156] = t[153] ? t[177] : t[219];
  assign t[157] = t[74] ^ t[39];
  assign t[158] = t[215] ^ t[178];
  assign t[159] = t[179] & t[180];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[181] & t[156];
  assign t[161] = ~(t[159] ^ t[182]);
  assign t[162] = t[183] ^ t[184];
  assign t[163] = t[216] ^ t[185];
  assign t[164] = t[217] ^ t[186];
  assign t[165] = t[166] ? x[98] : x[97];
  assign t[166] = ~(t[54]);
  assign t[167] = t[83] ? x[100] : x[99];
  assign t[168] = t[31] ? x[102] : x[101];
  assign t[169] = ~(t[187]);
  assign t[16] = t[194] | t[30];
  assign t[170] = ~(t[100]);
  assign t[171] = ~(t[101]);
  assign t[172] = t[218] ^ t[188];
  assign t[173] = ~(t[149] ^ t[189]);
  assign t[174] = t[190] ^ t[187];
  assign t[175] = t[191] ? x[104] : x[103];
  assign t[176] = t[191] ? x[106] : x[105];
  assign t[177] = t[219] ^ t[192];
  assign t[178] = t[191] ? x[108] : x[107];
  assign t[179] = ~(t[184]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = ~(t[131]);
  assign t[181] = ~(t[132]);
  assign t[182] = t[108] ^ t[131];
  assign t[183] = t[131] ^ t[137];
  assign t[184] = t[156] ^ t[132];
  assign t[185] = t[166] ? x[110] : x[109];
  assign t[186] = t[83] ? x[112] : x[111];
  assign t[187] = t[129] ^ t[101];
  assign t[188] = t[83] ? x[114] : x[113];
  assign t[189] = t[128] ^ t[100];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[100] ^ t[111];
  assign t[191] = ~(t[54]);
  assign t[192] = t[191] ? x[116] : x[115];
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[195] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[4];
  assign t[221] = t[248] ^ x[7];
  assign t[222] = t[249] ^ x[12];
  assign t[223] = t[250] ^ x[15];
  assign t[224] = t[251] ^ x[18];
  assign t[225] = t[252] ^ x[21];
  assign t[226] = t[253] ^ x[24];
  assign t[227] = t[254] ^ x[27];
  assign t[228] = t[255] ^ x[30];
  assign t[229] = t[256] ^ x[33];
  assign t[22] = t[39] ^ t[20];
  assign t[230] = t[257] ^ x[36];
  assign t[231] = t[258] ^ x[39];
  assign t[232] = t[259] ^ x[42];
  assign t[233] = t[260] ^ x[45];
  assign t[234] = t[261] ^ x[48];
  assign t[235] = t[262] ^ x[55];
  assign t[236] = t[263] ^ x[60];
  assign t[237] = t[264] ^ x[65];
  assign t[238] = t[265] ^ x[68];
  assign t[239] = t[266] ^ x[71];
  assign t[23] = t[40] & t[41];
  assign t[240] = t[267] ^ x[74];
  assign t[241] = t[268] ^ x[77];
  assign t[242] = t[269] ^ x[80];
  assign t[243] = t[270] ^ x[83];
  assign t[244] = t[271] ^ x[86];
  assign t[245] = t[272] ^ x[93];
  assign t[246] = t[273] ^ x[96];
  assign t[247] = (t[274] & ~t[275]);
  assign t[248] = (t[276] & ~t[277]);
  assign t[249] = (t[278] & ~t[279]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[280] & ~t[281]);
  assign t[251] = (t[282] & ~t[283]);
  assign t[252] = (t[284] & ~t[285]);
  assign t[253] = (t[286] & ~t[287]);
  assign t[254] = (t[288] & ~t[289]);
  assign t[255] = (t[290] & ~t[291]);
  assign t[256] = (t[292] & ~t[293]);
  assign t[257] = (t[294] & ~t[295]);
  assign t[258] = (t[296] & ~t[297]);
  assign t[259] = (t[298] & ~t[299]);
  assign t[25] = t[44] ^ t[45];
  assign t[260] = (t[300] & ~t[301]);
  assign t[261] = (t[302] & ~t[303]);
  assign t[262] = (t[304] & ~t[305]);
  assign t[263] = (t[306] & ~t[307]);
  assign t[264] = (t[308] & ~t[309]);
  assign t[265] = (t[310] & ~t[311]);
  assign t[266] = (t[312] & ~t[313]);
  assign t[267] = (t[314] & ~t[315]);
  assign t[268] = (t[316] & ~t[317]);
  assign t[269] = (t[318] & ~t[319]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[320] & ~t[321]);
  assign t[271] = (t[322] & ~t[323]);
  assign t[272] = (t[324] & ~t[325]);
  assign t[273] = (t[326] & ~t[327]);
  assign t[274] = t[328] ^ x[4];
  assign t[275] = t[329] ^ x[3];
  assign t[276] = t[330] ^ x[7];
  assign t[277] = t[331] ^ x[6];
  assign t[278] = t[332] ^ x[12];
  assign t[279] = t[333] ^ x[11];
  assign t[27] = ~(t[48] ^ t[49]);
  assign t[280] = t[334] ^ x[15];
  assign t[281] = t[335] ^ x[14];
  assign t[282] = t[336] ^ x[18];
  assign t[283] = t[337] ^ x[17];
  assign t[284] = t[338] ^ x[21];
  assign t[285] = t[339] ^ x[20];
  assign t[286] = t[340] ^ x[24];
  assign t[287] = t[341] ^ x[23];
  assign t[288] = t[342] ^ x[27];
  assign t[289] = t[343] ^ x[26];
  assign t[28] = ~(t[30] & t[50]);
  assign t[290] = t[344] ^ x[30];
  assign t[291] = t[345] ^ x[29];
  assign t[292] = t[346] ^ x[33];
  assign t[293] = t[347] ^ x[32];
  assign t[294] = t[348] ^ x[36];
  assign t[295] = t[349] ^ x[35];
  assign t[296] = t[350] ^ x[39];
  assign t[297] = t[351] ^ x[38];
  assign t[298] = t[352] ^ x[42];
  assign t[299] = t[353] ^ x[41];
  assign t[29] = ~(t[196] ^ t[51]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[45];
  assign t[301] = t[355] ^ x[44];
  assign t[302] = t[356] ^ x[48];
  assign t[303] = t[357] ^ x[47];
  assign t[304] = t[358] ^ x[55];
  assign t[305] = t[359] ^ x[54];
  assign t[306] = t[360] ^ x[60];
  assign t[307] = t[361] ^ x[59];
  assign t[308] = t[362] ^ x[65];
  assign t[309] = t[363] ^ x[64];
  assign t[30] = ~(t[52] & t[53]);
  assign t[310] = t[364] ^ x[68];
  assign t[311] = t[365] ^ x[67];
  assign t[312] = t[366] ^ x[71];
  assign t[313] = t[367] ^ x[70];
  assign t[314] = t[368] ^ x[74];
  assign t[315] = t[369] ^ x[73];
  assign t[316] = t[370] ^ x[77];
  assign t[317] = t[371] ^ x[76];
  assign t[318] = t[372] ^ x[80];
  assign t[319] = t[373] ^ x[79];
  assign t[31] = ~(t[54]);
  assign t[320] = t[374] ^ x[83];
  assign t[321] = t[375] ^ x[82];
  assign t[322] = t[376] ^ x[86];
  assign t[323] = t[377] ^ x[85];
  assign t[324] = t[378] ^ x[93];
  assign t[325] = t[379] ^ x[92];
  assign t[326] = t[380] ^ x[96];
  assign t[327] = t[381] ^ x[95];
  assign t[328] = (x[2]);
  assign t[329] = (x[2]);
  assign t[32] = ~(t[197]);
  assign t[330] = (x[5]);
  assign t[331] = (x[5]);
  assign t[332] = (x[10]);
  assign t[333] = (x[10]);
  assign t[334] = (x[13]);
  assign t[335] = (x[13]);
  assign t[336] = (x[16]);
  assign t[337] = (x[16]);
  assign t[338] = (x[19]);
  assign t[339] = (x[19]);
  assign t[33] = ~(t[198]);
  assign t[340] = (x[22]);
  assign t[341] = (x[22]);
  assign t[342] = (x[25]);
  assign t[343] = (x[25]);
  assign t[344] = (x[28]);
  assign t[345] = (x[28]);
  assign t[346] = (x[31]);
  assign t[347] = (x[31]);
  assign t[348] = (x[34]);
  assign t[349] = (x[34]);
  assign t[34] = ~(t[199]);
  assign t[350] = (x[37]);
  assign t[351] = (x[37]);
  assign t[352] = (x[40]);
  assign t[353] = (x[40]);
  assign t[354] = (x[43]);
  assign t[355] = (x[43]);
  assign t[356] = (x[46]);
  assign t[357] = (x[46]);
  assign t[358] = (x[53]);
  assign t[359] = (x[53]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[58]);
  assign t[361] = (x[58]);
  assign t[362] = (x[63]);
  assign t[363] = (x[63]);
  assign t[364] = (x[66]);
  assign t[365] = (x[66]);
  assign t[366] = (x[69]);
  assign t[367] = (x[69]);
  assign t[368] = (x[72]);
  assign t[369] = (x[72]);
  assign t[36] = t[57] ? t[58] : t[200];
  assign t[370] = (x[75]);
  assign t[371] = (x[75]);
  assign t[372] = (x[78]);
  assign t[373] = (x[78]);
  assign t[374] = (x[81]);
  assign t[375] = (x[81]);
  assign t[376] = (x[84]);
  assign t[377] = (x[84]);
  assign t[378] = (x[91]);
  assign t[379] = (x[91]);
  assign t[37] = t[59] ^ t[23];
  assign t[380] = (x[94]);
  assign t[381] = (x[94]);
  assign t[38] = t[60] & t[61];
  assign t[39] = t[57] ? t[62] : t[201];
  assign t[3] = t[6] ^ t[7];
  assign t[40] = ~(t[63]);
  assign t[41] = t[202] ^ t[64];
  assign t[42] = t[57] ? t[65] : t[203];
  assign t[43] = t[66] ^ t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] ^ t[73]);
  assign t[47] = t[74] ^ t[75];
  assign t[48] = t[76] ^ t[77];
  assign t[49] = ~(t[11] ^ t[78]);
  assign t[4] = t[8] ? t[9] : t[193];
  assign t[50] = ~(t[79] & t[80]);
  assign t[51] = t[81] ^ t[204];
  assign t[52] = ~(t[196]);
  assign t[53] = t[82] & t[81];
  assign t[54] = ~(t[83]);
  assign t[55] = ~(t[195]);
  assign t[56] = ~(t[84] & t[205]);
  assign t[57] = ~(t[85]);
  assign t[58] = t[200] ^ t[86];
  assign t[59] = t[87] & t[88];
  assign t[5] = ~(t[10]);
  assign t[60] = ~(t[89] ^ t[37]);
  assign t[61] = t[74] ^ t[41];
  assign t[62] = t[201] ^ t[90];
  assign t[63] = t[199] ^ t[91];
  assign t[64] = t[57] ? t[92] : t[206];
  assign t[65] = t[203] ^ t[93];
  assign t[66] = t[94] ^ t[95];
  assign t[67] = t[96] & t[97];
  assign t[68] = t[98] ^ t[42];
  assign t[69] = t[66] ^ t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[100] ^ t[101];
  assign t[71] = t[102] & t[103];
  assign t[72] = t[104] ^ t[24];
  assign t[73] = t[105] ^ t[106];
  assign t[74] = t[63] ^ t[20];
  assign t[75] = t[37] ^ t[107];
  assign t[76] = t[108] ^ t[109];
  assign t[77] = t[110] ^ t[95];
  assign t[78] = t[111] ^ t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[113] | t[52]);
  assign t[81] = ~(t[207]);
  assign t[82] = ~(t[204]);
  assign t[83] = ~(t[16]);
  assign t[84] = ~(t[202]);
  assign t[85] = ~(t[8]);
  assign t[86] = t[31] ? x[50] : x[49];
  assign t[87] = ~(t[114]);
  assign t[88] = ~(t[39]);
  assign t[89] = t[39] ^ t[63];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[31] ? x[52] : x[51];
  assign t[91] = t[57] ? t[115] : t[208];
  assign t[92] = t[206] ^ t[116];
  assign t[93] = t[83] ? x[57] : x[56];
  assign t[94] = t[117] & t[118];
  assign t[95] = t[119] & t[120];
  assign t[96] = ~(t[121] ^ t[66]);
  assign t[97] = t[68] ^ t[120];
  assign t[98] = t[57] ? t[122] : t[209];
  assign t[99] = t[123] & t[124];
  assign t[9] = t[193] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [116:0] x;
 output y;

 wire [381:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[125];
  assign t[101] = ~t[126];
  assign t[102] = ~(t[70] ^ t[127]);
  assign t[103] = t[128] ^ t[129];
  assign t[104] = t[128] ^ t[130];
  assign t[105] = t[131] ^ t[132];
  assign t[106] = t[133] & t[134];
  assign t[107] = t[135] & t[136];
  assign t[108] = t[132] ^ t[137];
  assign t[109] = t[138] ^ t[139];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[140] ^ t[42];
  assign t[111] = t[141];
  assign t[112] = t[127] ^ t[71];
  assign t[113] = ~(t[194]);
  assign t[114] = t[41] ^ t[63];
  assign t[115] = t[208] ^ t[142];
  assign t[116] = t[31] ? x[62] : x[61];
  assign t[117] = ~(t[143]);
  assign t[118] = ~(t[140]);
  assign t[119] = ~(t[98]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[57] ? t[144] : t[210];
  assign t[121] = t[140] ^ t[98];
  assign t[122] = t[209] ^ t[145];
  assign t[123] = ~(t[94] ^ t[146]);
  assign t[124] = t[110] ^ t[143];
  assign t[125] = t[57] ? t[147] : t[211];
  assign t[126] = t[57] ? t[148] : t[212];
  assign t[127] = t[149] ^ t[150];
  assign t[128] = t[101] ^ t[111];
  assign t[129] = t[151];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[127] ^ t[152];
  assign t[131] = t[153] ? t[154] : t[213];
  assign t[132] = t[153] ? t[155] : t[214];
  assign t[133] = ~(t[105] ^ t[138]);
  assign t[134] = t[108] ^ t[156];
  assign t[135] = ~(t[59] ^ t[157]);
  assign t[136] = t[22] ^ t[114];
  assign t[137] = t[153] ? t[158] : t[215];
  assign t[138] = t[159] ^ t[160];
  assign t[139] = t[161] & t[162];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[57] ? t[163] : t[216];
  assign t[141] = t[57] ? t[164] : t[217];
  assign t[142] = t[31] ? x[88] : x[87];
  assign t[143] = t[120] ^ t[98];
  assign t[144] = t[210] ^ t[165];
  assign t[145] = t[166] ? x[90] : x[89];
  assign t[146] = t[68] ^ t[140];
  assign t[147] = t[211] ^ t[167];
  assign t[148] = t[212] ^ t[168];
  assign t[149] = t[169] & t[170];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[171] & t[129];
  assign t[151] = t[57] ? t[172] : t[218];
  assign t[152] = t[173] & t[174];
  assign t[153] = ~(t[85]);
  assign t[154] = t[213] ^ t[175];
  assign t[155] = t[214] ^ t[176];
  assign t[156] = t[153] ? t[177] : t[219];
  assign t[157] = t[74] ^ t[39];
  assign t[158] = t[215] ^ t[178];
  assign t[159] = t[179] & t[180];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[181] & t[156];
  assign t[161] = ~(t[159] ^ t[182]);
  assign t[162] = t[183] ^ t[184];
  assign t[163] = t[216] ^ t[185];
  assign t[164] = t[217] ^ t[186];
  assign t[165] = t[166] ? x[98] : x[97];
  assign t[166] = ~(t[54]);
  assign t[167] = t[83] ? x[100] : x[99];
  assign t[168] = t[31] ? x[102] : x[101];
  assign t[169] = ~(t[187]);
  assign t[16] = t[194] | t[30];
  assign t[170] = ~(t[100]);
  assign t[171] = ~(t[101]);
  assign t[172] = t[218] ^ t[188];
  assign t[173] = ~(t[149] ^ t[189]);
  assign t[174] = t[190] ^ t[187];
  assign t[175] = t[191] ? x[104] : x[103];
  assign t[176] = t[191] ? x[106] : x[105];
  assign t[177] = t[219] ^ t[192];
  assign t[178] = t[191] ? x[108] : x[107];
  assign t[179] = ~(t[184]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = ~(t[131]);
  assign t[181] = ~(t[132]);
  assign t[182] = t[108] ^ t[131];
  assign t[183] = t[131] ^ t[137];
  assign t[184] = t[156] ^ t[132];
  assign t[185] = t[166] ? x[110] : x[109];
  assign t[186] = t[83] ? x[112] : x[111];
  assign t[187] = t[129] ^ t[101];
  assign t[188] = t[83] ? x[114] : x[113];
  assign t[189] = t[128] ^ t[100];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = t[100] ^ t[111];
  assign t[191] = ~(t[54]);
  assign t[192] = t[191] ? x[116] : x[115];
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[195] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[4];
  assign t[221] = t[248] ^ x[7];
  assign t[222] = t[249] ^ x[12];
  assign t[223] = t[250] ^ x[15];
  assign t[224] = t[251] ^ x[18];
  assign t[225] = t[252] ^ x[21];
  assign t[226] = t[253] ^ x[24];
  assign t[227] = t[254] ^ x[27];
  assign t[228] = t[255] ^ x[30];
  assign t[229] = t[256] ^ x[33];
  assign t[22] = t[39] ^ t[20];
  assign t[230] = t[257] ^ x[36];
  assign t[231] = t[258] ^ x[39];
  assign t[232] = t[259] ^ x[42];
  assign t[233] = t[260] ^ x[45];
  assign t[234] = t[261] ^ x[48];
  assign t[235] = t[262] ^ x[55];
  assign t[236] = t[263] ^ x[60];
  assign t[237] = t[264] ^ x[65];
  assign t[238] = t[265] ^ x[68];
  assign t[239] = t[266] ^ x[71];
  assign t[23] = t[40] & t[41];
  assign t[240] = t[267] ^ x[74];
  assign t[241] = t[268] ^ x[77];
  assign t[242] = t[269] ^ x[80];
  assign t[243] = t[270] ^ x[83];
  assign t[244] = t[271] ^ x[86];
  assign t[245] = t[272] ^ x[93];
  assign t[246] = t[273] ^ x[96];
  assign t[247] = (t[274] & ~t[275]);
  assign t[248] = (t[276] & ~t[277]);
  assign t[249] = (t[278] & ~t[279]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[280] & ~t[281]);
  assign t[251] = (t[282] & ~t[283]);
  assign t[252] = (t[284] & ~t[285]);
  assign t[253] = (t[286] & ~t[287]);
  assign t[254] = (t[288] & ~t[289]);
  assign t[255] = (t[290] & ~t[291]);
  assign t[256] = (t[292] & ~t[293]);
  assign t[257] = (t[294] & ~t[295]);
  assign t[258] = (t[296] & ~t[297]);
  assign t[259] = (t[298] & ~t[299]);
  assign t[25] = t[44] ^ t[45];
  assign t[260] = (t[300] & ~t[301]);
  assign t[261] = (t[302] & ~t[303]);
  assign t[262] = (t[304] & ~t[305]);
  assign t[263] = (t[306] & ~t[307]);
  assign t[264] = (t[308] & ~t[309]);
  assign t[265] = (t[310] & ~t[311]);
  assign t[266] = (t[312] & ~t[313]);
  assign t[267] = (t[314] & ~t[315]);
  assign t[268] = (t[316] & ~t[317]);
  assign t[269] = (t[318] & ~t[319]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[320] & ~t[321]);
  assign t[271] = (t[322] & ~t[323]);
  assign t[272] = (t[324] & ~t[325]);
  assign t[273] = (t[326] & ~t[327]);
  assign t[274] = t[328] ^ x[4];
  assign t[275] = t[329] ^ x[3];
  assign t[276] = t[330] ^ x[7];
  assign t[277] = t[331] ^ x[6];
  assign t[278] = t[332] ^ x[12];
  assign t[279] = t[333] ^ x[11];
  assign t[27] = ~(t[48] ^ t[49]);
  assign t[280] = t[334] ^ x[15];
  assign t[281] = t[335] ^ x[14];
  assign t[282] = t[336] ^ x[18];
  assign t[283] = t[337] ^ x[17];
  assign t[284] = t[338] ^ x[21];
  assign t[285] = t[339] ^ x[20];
  assign t[286] = t[340] ^ x[24];
  assign t[287] = t[341] ^ x[23];
  assign t[288] = t[342] ^ x[27];
  assign t[289] = t[343] ^ x[26];
  assign t[28] = ~(t[30] & t[50]);
  assign t[290] = t[344] ^ x[30];
  assign t[291] = t[345] ^ x[29];
  assign t[292] = t[346] ^ x[33];
  assign t[293] = t[347] ^ x[32];
  assign t[294] = t[348] ^ x[36];
  assign t[295] = t[349] ^ x[35];
  assign t[296] = t[350] ^ x[39];
  assign t[297] = t[351] ^ x[38];
  assign t[298] = t[352] ^ x[42];
  assign t[299] = t[353] ^ x[41];
  assign t[29] = ~(t[196] ^ t[51]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[45];
  assign t[301] = t[355] ^ x[44];
  assign t[302] = t[356] ^ x[48];
  assign t[303] = t[357] ^ x[47];
  assign t[304] = t[358] ^ x[55];
  assign t[305] = t[359] ^ x[54];
  assign t[306] = t[360] ^ x[60];
  assign t[307] = t[361] ^ x[59];
  assign t[308] = t[362] ^ x[65];
  assign t[309] = t[363] ^ x[64];
  assign t[30] = ~(t[52] & t[53]);
  assign t[310] = t[364] ^ x[68];
  assign t[311] = t[365] ^ x[67];
  assign t[312] = t[366] ^ x[71];
  assign t[313] = t[367] ^ x[70];
  assign t[314] = t[368] ^ x[74];
  assign t[315] = t[369] ^ x[73];
  assign t[316] = t[370] ^ x[77];
  assign t[317] = t[371] ^ x[76];
  assign t[318] = t[372] ^ x[80];
  assign t[319] = t[373] ^ x[79];
  assign t[31] = ~(t[54]);
  assign t[320] = t[374] ^ x[83];
  assign t[321] = t[375] ^ x[82];
  assign t[322] = t[376] ^ x[86];
  assign t[323] = t[377] ^ x[85];
  assign t[324] = t[378] ^ x[93];
  assign t[325] = t[379] ^ x[92];
  assign t[326] = t[380] ^ x[96];
  assign t[327] = t[381] ^ x[95];
  assign t[328] = (x[2]);
  assign t[329] = (x[2]);
  assign t[32] = ~(t[197]);
  assign t[330] = (x[5]);
  assign t[331] = (x[5]);
  assign t[332] = (x[10]);
  assign t[333] = (x[10]);
  assign t[334] = (x[13]);
  assign t[335] = (x[13]);
  assign t[336] = (x[16]);
  assign t[337] = (x[16]);
  assign t[338] = (x[19]);
  assign t[339] = (x[19]);
  assign t[33] = ~(t[198]);
  assign t[340] = (x[22]);
  assign t[341] = (x[22]);
  assign t[342] = (x[25]);
  assign t[343] = (x[25]);
  assign t[344] = (x[28]);
  assign t[345] = (x[28]);
  assign t[346] = (x[31]);
  assign t[347] = (x[31]);
  assign t[348] = (x[34]);
  assign t[349] = (x[34]);
  assign t[34] = ~(t[199]);
  assign t[350] = (x[37]);
  assign t[351] = (x[37]);
  assign t[352] = (x[40]);
  assign t[353] = (x[40]);
  assign t[354] = (x[43]);
  assign t[355] = (x[43]);
  assign t[356] = (x[46]);
  assign t[357] = (x[46]);
  assign t[358] = (x[53]);
  assign t[359] = (x[53]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[58]);
  assign t[361] = (x[58]);
  assign t[362] = (x[63]);
  assign t[363] = (x[63]);
  assign t[364] = (x[66]);
  assign t[365] = (x[66]);
  assign t[366] = (x[69]);
  assign t[367] = (x[69]);
  assign t[368] = (x[72]);
  assign t[369] = (x[72]);
  assign t[36] = t[57] ? t[58] : t[200];
  assign t[370] = (x[75]);
  assign t[371] = (x[75]);
  assign t[372] = (x[78]);
  assign t[373] = (x[78]);
  assign t[374] = (x[81]);
  assign t[375] = (x[81]);
  assign t[376] = (x[84]);
  assign t[377] = (x[84]);
  assign t[378] = (x[91]);
  assign t[379] = (x[91]);
  assign t[37] = t[59] ^ t[23];
  assign t[380] = (x[94]);
  assign t[381] = (x[94]);
  assign t[38] = t[60] & t[61];
  assign t[39] = t[57] ? t[62] : t[201];
  assign t[3] = t[6] ^ t[7];
  assign t[40] = ~(t[63]);
  assign t[41] = t[202] ^ t[64];
  assign t[42] = t[57] ? t[65] : t[203];
  assign t[43] = t[66] ^ t[67];
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[72] ^ t[73]);
  assign t[47] = t[74] ^ t[75];
  assign t[48] = t[76] ^ t[77];
  assign t[49] = ~(t[11] ^ t[78]);
  assign t[4] = t[8] ? t[9] : t[193];
  assign t[50] = ~(t[79] & t[80]);
  assign t[51] = t[81] ^ t[204];
  assign t[52] = ~(t[196]);
  assign t[53] = t[82] & t[81];
  assign t[54] = ~(t[83]);
  assign t[55] = ~(t[195]);
  assign t[56] = ~(t[84] & t[205]);
  assign t[57] = ~(t[85]);
  assign t[58] = t[200] ^ t[86];
  assign t[59] = t[87] & t[88];
  assign t[5] = ~(t[10]);
  assign t[60] = ~(t[89] ^ t[37]);
  assign t[61] = t[74] ^ t[41];
  assign t[62] = t[201] ^ t[90];
  assign t[63] = t[199] ^ t[91];
  assign t[64] = t[57] ? t[92] : t[206];
  assign t[65] = t[203] ^ t[93];
  assign t[66] = t[94] ^ t[95];
  assign t[67] = t[96] & t[97];
  assign t[68] = t[98] ^ t[42];
  assign t[69] = t[66] ^ t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[100] ^ t[101];
  assign t[71] = t[102] & t[103];
  assign t[72] = t[104] ^ t[24];
  assign t[73] = t[105] ^ t[106];
  assign t[74] = t[63] ^ t[20];
  assign t[75] = t[37] ^ t[107];
  assign t[76] = t[108] ^ t[109];
  assign t[77] = t[110] ^ t[95];
  assign t[78] = t[111] ^ t[112];
  assign t[79] = ~(t[82] | t[81]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[113] | t[52]);
  assign t[81] = ~(t[207]);
  assign t[82] = ~(t[204]);
  assign t[83] = ~(t[16]);
  assign t[84] = ~(t[202]);
  assign t[85] = ~(t[8]);
  assign t[86] = t[31] ? x[50] : x[49];
  assign t[87] = ~(t[114]);
  assign t[88] = ~(t[39]);
  assign t[89] = t[39] ^ t[63];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[31] ? x[52] : x[51];
  assign t[91] = t[57] ? t[115] : t[208];
  assign t[92] = t[206] ^ t[116];
  assign t[93] = t[83] ? x[57] : x[56];
  assign t[94] = t[117] & t[118];
  assign t[95] = t[119] & t[120];
  assign t[96] = ~(t[121] ^ t[66]);
  assign t[97] = t[68] ^ t[120];
  assign t[98] = t[57] ? t[122] : t[209];
  assign t[99] = t[123] & t[124];
  assign t[9] = t[193] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind76(x, y);
 input [116:0] x;
 output y;

 wire [370:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[31] ? x[61] : x[60];
  assign t[101] = t[195] ^ t[129];
  assign t[102] = t[128] ? x[63] : x[62];
  assign t[103] = t[65] ? t[130] : t[200];
  assign t[104] = t[131] & t[132];
  assign t[105] = ~(t[104] ^ t[133]);
  assign t[106] = t[61] ^ t[134];
  assign t[107] = t[135] & t[136];
  assign t[108] = ~(t[117] ^ t[73]);
  assign t[109] = t[137] ^ t[43];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[138] ? x[68] : x[67];
  assign t[111] = t[196] ^ t[139];
  assign t[112] = t[140] & t[141];
  assign t[113] = t[65] ? t[142] : t[201];
  assign t[114] = ~(t[183]);
  assign t[115] = t[65] ? t[143] : t[202];
  assign t[116] = ~(t[48]);
  assign t[117] = t[40] ^ t[68];
  assign t[118] = t[144] ? t[145] : t[203];
  assign t[119] = t[121] ^ t[146];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[144] ? t[147] : t[204];
  assign t[121] = t[148] ^ t[149];
  assign t[122] = t[150] & t[151];
  assign t[123] = t[65] ? t[152] : t[205];
  assign t[124] = t[65] ? t[153] : t[206];
  assign t[125] = t[199] ^ t[154];
  assign t[126] = ~(t[155] ^ t[71]);
  assign t[127] = t[44] ^ t[95];
  assign t[128] = ~(t[156]);
  assign t[129] = t[128] ? x[88] : x[87];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[200] ^ t[157];
  assign t[131] = ~(t[134]);
  assign t[132] = ~(t[93]);
  assign t[133] = t[44] ^ t[93];
  assign t[134] = t[95] ^ t[70];
  assign t[135] = ~(t[158]);
  assign t[136] = ~(t[40]);
  assign t[137] = t[68] ^ t[41];
  assign t[138] = ~(t[156]);
  assign t[139] = t[138] ? x[90] : x[89];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[159]);
  assign t[141] = ~(t[47]);
  assign t[142] = t[201] ^ t[160];
  assign t[143] = t[202] ^ t[161];
  assign t[144] = ~(t[98]);
  assign t[145] = t[203] ^ t[162];
  assign t[146] = t[163] & t[164];
  assign t[147] = t[204] ^ t[165];
  assign t[148] = t[166] & t[167];
  assign t[149] = t[168] & t[169];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = ~(t[148] ^ t[170]);
  assign t[151] = t[171] ^ t[172];
  assign t[152] = t[205] ^ t[173];
  assign t[153] = t[206] ^ t[174];
  assign t[154] = t[31] ? x[92] : x[91];
  assign t[155] = t[93] ^ t[70];
  assign t[156] = ~(t[31]);
  assign t[157] = t[138] ? x[94] : x[93];
  assign t[158] = t[43] ^ t[68];
  assign t[159] = t[79] ^ t[48];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[138] ? x[96] : x[95];
  assign t[161] = t[138] ? x[98] : x[97];
  assign t[162] = t[175] ? x[100] : x[99];
  assign t[163] = ~(t[176] ^ t[121]);
  assign t[164] = t[91] ^ t[169];
  assign t[165] = t[175] ? x[102] : x[101];
  assign t[166] = ~(t[172]);
  assign t[167] = ~(t[177]);
  assign t[168] = ~(t[120]);
  assign t[169] = t[144] ? t[178] : t[207];
  assign t[16] = t[183] | t[30];
  assign t[170] = t[91] ^ t[177];
  assign t[171] = t[177] ^ t[118];
  assign t[172] = t[169] ^ t[120];
  assign t[173] = t[31] ? x[107] : x[106];
  assign t[174] = t[31] ? x[109] : x[108];
  assign t[175] = ~(t[156]);
  assign t[176] = t[177] ^ t[120];
  assign t[177] = t[144] ? t[179] : t[208];
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[208] ^ t[181];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[175] ? x[114] : x[113];
  assign t[181] = t[175] ? x[116] : x[115];
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = t[236] ^ x[4];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[7];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[66];
  assign t[228] = t[255] ^ x[71];
  assign t[229] = t[256] ^ x[74];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[77];
  assign t[231] = t[258] ^ x[80];
  assign t[232] = t[259] ^ x[83];
  assign t[233] = t[260] ^ x[86];
  assign t[234] = t[261] ^ x[105];
  assign t[235] = t[262] ^ x[112];
  assign t[236] = (t[263] & ~t[264]);
  assign t[237] = (t[265] & ~t[266]);
  assign t[238] = (t[267] & ~t[268]);
  assign t[239] = (t[269] & ~t[270]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[271] & ~t[272]);
  assign t[241] = (t[273] & ~t[274]);
  assign t[242] = (t[275] & ~t[276]);
  assign t[243] = (t[277] & ~t[278]);
  assign t[244] = (t[279] & ~t[280]);
  assign t[245] = (t[281] & ~t[282]);
  assign t[246] = (t[283] & ~t[284]);
  assign t[247] = (t[285] & ~t[286]);
  assign t[248] = (t[287] & ~t[288]);
  assign t[249] = (t[289] & ~t[290]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[291] & ~t[292]);
  assign t[251] = (t[293] & ~t[294]);
  assign t[252] = (t[295] & ~t[296]);
  assign t[253] = (t[297] & ~t[298]);
  assign t[254] = (t[299] & ~t[300]);
  assign t[255] = (t[301] & ~t[302]);
  assign t[256] = (t[303] & ~t[304]);
  assign t[257] = (t[305] & ~t[306]);
  assign t[258] = (t[307] & ~t[308]);
  assign t[259] = (t[309] & ~t[310]);
  assign t[25] = t[41] ^ t[46];
  assign t[260] = (t[311] & ~t[312]);
  assign t[261] = (t[313] & ~t[314]);
  assign t[262] = (t[315] & ~t[316]);
  assign t[263] = t[317] ^ x[4];
  assign t[264] = t[318] ^ x[3];
  assign t[265] = t[319] ^ x[7];
  assign t[266] = t[320] ^ x[6];
  assign t[267] = t[321] ^ x[12];
  assign t[268] = t[322] ^ x[11];
  assign t[269] = t[323] ^ x[15];
  assign t[26] = t[47] ^ t[48];
  assign t[270] = t[324] ^ x[14];
  assign t[271] = t[325] ^ x[18];
  assign t[272] = t[326] ^ x[17];
  assign t[273] = t[327] ^ x[21];
  assign t[274] = t[328] ^ x[20];
  assign t[275] = t[329] ^ x[24];
  assign t[276] = t[330] ^ x[23];
  assign t[277] = t[331] ^ x[27];
  assign t[278] = t[332] ^ x[26];
  assign t[279] = t[333] ^ x[30];
  assign t[27] = t[49] & t[50];
  assign t[280] = t[334] ^ x[29];
  assign t[281] = t[335] ^ x[33];
  assign t[282] = t[336] ^ x[32];
  assign t[283] = t[337] ^ x[36];
  assign t[284] = t[338] ^ x[35];
  assign t[285] = t[339] ^ x[39];
  assign t[286] = t[340] ^ x[38];
  assign t[287] = t[341] ^ x[42];
  assign t[288] = t[342] ^ x[41];
  assign t[289] = t[343] ^ x[45];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[44];
  assign t[291] = t[345] ^ x[48];
  assign t[292] = t[346] ^ x[47];
  assign t[293] = t[347] ^ x[51];
  assign t[294] = t[348] ^ x[50];
  assign t[295] = t[349] ^ x[54];
  assign t[296] = t[350] ^ x[53];
  assign t[297] = t[351] ^ x[57];
  assign t[298] = t[352] ^ x[56];
  assign t[299] = t[353] ^ x[66];
  assign t[29] = ~(t[184] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[65];
  assign t[301] = t[355] ^ x[71];
  assign t[302] = t[356] ^ x[70];
  assign t[303] = t[357] ^ x[74];
  assign t[304] = t[358] ^ x[73];
  assign t[305] = t[359] ^ x[77];
  assign t[306] = t[360] ^ x[76];
  assign t[307] = t[361] ^ x[80];
  assign t[308] = t[362] ^ x[79];
  assign t[309] = t[363] ^ x[83];
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = t[364] ^ x[82];
  assign t[311] = t[365] ^ x[86];
  assign t[312] = t[366] ^ x[85];
  assign t[313] = t[367] ^ x[105];
  assign t[314] = t[368] ^ x[104];
  assign t[315] = t[369] ^ x[112];
  assign t[316] = t[370] ^ x[111];
  assign t[317] = (x[2]);
  assign t[318] = (x[2]);
  assign t[319] = (x[5]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[5]);
  assign t[321] = (x[10]);
  assign t[322] = (x[10]);
  assign t[323] = (x[13]);
  assign t[324] = (x[13]);
  assign t[325] = (x[16]);
  assign t[326] = (x[16]);
  assign t[327] = (x[19]);
  assign t[328] = (x[19]);
  assign t[329] = (x[22]);
  assign t[32] = ~(t[185]);
  assign t[330] = (x[22]);
  assign t[331] = (x[25]);
  assign t[332] = (x[25]);
  assign t[333] = (x[28]);
  assign t[334] = (x[28]);
  assign t[335] = (x[31]);
  assign t[336] = (x[31]);
  assign t[337] = (x[34]);
  assign t[338] = (x[34]);
  assign t[339] = (x[37]);
  assign t[33] = ~(t[186]);
  assign t[340] = (x[37]);
  assign t[341] = (x[40]);
  assign t[342] = (x[40]);
  assign t[343] = (x[43]);
  assign t[344] = (x[43]);
  assign t[345] = (x[46]);
  assign t[346] = (x[46]);
  assign t[347] = (x[49]);
  assign t[348] = (x[49]);
  assign t[349] = (x[52]);
  assign t[34] = ~(t[187]);
  assign t[350] = (x[52]);
  assign t[351] = (x[55]);
  assign t[352] = (x[55]);
  assign t[353] = (x[64]);
  assign t[354] = (x[64]);
  assign t[355] = (x[69]);
  assign t[356] = (x[69]);
  assign t[357] = (x[72]);
  assign t[358] = (x[72]);
  assign t[359] = (x[75]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[75]);
  assign t[361] = (x[78]);
  assign t[362] = (x[78]);
  assign t[363] = (x[81]);
  assign t[364] = (x[81]);
  assign t[365] = (x[84]);
  assign t[366] = (x[84]);
  assign t[367] = (x[103]);
  assign t[368] = (x[103]);
  assign t[369] = (x[110]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[110]);
  assign t[37] = ~(t[59] ^ t[60]);
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[64];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[65] ? t[66] : t[188];
  assign t[41] = t[65] ? t[67] : t[189];
  assign t[42] = ~(t[68]);
  assign t[43] = t[65] ? t[69] : t[190];
  assign t[44] = t[70] ^ t[63];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = t[73] ^ t[74];
  assign t[47] = t[65] ? t[75] : t[191];
  assign t[48] = t[187] ^ t[76];
  assign t[49] = ~(t[26] ^ t[77]);
  assign t[4] = t[8] ? t[9] : t[182];
  assign t[50] = t[78] ^ t[79];
  assign t[51] = ~(t[80] & t[81]);
  assign t[52] = t[82] ^ t[192];
  assign t[53] = ~(t[184]);
  assign t[54] = t[83] & t[82];
  assign t[55] = ~(t[193]);
  assign t[56] = ~(t[84] & t[194]);
  assign t[57] = t[85] ^ t[86];
  assign t[58] = t[87] ^ t[88];
  assign t[59] = ~(t[89] ^ t[90]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[91] ^ t[92];
  assign t[61] = t[93] ^ t[63];
  assign t[62] = t[94] & t[95];
  assign t[63] = t[96];
  assign t[64] = t[71] ^ t[97];
  assign t[65] = ~(t[98]);
  assign t[66] = t[188] ^ t[99];
  assign t[67] = t[189] ^ t[100];
  assign t[68] = t[65] ? t[101] : t[195];
  assign t[69] = t[190] ^ t[102];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~t[103];
  assign t[71] = t[104] ^ t[62];
  assign t[72] = t[105] & t[106];
  assign t[73] = t[107] ^ t[23];
  assign t[74] = t[108] & t[109];
  assign t[75] = t[191] ^ t[110];
  assign t[76] = t[65] ? t[111] : t[196];
  assign t[77] = t[112] ^ t[88];
  assign t[78] = t[48] ^ t[85];
  assign t[79] = t[197] ^ t[113];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[83] | t[82]);
  assign t[81] = ~(t[114] | t[53]);
  assign t[82] = ~(t[198]);
  assign t[83] = ~(t[192]);
  assign t[84] = ~(t[197]);
  assign t[85] = t[193] ^ t[115];
  assign t[86] = t[77] ^ t[27];
  assign t[87] = t[47] ^ t[85];
  assign t[88] = t[116] & t[79];
  assign t[89] = t[117] ^ t[74];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[118] ^ t[119];
  assign t[91] = t[120] ^ t[118];
  assign t[92] = t[121] ^ t[122];
  assign t[93] = t[123];
  assign t[94] = ~(t[70]);
  assign t[95] = t[124];
  assign t[96] = t[65] ? t[125] : t[199];
  assign t[97] = t[126] & t[127];
  assign t[98] = ~(t[8]);
  assign t[99] = t[128] ? x[59] : x[58];
  assign t[9] = t[182] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [116:0] x;
 output y;

 wire [370:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[31] ? x[61] : x[60];
  assign t[101] = t[195] ^ t[129];
  assign t[102] = t[128] ? x[63] : x[62];
  assign t[103] = t[65] ? t[130] : t[200];
  assign t[104] = t[131] & t[132];
  assign t[105] = ~(t[104] ^ t[133]);
  assign t[106] = t[61] ^ t[134];
  assign t[107] = t[135] & t[136];
  assign t[108] = ~(t[117] ^ t[73]);
  assign t[109] = t[137] ^ t[43];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[138] ? x[68] : x[67];
  assign t[111] = t[196] ^ t[139];
  assign t[112] = t[140] & t[141];
  assign t[113] = t[65] ? t[142] : t[201];
  assign t[114] = ~(t[183]);
  assign t[115] = t[65] ? t[143] : t[202];
  assign t[116] = ~(t[48]);
  assign t[117] = t[40] ^ t[68];
  assign t[118] = t[144] ? t[145] : t[203];
  assign t[119] = t[121] ^ t[146];
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = t[144] ? t[147] : t[204];
  assign t[121] = t[148] ^ t[149];
  assign t[122] = t[150] & t[151];
  assign t[123] = t[65] ? t[152] : t[205];
  assign t[124] = t[65] ? t[153] : t[206];
  assign t[125] = t[199] ^ t[154];
  assign t[126] = ~(t[155] ^ t[71]);
  assign t[127] = t[44] ^ t[95];
  assign t[128] = ~(t[156]);
  assign t[129] = t[128] ? x[88] : x[87];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[200] ^ t[157];
  assign t[131] = ~(t[134]);
  assign t[132] = ~(t[93]);
  assign t[133] = t[44] ^ t[93];
  assign t[134] = t[95] ^ t[70];
  assign t[135] = ~(t[158]);
  assign t[136] = ~(t[40]);
  assign t[137] = t[68] ^ t[41];
  assign t[138] = ~(t[156]);
  assign t[139] = t[138] ? x[90] : x[89];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = ~(t[159]);
  assign t[141] = ~(t[47]);
  assign t[142] = t[201] ^ t[160];
  assign t[143] = t[202] ^ t[161];
  assign t[144] = ~(t[98]);
  assign t[145] = t[203] ^ t[162];
  assign t[146] = t[163] & t[164];
  assign t[147] = t[204] ^ t[165];
  assign t[148] = t[166] & t[167];
  assign t[149] = t[168] & t[169];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = ~(t[148] ^ t[170]);
  assign t[151] = t[171] ^ t[172];
  assign t[152] = t[205] ^ t[173];
  assign t[153] = t[206] ^ t[174];
  assign t[154] = t[31] ? x[92] : x[91];
  assign t[155] = t[93] ^ t[70];
  assign t[156] = ~(t[31]);
  assign t[157] = t[138] ? x[94] : x[93];
  assign t[158] = t[43] ^ t[68];
  assign t[159] = t[79] ^ t[48];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[138] ? x[96] : x[95];
  assign t[161] = t[138] ? x[98] : x[97];
  assign t[162] = t[175] ? x[100] : x[99];
  assign t[163] = ~(t[176] ^ t[121]);
  assign t[164] = t[91] ^ t[169];
  assign t[165] = t[175] ? x[102] : x[101];
  assign t[166] = ~(t[172]);
  assign t[167] = ~(t[177]);
  assign t[168] = ~(t[120]);
  assign t[169] = t[144] ? t[178] : t[207];
  assign t[16] = t[183] | t[30];
  assign t[170] = t[91] ^ t[177];
  assign t[171] = t[177] ^ t[118];
  assign t[172] = t[169] ^ t[120];
  assign t[173] = t[31] ? x[107] : x[106];
  assign t[174] = t[31] ? x[109] : x[108];
  assign t[175] = ~(t[156]);
  assign t[176] = t[177] ^ t[120];
  assign t[177] = t[144] ? t[179] : t[208];
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[208] ^ t[181];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[175] ? x[114] : x[113];
  assign t[181] = t[175] ? x[116] : x[115];
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = t[236] ^ x[4];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[7];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[66];
  assign t[228] = t[255] ^ x[71];
  assign t[229] = t[256] ^ x[74];
  assign t[22] = t[40] ^ t[41];
  assign t[230] = t[257] ^ x[77];
  assign t[231] = t[258] ^ x[80];
  assign t[232] = t[259] ^ x[83];
  assign t[233] = t[260] ^ x[86];
  assign t[234] = t[261] ^ x[105];
  assign t[235] = t[262] ^ x[112];
  assign t[236] = (t[263] & ~t[264]);
  assign t[237] = (t[265] & ~t[266]);
  assign t[238] = (t[267] & ~t[268]);
  assign t[239] = (t[269] & ~t[270]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[271] & ~t[272]);
  assign t[241] = (t[273] & ~t[274]);
  assign t[242] = (t[275] & ~t[276]);
  assign t[243] = (t[277] & ~t[278]);
  assign t[244] = (t[279] & ~t[280]);
  assign t[245] = (t[281] & ~t[282]);
  assign t[246] = (t[283] & ~t[284]);
  assign t[247] = (t[285] & ~t[286]);
  assign t[248] = (t[287] & ~t[288]);
  assign t[249] = (t[289] & ~t[290]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[291] & ~t[292]);
  assign t[251] = (t[293] & ~t[294]);
  assign t[252] = (t[295] & ~t[296]);
  assign t[253] = (t[297] & ~t[298]);
  assign t[254] = (t[299] & ~t[300]);
  assign t[255] = (t[301] & ~t[302]);
  assign t[256] = (t[303] & ~t[304]);
  assign t[257] = (t[305] & ~t[306]);
  assign t[258] = (t[307] & ~t[308]);
  assign t[259] = (t[309] & ~t[310]);
  assign t[25] = t[41] ^ t[46];
  assign t[260] = (t[311] & ~t[312]);
  assign t[261] = (t[313] & ~t[314]);
  assign t[262] = (t[315] & ~t[316]);
  assign t[263] = t[317] ^ x[4];
  assign t[264] = t[318] ^ x[3];
  assign t[265] = t[319] ^ x[7];
  assign t[266] = t[320] ^ x[6];
  assign t[267] = t[321] ^ x[12];
  assign t[268] = t[322] ^ x[11];
  assign t[269] = t[323] ^ x[15];
  assign t[26] = t[47] ^ t[48];
  assign t[270] = t[324] ^ x[14];
  assign t[271] = t[325] ^ x[18];
  assign t[272] = t[326] ^ x[17];
  assign t[273] = t[327] ^ x[21];
  assign t[274] = t[328] ^ x[20];
  assign t[275] = t[329] ^ x[24];
  assign t[276] = t[330] ^ x[23];
  assign t[277] = t[331] ^ x[27];
  assign t[278] = t[332] ^ x[26];
  assign t[279] = t[333] ^ x[30];
  assign t[27] = t[49] & t[50];
  assign t[280] = t[334] ^ x[29];
  assign t[281] = t[335] ^ x[33];
  assign t[282] = t[336] ^ x[32];
  assign t[283] = t[337] ^ x[36];
  assign t[284] = t[338] ^ x[35];
  assign t[285] = t[339] ^ x[39];
  assign t[286] = t[340] ^ x[38];
  assign t[287] = t[341] ^ x[42];
  assign t[288] = t[342] ^ x[41];
  assign t[289] = t[343] ^ x[45];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[44];
  assign t[291] = t[345] ^ x[48];
  assign t[292] = t[346] ^ x[47];
  assign t[293] = t[347] ^ x[51];
  assign t[294] = t[348] ^ x[50];
  assign t[295] = t[349] ^ x[54];
  assign t[296] = t[350] ^ x[53];
  assign t[297] = t[351] ^ x[57];
  assign t[298] = t[352] ^ x[56];
  assign t[299] = t[353] ^ x[66];
  assign t[29] = ~(t[184] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[65];
  assign t[301] = t[355] ^ x[71];
  assign t[302] = t[356] ^ x[70];
  assign t[303] = t[357] ^ x[74];
  assign t[304] = t[358] ^ x[73];
  assign t[305] = t[359] ^ x[77];
  assign t[306] = t[360] ^ x[76];
  assign t[307] = t[361] ^ x[80];
  assign t[308] = t[362] ^ x[79];
  assign t[309] = t[363] ^ x[83];
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = t[364] ^ x[82];
  assign t[311] = t[365] ^ x[86];
  assign t[312] = t[366] ^ x[85];
  assign t[313] = t[367] ^ x[105];
  assign t[314] = t[368] ^ x[104];
  assign t[315] = t[369] ^ x[112];
  assign t[316] = t[370] ^ x[111];
  assign t[317] = (x[2]);
  assign t[318] = (x[2]);
  assign t[319] = (x[5]);
  assign t[31] = ~(t[16]);
  assign t[320] = (x[5]);
  assign t[321] = (x[10]);
  assign t[322] = (x[10]);
  assign t[323] = (x[13]);
  assign t[324] = (x[13]);
  assign t[325] = (x[16]);
  assign t[326] = (x[16]);
  assign t[327] = (x[19]);
  assign t[328] = (x[19]);
  assign t[329] = (x[22]);
  assign t[32] = ~(t[185]);
  assign t[330] = (x[22]);
  assign t[331] = (x[25]);
  assign t[332] = (x[25]);
  assign t[333] = (x[28]);
  assign t[334] = (x[28]);
  assign t[335] = (x[31]);
  assign t[336] = (x[31]);
  assign t[337] = (x[34]);
  assign t[338] = (x[34]);
  assign t[339] = (x[37]);
  assign t[33] = ~(t[186]);
  assign t[340] = (x[37]);
  assign t[341] = (x[40]);
  assign t[342] = (x[40]);
  assign t[343] = (x[43]);
  assign t[344] = (x[43]);
  assign t[345] = (x[46]);
  assign t[346] = (x[46]);
  assign t[347] = (x[49]);
  assign t[348] = (x[49]);
  assign t[349] = (x[52]);
  assign t[34] = ~(t[187]);
  assign t[350] = (x[52]);
  assign t[351] = (x[55]);
  assign t[352] = (x[55]);
  assign t[353] = (x[64]);
  assign t[354] = (x[64]);
  assign t[355] = (x[69]);
  assign t[356] = (x[69]);
  assign t[357] = (x[72]);
  assign t[358] = (x[72]);
  assign t[359] = (x[75]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[75]);
  assign t[361] = (x[78]);
  assign t[362] = (x[78]);
  assign t[363] = (x[81]);
  assign t[364] = (x[81]);
  assign t[365] = (x[84]);
  assign t[366] = (x[84]);
  assign t[367] = (x[103]);
  assign t[368] = (x[103]);
  assign t[369] = (x[110]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[110]);
  assign t[37] = ~(t[59] ^ t[60]);
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[64];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[65] ? t[66] : t[188];
  assign t[41] = t[65] ? t[67] : t[189];
  assign t[42] = ~(t[68]);
  assign t[43] = t[65] ? t[69] : t[190];
  assign t[44] = t[70] ^ t[63];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = t[73] ^ t[74];
  assign t[47] = t[65] ? t[75] : t[191];
  assign t[48] = t[187] ^ t[76];
  assign t[49] = ~(t[26] ^ t[77]);
  assign t[4] = t[8] ? t[9] : t[182];
  assign t[50] = t[78] ^ t[79];
  assign t[51] = ~(t[80] & t[81]);
  assign t[52] = t[82] ^ t[192];
  assign t[53] = ~(t[184]);
  assign t[54] = t[83] & t[82];
  assign t[55] = ~(t[193]);
  assign t[56] = ~(t[84] & t[194]);
  assign t[57] = t[85] ^ t[86];
  assign t[58] = t[87] ^ t[88];
  assign t[59] = ~(t[89] ^ t[90]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[91] ^ t[92];
  assign t[61] = t[93] ^ t[63];
  assign t[62] = t[94] & t[95];
  assign t[63] = t[96];
  assign t[64] = t[71] ^ t[97];
  assign t[65] = ~(t[98]);
  assign t[66] = t[188] ^ t[99];
  assign t[67] = t[189] ^ t[100];
  assign t[68] = t[65] ? t[101] : t[195];
  assign t[69] = t[190] ^ t[102];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~t[103];
  assign t[71] = t[104] ^ t[62];
  assign t[72] = t[105] & t[106];
  assign t[73] = t[107] ^ t[23];
  assign t[74] = t[108] & t[109];
  assign t[75] = t[191] ^ t[110];
  assign t[76] = t[65] ? t[111] : t[196];
  assign t[77] = t[112] ^ t[88];
  assign t[78] = t[48] ^ t[85];
  assign t[79] = t[197] ^ t[113];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[83] | t[82]);
  assign t[81] = ~(t[114] | t[53]);
  assign t[82] = ~(t[198]);
  assign t[83] = ~(t[192]);
  assign t[84] = ~(t[197]);
  assign t[85] = t[193] ^ t[115];
  assign t[86] = t[77] ^ t[27];
  assign t[87] = t[47] ^ t[85];
  assign t[88] = t[116] & t[79];
  assign t[89] = t[117] ^ t[74];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[118] ^ t[119];
  assign t[91] = t[120] ^ t[118];
  assign t[92] = t[121] ^ t[122];
  assign t[93] = t[123];
  assign t[94] = ~(t[70]);
  assign t[95] = t[124];
  assign t[96] = t[65] ? t[125] : t[199];
  assign t[97] = t[126] & t[127];
  assign t[98] = ~(t[8]);
  assign t[99] = t[128] ? x[59] : x[58];
  assign t[9] = t[182] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [116:0] x;
 output y;

 wire [361:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[133] & t[134];
  assign t[101] = ~(t[8]);
  assign t[102] = t[135] ? x[68] : x[67];
  assign t[103] = t[135] ? x[70] : x[69];
  assign t[104] = t[136] & t[137];
  assign t[105] = t[138] & t[71];
  assign t[106] = t[66] ? t[139] : t[194];
  assign t[107] = t[186] ^ t[140];
  assign t[108] = t[187] ^ t[141];
  assign t[109] = t[188] ^ t[142];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[116]);
  assign t[111] = ~(t[92]);
  assign t[112] = ~(t[44]);
  assign t[113] = t[190] ^ t[143];
  assign t[114] = t[24] ^ t[92];
  assign t[115] = t[92] ^ t[45];
  assign t[116] = t[113] ^ t[44];
  assign t[117] = t[87] ? x[75] : x[74];
  assign t[118] = ~(t[144]);
  assign t[119] = ~(t[129]);
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = ~(t[130]);
  assign t[121] = t[145];
  assign t[122] = t[130] ^ t[26];
  assign t[123] = ~(t[174]);
  assign t[124] = t[191] ^ t[146];
  assign t[125] = t[97] ? t[147] : t[195];
  assign t[126] = t[192] ^ t[148];
  assign t[127] = t[193] ^ t[149];
  assign t[128] = t[150] & t[151];
  assign t[129] = t[152];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = ~t[153];
  assign t[131] = t[154] ? x[80] : x[79];
  assign t[132] = t[155] & t[156];
  assign t[133] = ~(t[157] ^ t[99]);
  assign t[134] = t[158] ^ t[91];
  assign t[135] = ~(t[55]);
  assign t[136] = ~(t[159]);
  assign t[137] = ~(t[40]);
  assign t[138] = ~(t[41]);
  assign t[139] = t[194] ^ t[160];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[135] ? x[82] : x[81];
  assign t[141] = t[31] ? x[84] : x[83];
  assign t[142] = t[31] ? x[86] : x[85];
  assign t[143] = t[66] ? t[161] : t[196];
  assign t[144] = t[121] ^ t[130];
  assign t[145] = t[66] ? t[162] : t[197];
  assign t[146] = t[154] ? x[94] : x[93];
  assign t[147] = t[195] ^ t[163];
  assign t[148] = t[154] ? x[96] : x[95];
  assign t[149] = t[31] ? x[98] : x[97];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = ~(t[104] ^ t[164]);
  assign t[151] = t[165] ^ t[159];
  assign t[152] = t[66] ? t[166] : t[198];
  assign t[153] = t[66] ? t[167] : t[199];
  assign t[154] = ~(t[55]);
  assign t[155] = ~(t[168]);
  assign t[156] = ~(t[89]);
  assign t[157] = t[89] ^ t[125];
  assign t[158] = t[125] ^ t[64];
  assign t[159] = t[71] ^ t[41];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[87] ? x[106] : x[105];
  assign t[161] = t[196] ^ t[169];
  assign t[162] = t[197] ^ t[170];
  assign t[163] = t[154] ? x[108] : x[107];
  assign t[164] = t[70] ^ t[40];
  assign t[165] = t[40] ^ t[106];
  assign t[166] = t[198] ^ t[171];
  assign t[167] = t[199] ^ t[172];
  assign t[168] = t[91] ^ t[125];
  assign t[169] = t[31] ? x[110] : x[109];
  assign t[16] = t[174] | t[30];
  assign t[170] = t[87] ? x[112] : x[111];
  assign t[171] = t[87] ? x[114] : x[113];
  assign t[172] = t[31] ? x[116] : x[115];
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[4];
  assign t[201] = t[228] ^ x[7];
  assign t[202] = t[229] ^ x[12];
  assign t[203] = t[230] ^ x[15];
  assign t[204] = t[231] ^ x[18];
  assign t[205] = t[232] ^ x[21];
  assign t[206] = t[233] ^ x[24];
  assign t[207] = t[234] ^ x[27];
  assign t[208] = t[235] ^ x[30];
  assign t[209] = t[236] ^ x[33];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[36];
  assign t[211] = t[238] ^ x[39];
  assign t[212] = t[239] ^ x[42];
  assign t[213] = t[240] ^ x[45];
  assign t[214] = t[241] ^ x[48];
  assign t[215] = t[242] ^ x[51];
  assign t[216] = t[243] ^ x[54];
  assign t[217] = t[244] ^ x[57];
  assign t[218] = t[245] ^ x[60];
  assign t[219] = t[246] ^ x[63];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[66];
  assign t[221] = t[248] ^ x[73];
  assign t[222] = t[249] ^ x[78];
  assign t[223] = t[250] ^ x[89];
  assign t[224] = t[251] ^ x[92];
  assign t[225] = t[252] ^ x[101];
  assign t[226] = t[253] ^ x[104];
  assign t[227] = (t[254] & ~t[255]);
  assign t[228] = (t[256] & ~t[257]);
  assign t[229] = (t[258] & ~t[259]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[260] & ~t[261]);
  assign t[231] = (t[262] & ~t[263]);
  assign t[232] = (t[264] & ~t[265]);
  assign t[233] = (t[266] & ~t[267]);
  assign t[234] = (t[268] & ~t[269]);
  assign t[235] = (t[270] & ~t[271]);
  assign t[236] = (t[272] & ~t[273]);
  assign t[237] = (t[274] & ~t[275]);
  assign t[238] = (t[276] & ~t[277]);
  assign t[239] = (t[278] & ~t[279]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[280] & ~t[281]);
  assign t[241] = (t[282] & ~t[283]);
  assign t[242] = (t[284] & ~t[285]);
  assign t[243] = (t[286] & ~t[287]);
  assign t[244] = (t[288] & ~t[289]);
  assign t[245] = (t[290] & ~t[291]);
  assign t[246] = (t[292] & ~t[293]);
  assign t[247] = (t[294] & ~t[295]);
  assign t[248] = (t[296] & ~t[297]);
  assign t[249] = (t[298] & ~t[299]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[300] & ~t[301]);
  assign t[251] = (t[302] & ~t[303]);
  assign t[252] = (t[304] & ~t[305]);
  assign t[253] = (t[306] & ~t[307]);
  assign t[254] = t[308] ^ x[4];
  assign t[255] = t[309] ^ x[3];
  assign t[256] = t[310] ^ x[7];
  assign t[257] = t[311] ^ x[6];
  assign t[258] = t[312] ^ x[12];
  assign t[259] = t[313] ^ x[11];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[314] ^ x[15];
  assign t[261] = t[315] ^ x[14];
  assign t[262] = t[316] ^ x[18];
  assign t[263] = t[317] ^ x[17];
  assign t[264] = t[318] ^ x[21];
  assign t[265] = t[319] ^ x[20];
  assign t[266] = t[320] ^ x[24];
  assign t[267] = t[321] ^ x[23];
  assign t[268] = t[322] ^ x[27];
  assign t[269] = t[323] ^ x[26];
  assign t[26] = t[48];
  assign t[270] = t[324] ^ x[30];
  assign t[271] = t[325] ^ x[29];
  assign t[272] = t[326] ^ x[33];
  assign t[273] = t[327] ^ x[32];
  assign t[274] = t[328] ^ x[36];
  assign t[275] = t[329] ^ x[35];
  assign t[276] = t[330] ^ x[39];
  assign t[277] = t[331] ^ x[38];
  assign t[278] = t[332] ^ x[42];
  assign t[279] = t[333] ^ x[41];
  assign t[27] = t[49] ^ t[50];
  assign t[280] = t[334] ^ x[45];
  assign t[281] = t[335] ^ x[44];
  assign t[282] = t[336] ^ x[48];
  assign t[283] = t[337] ^ x[47];
  assign t[284] = t[338] ^ x[51];
  assign t[285] = t[339] ^ x[50];
  assign t[286] = t[340] ^ x[54];
  assign t[287] = t[341] ^ x[53];
  assign t[288] = t[342] ^ x[57];
  assign t[289] = t[343] ^ x[56];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[60];
  assign t[291] = t[345] ^ x[59];
  assign t[292] = t[346] ^ x[63];
  assign t[293] = t[347] ^ x[62];
  assign t[294] = t[348] ^ x[66];
  assign t[295] = t[349] ^ x[65];
  assign t[296] = t[350] ^ x[73];
  assign t[297] = t[351] ^ x[72];
  assign t[298] = t[352] ^ x[78];
  assign t[299] = t[353] ^ x[77];
  assign t[29] = ~(t[175] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[89];
  assign t[301] = t[355] ^ x[88];
  assign t[302] = t[356] ^ x[92];
  assign t[303] = t[357] ^ x[91];
  assign t[304] = t[358] ^ x[101];
  assign t[305] = t[359] ^ x[100];
  assign t[306] = t[360] ^ x[104];
  assign t[307] = t[361] ^ x[103];
  assign t[308] = (x[2]);
  assign t[309] = (x[2]);
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = (x[5]);
  assign t[311] = (x[5]);
  assign t[312] = (x[10]);
  assign t[313] = (x[10]);
  assign t[314] = (x[13]);
  assign t[315] = (x[13]);
  assign t[316] = (x[16]);
  assign t[317] = (x[16]);
  assign t[318] = (x[19]);
  assign t[319] = (x[19]);
  assign t[31] = ~(t[55]);
  assign t[320] = (x[22]);
  assign t[321] = (x[22]);
  assign t[322] = (x[25]);
  assign t[323] = (x[25]);
  assign t[324] = (x[28]);
  assign t[325] = (x[28]);
  assign t[326] = (x[31]);
  assign t[327] = (x[31]);
  assign t[328] = (x[34]);
  assign t[329] = (x[34]);
  assign t[32] = ~(t[176]);
  assign t[330] = (x[37]);
  assign t[331] = (x[37]);
  assign t[332] = (x[40]);
  assign t[333] = (x[40]);
  assign t[334] = (x[43]);
  assign t[335] = (x[43]);
  assign t[336] = (x[46]);
  assign t[337] = (x[46]);
  assign t[338] = (x[49]);
  assign t[339] = (x[49]);
  assign t[33] = ~(t[177]);
  assign t[340] = (x[52]);
  assign t[341] = (x[52]);
  assign t[342] = (x[55]);
  assign t[343] = (x[55]);
  assign t[344] = (x[58]);
  assign t[345] = (x[58]);
  assign t[346] = (x[61]);
  assign t[347] = (x[61]);
  assign t[348] = (x[64]);
  assign t[349] = (x[64]);
  assign t[34] = ~(t[178]);
  assign t[350] = (x[71]);
  assign t[351] = (x[71]);
  assign t[352] = (x[76]);
  assign t[353] = (x[76]);
  assign t[354] = (x[87]);
  assign t[355] = (x[87]);
  assign t[356] = (x[90]);
  assign t[357] = (x[90]);
  assign t[358] = (x[99]);
  assign t[359] = (x[99]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = (x[102]);
  assign t[361] = (x[102]);
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[62] ^ t[63];
  assign t[39] = t[64] ^ t[65];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[66] ? t[67] : t[179];
  assign t[41] = t[66] ? t[68] : t[180];
  assign t[42] = ~(t[22] ^ t[69]);
  assign t[43] = t[70] ^ t[71];
  assign t[44] = t[178] ^ t[72];
  assign t[45] = t[181] ^ t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = t[76] & t[77];
  assign t[48] = t[66] ? t[78] : t[182];
  assign t[49] = t[79] ^ t[80];
  assign t[4] = t[8] ? t[9] : t[173];
  assign t[50] = t[81] & t[82];
  assign t[51] = ~(t[83] & t[84]);
  assign t[52] = t[85] ^ t[183];
  assign t[53] = ~(t[175]);
  assign t[54] = t[86] & t[85];
  assign t[55] = ~(t[87]);
  assign t[56] = ~(t[181]);
  assign t[57] = ~(t[88] & t[184]);
  assign t[58] = t[89] ^ t[64];
  assign t[59] = t[90] & t[91];
  assign t[5] = ~(t[10]);
  assign t[60] = t[92] ^ t[44];
  assign t[61] = t[93] & t[94];
  assign t[62] = t[70] ^ t[95];
  assign t[63] = t[96] ^ t[50];
  assign t[64] = t[97] ? t[98] : t[185];
  assign t[65] = t[99] ^ t[100];
  assign t[66] = ~(t[101]);
  assign t[67] = t[179] ^ t[102];
  assign t[68] = t[180] ^ t[103];
  assign t[69] = t[104] ^ t[105];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[41] ^ t[106];
  assign t[71] = t[66] ? t[107] : t[186];
  assign t[72] = t[66] ? t[108] : t[187];
  assign t[73] = t[66] ? t[109] : t[188];
  assign t[74] = t[110] & t[111];
  assign t[75] = t[112] & t[113];
  assign t[76] = ~(t[74] ^ t[114]);
  assign t[77] = t[115] ^ t[116];
  assign t[78] = t[182] ^ t[117];
  assign t[79] = t[118] & t[119];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[120] & t[121];
  assign t[81] = ~(t[96] ^ t[49]);
  assign t[82] = t[122] ^ t[121];
  assign t[83] = ~(t[86] | t[85]);
  assign t[84] = ~(t[123] | t[53]);
  assign t[85] = ~(t[189]);
  assign t[86] = ~(t[183]);
  assign t[87] = ~(t[16]);
  assign t[88] = ~(t[190]);
  assign t[89] = t[97] ? t[124] : t[191];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = ~(t[125]);
  assign t[91] = t[97] ? t[126] : t[192];
  assign t[92] = t[66] ? t[127] : t[193];
  assign t[93] = ~(t[60] ^ t[46]);
  assign t[94] = t[24] ^ t[113];
  assign t[95] = t[69] ^ t[128];
  assign t[96] = t[129] ^ t[130];
  assign t[97] = ~(t[101]);
  assign t[98] = t[185] ^ t[131];
  assign t[99] = t[132] ^ t[59];
  assign t[9] = t[173] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [116:0] x;
 output y;

 wire [361:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[133] & t[134];
  assign t[101] = ~(t[8]);
  assign t[102] = t[135] ? x[68] : x[67];
  assign t[103] = t[135] ? x[70] : x[69];
  assign t[104] = t[136] & t[137];
  assign t[105] = t[138] & t[71];
  assign t[106] = t[66] ? t[139] : t[194];
  assign t[107] = t[186] ^ t[140];
  assign t[108] = t[187] ^ t[141];
  assign t[109] = t[188] ^ t[142];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = ~(t[116]);
  assign t[111] = ~(t[92]);
  assign t[112] = ~(t[44]);
  assign t[113] = t[190] ^ t[143];
  assign t[114] = t[24] ^ t[92];
  assign t[115] = t[92] ^ t[45];
  assign t[116] = t[113] ^ t[44];
  assign t[117] = t[87] ? x[75] : x[74];
  assign t[118] = ~(t[144]);
  assign t[119] = ~(t[129]);
  assign t[11] = ~(t[20] ^ t[21]);
  assign t[120] = ~(t[130]);
  assign t[121] = t[145];
  assign t[122] = t[130] ^ t[26];
  assign t[123] = ~(t[174]);
  assign t[124] = t[191] ^ t[146];
  assign t[125] = t[97] ? t[147] : t[195];
  assign t[126] = t[192] ^ t[148];
  assign t[127] = t[193] ^ t[149];
  assign t[128] = t[150] & t[151];
  assign t[129] = t[152];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = ~t[153];
  assign t[131] = t[154] ? x[80] : x[79];
  assign t[132] = t[155] & t[156];
  assign t[133] = ~(t[157] ^ t[99]);
  assign t[134] = t[158] ^ t[91];
  assign t[135] = ~(t[55]);
  assign t[136] = ~(t[159]);
  assign t[137] = ~(t[40]);
  assign t[138] = ~(t[41]);
  assign t[139] = t[194] ^ t[160];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[135] ? x[82] : x[81];
  assign t[141] = t[31] ? x[84] : x[83];
  assign t[142] = t[31] ? x[86] : x[85];
  assign t[143] = t[66] ? t[161] : t[196];
  assign t[144] = t[121] ^ t[130];
  assign t[145] = t[66] ? t[162] : t[197];
  assign t[146] = t[154] ? x[94] : x[93];
  assign t[147] = t[195] ^ t[163];
  assign t[148] = t[154] ? x[96] : x[95];
  assign t[149] = t[31] ? x[98] : x[97];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = ~(t[104] ^ t[164]);
  assign t[151] = t[165] ^ t[159];
  assign t[152] = t[66] ? t[166] : t[198];
  assign t[153] = t[66] ? t[167] : t[199];
  assign t[154] = ~(t[55]);
  assign t[155] = ~(t[168]);
  assign t[156] = ~(t[89]);
  assign t[157] = t[89] ^ t[125];
  assign t[158] = t[125] ^ t[64];
  assign t[159] = t[71] ^ t[41];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[87] ? x[106] : x[105];
  assign t[161] = t[196] ^ t[169];
  assign t[162] = t[197] ^ t[170];
  assign t[163] = t[154] ? x[108] : x[107];
  assign t[164] = t[70] ^ t[40];
  assign t[165] = t[40] ^ t[106];
  assign t[166] = t[198] ^ t[171];
  assign t[167] = t[199] ^ t[172];
  assign t[168] = t[91] ^ t[125];
  assign t[169] = t[31] ? x[110] : x[109];
  assign t[16] = t[174] | t[30];
  assign t[170] = t[87] ? x[112] : x[111];
  assign t[171] = t[87] ? x[114] : x[113];
  assign t[172] = t[31] ? x[116] : x[115];
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[4];
  assign t[201] = t[228] ^ x[7];
  assign t[202] = t[229] ^ x[12];
  assign t[203] = t[230] ^ x[15];
  assign t[204] = t[231] ^ x[18];
  assign t[205] = t[232] ^ x[21];
  assign t[206] = t[233] ^ x[24];
  assign t[207] = t[234] ^ x[27];
  assign t[208] = t[235] ^ x[30];
  assign t[209] = t[236] ^ x[33];
  assign t[20] = t[36] ^ t[37];
  assign t[210] = t[237] ^ x[36];
  assign t[211] = t[238] ^ x[39];
  assign t[212] = t[239] ^ x[42];
  assign t[213] = t[240] ^ x[45];
  assign t[214] = t[241] ^ x[48];
  assign t[215] = t[242] ^ x[51];
  assign t[216] = t[243] ^ x[54];
  assign t[217] = t[244] ^ x[57];
  assign t[218] = t[245] ^ x[60];
  assign t[219] = t[246] ^ x[63];
  assign t[21] = ~(t[38] ^ t[39]);
  assign t[220] = t[247] ^ x[66];
  assign t[221] = t[248] ^ x[73];
  assign t[222] = t[249] ^ x[78];
  assign t[223] = t[250] ^ x[89];
  assign t[224] = t[251] ^ x[92];
  assign t[225] = t[252] ^ x[101];
  assign t[226] = t[253] ^ x[104];
  assign t[227] = (t[254] & ~t[255]);
  assign t[228] = (t[256] & ~t[257]);
  assign t[229] = (t[258] & ~t[259]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[260] & ~t[261]);
  assign t[231] = (t[262] & ~t[263]);
  assign t[232] = (t[264] & ~t[265]);
  assign t[233] = (t[266] & ~t[267]);
  assign t[234] = (t[268] & ~t[269]);
  assign t[235] = (t[270] & ~t[271]);
  assign t[236] = (t[272] & ~t[273]);
  assign t[237] = (t[274] & ~t[275]);
  assign t[238] = (t[276] & ~t[277]);
  assign t[239] = (t[278] & ~t[279]);
  assign t[23] = t[42] & t[43];
  assign t[240] = (t[280] & ~t[281]);
  assign t[241] = (t[282] & ~t[283]);
  assign t[242] = (t[284] & ~t[285]);
  assign t[243] = (t[286] & ~t[287]);
  assign t[244] = (t[288] & ~t[289]);
  assign t[245] = (t[290] & ~t[291]);
  assign t[246] = (t[292] & ~t[293]);
  assign t[247] = (t[294] & ~t[295]);
  assign t[248] = (t[296] & ~t[297]);
  assign t[249] = (t[298] & ~t[299]);
  assign t[24] = t[44] ^ t[45];
  assign t[250] = (t[300] & ~t[301]);
  assign t[251] = (t[302] & ~t[303]);
  assign t[252] = (t[304] & ~t[305]);
  assign t[253] = (t[306] & ~t[307]);
  assign t[254] = t[308] ^ x[4];
  assign t[255] = t[309] ^ x[3];
  assign t[256] = t[310] ^ x[7];
  assign t[257] = t[311] ^ x[6];
  assign t[258] = t[312] ^ x[12];
  assign t[259] = t[313] ^ x[11];
  assign t[25] = t[46] ^ t[47];
  assign t[260] = t[314] ^ x[15];
  assign t[261] = t[315] ^ x[14];
  assign t[262] = t[316] ^ x[18];
  assign t[263] = t[317] ^ x[17];
  assign t[264] = t[318] ^ x[21];
  assign t[265] = t[319] ^ x[20];
  assign t[266] = t[320] ^ x[24];
  assign t[267] = t[321] ^ x[23];
  assign t[268] = t[322] ^ x[27];
  assign t[269] = t[323] ^ x[26];
  assign t[26] = t[48];
  assign t[270] = t[324] ^ x[30];
  assign t[271] = t[325] ^ x[29];
  assign t[272] = t[326] ^ x[33];
  assign t[273] = t[327] ^ x[32];
  assign t[274] = t[328] ^ x[36];
  assign t[275] = t[329] ^ x[35];
  assign t[276] = t[330] ^ x[39];
  assign t[277] = t[331] ^ x[38];
  assign t[278] = t[332] ^ x[42];
  assign t[279] = t[333] ^ x[41];
  assign t[27] = t[49] ^ t[50];
  assign t[280] = t[334] ^ x[45];
  assign t[281] = t[335] ^ x[44];
  assign t[282] = t[336] ^ x[48];
  assign t[283] = t[337] ^ x[47];
  assign t[284] = t[338] ^ x[51];
  assign t[285] = t[339] ^ x[50];
  assign t[286] = t[340] ^ x[54];
  assign t[287] = t[341] ^ x[53];
  assign t[288] = t[342] ^ x[57];
  assign t[289] = t[343] ^ x[56];
  assign t[28] = ~(t[30] & t[51]);
  assign t[290] = t[344] ^ x[60];
  assign t[291] = t[345] ^ x[59];
  assign t[292] = t[346] ^ x[63];
  assign t[293] = t[347] ^ x[62];
  assign t[294] = t[348] ^ x[66];
  assign t[295] = t[349] ^ x[65];
  assign t[296] = t[350] ^ x[73];
  assign t[297] = t[351] ^ x[72];
  assign t[298] = t[352] ^ x[78];
  assign t[299] = t[353] ^ x[77];
  assign t[29] = ~(t[175] ^ t[52]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[89];
  assign t[301] = t[355] ^ x[88];
  assign t[302] = t[356] ^ x[92];
  assign t[303] = t[357] ^ x[91];
  assign t[304] = t[358] ^ x[101];
  assign t[305] = t[359] ^ x[100];
  assign t[306] = t[360] ^ x[104];
  assign t[307] = t[361] ^ x[103];
  assign t[308] = (x[2]);
  assign t[309] = (x[2]);
  assign t[30] = ~(t[53] & t[54]);
  assign t[310] = (x[5]);
  assign t[311] = (x[5]);
  assign t[312] = (x[10]);
  assign t[313] = (x[10]);
  assign t[314] = (x[13]);
  assign t[315] = (x[13]);
  assign t[316] = (x[16]);
  assign t[317] = (x[16]);
  assign t[318] = (x[19]);
  assign t[319] = (x[19]);
  assign t[31] = ~(t[55]);
  assign t[320] = (x[22]);
  assign t[321] = (x[22]);
  assign t[322] = (x[25]);
  assign t[323] = (x[25]);
  assign t[324] = (x[28]);
  assign t[325] = (x[28]);
  assign t[326] = (x[31]);
  assign t[327] = (x[31]);
  assign t[328] = (x[34]);
  assign t[329] = (x[34]);
  assign t[32] = ~(t[176]);
  assign t[330] = (x[37]);
  assign t[331] = (x[37]);
  assign t[332] = (x[40]);
  assign t[333] = (x[40]);
  assign t[334] = (x[43]);
  assign t[335] = (x[43]);
  assign t[336] = (x[46]);
  assign t[337] = (x[46]);
  assign t[338] = (x[49]);
  assign t[339] = (x[49]);
  assign t[33] = ~(t[177]);
  assign t[340] = (x[52]);
  assign t[341] = (x[52]);
  assign t[342] = (x[55]);
  assign t[343] = (x[55]);
  assign t[344] = (x[58]);
  assign t[345] = (x[58]);
  assign t[346] = (x[61]);
  assign t[347] = (x[61]);
  assign t[348] = (x[64]);
  assign t[349] = (x[64]);
  assign t[34] = ~(t[178]);
  assign t[350] = (x[71]);
  assign t[351] = (x[71]);
  assign t[352] = (x[76]);
  assign t[353] = (x[76]);
  assign t[354] = (x[87]);
  assign t[355] = (x[87]);
  assign t[356] = (x[90]);
  assign t[357] = (x[90]);
  assign t[358] = (x[99]);
  assign t[359] = (x[99]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = (x[102]);
  assign t[361] = (x[102]);
  assign t[36] = t[58] ^ t[59];
  assign t[37] = t[60] ^ t[61];
  assign t[38] = t[62] ^ t[63];
  assign t[39] = t[64] ^ t[65];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[66] ? t[67] : t[179];
  assign t[41] = t[66] ? t[68] : t[180];
  assign t[42] = ~(t[22] ^ t[69]);
  assign t[43] = t[70] ^ t[71];
  assign t[44] = t[178] ^ t[72];
  assign t[45] = t[181] ^ t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = t[76] & t[77];
  assign t[48] = t[66] ? t[78] : t[182];
  assign t[49] = t[79] ^ t[80];
  assign t[4] = t[8] ? t[9] : t[173];
  assign t[50] = t[81] & t[82];
  assign t[51] = ~(t[83] & t[84]);
  assign t[52] = t[85] ^ t[183];
  assign t[53] = ~(t[175]);
  assign t[54] = t[86] & t[85];
  assign t[55] = ~(t[87]);
  assign t[56] = ~(t[181]);
  assign t[57] = ~(t[88] & t[184]);
  assign t[58] = t[89] ^ t[64];
  assign t[59] = t[90] & t[91];
  assign t[5] = ~(t[10]);
  assign t[60] = t[92] ^ t[44];
  assign t[61] = t[93] & t[94];
  assign t[62] = t[70] ^ t[95];
  assign t[63] = t[96] ^ t[50];
  assign t[64] = t[97] ? t[98] : t[185];
  assign t[65] = t[99] ^ t[100];
  assign t[66] = ~(t[101]);
  assign t[67] = t[179] ^ t[102];
  assign t[68] = t[180] ^ t[103];
  assign t[69] = t[104] ^ t[105];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[41] ^ t[106];
  assign t[71] = t[66] ? t[107] : t[186];
  assign t[72] = t[66] ? t[108] : t[187];
  assign t[73] = t[66] ? t[109] : t[188];
  assign t[74] = t[110] & t[111];
  assign t[75] = t[112] & t[113];
  assign t[76] = ~(t[74] ^ t[114]);
  assign t[77] = t[115] ^ t[116];
  assign t[78] = t[182] ^ t[117];
  assign t[79] = t[118] & t[119];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[120] & t[121];
  assign t[81] = ~(t[96] ^ t[49]);
  assign t[82] = t[122] ^ t[121];
  assign t[83] = ~(t[86] | t[85]);
  assign t[84] = ~(t[123] | t[53]);
  assign t[85] = ~(t[189]);
  assign t[86] = ~(t[183]);
  assign t[87] = ~(t[16]);
  assign t[88] = ~(t[190]);
  assign t[89] = t[97] ? t[124] : t[191];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = ~(t[125]);
  assign t[91] = t[97] ? t[126] : t[192];
  assign t[92] = t[66] ? t[127] : t[193];
  assign t[93] = ~(t[60] ^ t[46]);
  assign t[94] = t[24] ^ t[113];
  assign t[95] = t[69] ^ t[128];
  assign t[96] = t[129] ^ t[130];
  assign t[97] = ~(t[101]);
  assign t[98] = t[185] ^ t[131];
  assign t[99] = t[132] ^ t[59];
  assign t[9] = t[173] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [116:0] x;
 output y;

 wire [360:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[130]);
  assign t[101] = ~(t[129]);
  assign t[102] = ~(t[131]);
  assign t[103] = ~(t[66]);
  assign t[104] = t[8] ? t[132] : t[191];
  assign t[105] = t[131] ^ t[66];
  assign t[106] = ~(t[133] & t[134]);
  assign t[107] = t[135] ^ t[192];
  assign t[108] = ~(t[186]);
  assign t[109] = t[136] & t[135];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[28] ? x[72] : x[71];
  assign t[111] = t[188] ^ t[137];
  assign t[112] = t[138] ? x[74] : x[73];
  assign t[113] = t[138] ? x[76] : x[75];
  assign t[114] = t[28] ? x[78] : x[77];
  assign t[115] = ~t[139];
  assign t[116] = t[27] ? t[140] : t[193];
  assign t[117] = t[141] ^ t[20];
  assign t[118] = t[142] & t[143];
  assign t[119] = t[144] & t[145];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[15]);
  assign t[121] = t[189] ^ t[146];
  assign t[122] = t[190] ^ t[147];
  assign t[123] = t[148] ^ t[149];
  assign t[124] = t[94] ^ t[150];
  assign t[125] = t[120] ? t[151] : t[194];
  assign t[126] = t[100] ? x[86] : x[85];
  assign t[127] = t[43] ^ t[131];
  assign t[128] = t[131] ^ t[25];
  assign t[129] = t[104] ^ t[66];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = ~(t[28]);
  assign t[131] = t[8] ? t[152] : t[195];
  assign t[132] = t[191] ^ t[153];
  assign t[133] = ~(t[136] | t[135]);
  assign t[134] = ~(t[154] | t[108]);
  assign t[135] = ~(t[196]);
  assign t[136] = ~(t[192]);
  assign t[137] = t[138] ? x[94] : x[93];
  assign t[138] = ~(t[130]);
  assign t[139] = t[27] ? t[155] : t[197];
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[193] ^ t[156];
  assign t[141] = t[157] & t[158];
  assign t[142] = ~(t[141] ^ t[159]);
  assign t[143] = t[19] ^ t[160];
  assign t[144] = ~(t[161] ^ t[39]);
  assign t[145] = t[21] ^ t[86];
  assign t[146] = t[162] ? x[99] : x[98];
  assign t[147] = t[162] ? x[101] : x[100];
  assign t[148] = t[163] & t[164];
  assign t[149] = t[165] & t[125];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[120] ? t[166] : t[198];
  assign t[151] = t[194] ^ t[167];
  assign t[152] = t[195] ^ t[168];
  assign t[153] = t[100] ? x[106] : x[105];
  assign t[154] = ~(t[179]);
  assign t[155] = t[197] ^ t[169];
  assign t[156] = t[100] ? x[108] : x[107];
  assign t[157] = ~(t[160]);
  assign t[158] = ~(t[33]);
  assign t[159] = t[90] ^ t[33];
  assign t[15] = ~(t[27]);
  assign t[160] = t[36] ^ t[54];
  assign t[161] = t[115] ^ t[37];
  assign t[162] = ~(t[130]);
  assign t[163] = ~(t[170]);
  assign t[164] = ~(t[93]);
  assign t[165] = ~(t[94]);
  assign t[166] = t[198] ^ t[171];
  assign t[167] = t[162] ? x[110] : x[109];
  assign t[168] = t[100] ? x[112] : x[111];
  assign t[169] = t[28] ? x[114] : x[113];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[125] ^ t[94];
  assign t[171] = t[162] ? x[116] : x[115];
  assign t[172] = (t[199]);
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = t[226] ^ x[4];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[9];
  assign t[201] = t[228] ^ x[12];
  assign t[202] = t[229] ^ x[15];
  assign t[203] = t[230] ^ x[18];
  assign t[204] = t[231] ^ x[21];
  assign t[205] = t[232] ^ x[24];
  assign t[206] = t[233] ^ x[27];
  assign t[207] = t[234] ^ x[30];
  assign t[208] = t[235] ^ x[33];
  assign t[209] = t[236] ^ x[36];
  assign t[20] = t[35] & t[36];
  assign t[210] = t[237] ^ x[39];
  assign t[211] = t[238] ^ x[42];
  assign t[212] = t[239] ^ x[45];
  assign t[213] = t[240] ^ x[50];
  assign t[214] = t[241] ^ x[53];
  assign t[215] = t[242] ^ x[58];
  assign t[216] = t[243] ^ x[61];
  assign t[217] = t[244] ^ x[64];
  assign t[218] = t[245] ^ x[67];
  assign t[219] = t[246] ^ x[70];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[81];
  assign t[221] = t[248] ^ x[84];
  assign t[222] = t[249] ^ x[89];
  assign t[223] = t[250] ^ x[92];
  assign t[224] = t[251] ^ x[97];
  assign t[225] = t[252] ^ x[104];
  assign t[226] = (t[253] & ~t[254]);
  assign t[227] = (t[255] & ~t[256]);
  assign t[228] = (t[257] & ~t[258]);
  assign t[229] = (t[259] & ~t[260]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[261] & ~t[262]);
  assign t[231] = (t[263] & ~t[264]);
  assign t[232] = (t[265] & ~t[266]);
  assign t[233] = (t[267] & ~t[268]);
  assign t[234] = (t[269] & ~t[270]);
  assign t[235] = (t[271] & ~t[272]);
  assign t[236] = (t[273] & ~t[274]);
  assign t[237] = (t[275] & ~t[276]);
  assign t[238] = (t[277] & ~t[278]);
  assign t[239] = (t[279] & ~t[280]);
  assign t[23] = ~(t[41] ^ t[42]);
  assign t[240] = (t[281] & ~t[282]);
  assign t[241] = (t[283] & ~t[284]);
  assign t[242] = (t[285] & ~t[286]);
  assign t[243] = (t[287] & ~t[288]);
  assign t[244] = (t[289] & ~t[290]);
  assign t[245] = (t[291] & ~t[292]);
  assign t[246] = (t[293] & ~t[294]);
  assign t[247] = (t[295] & ~t[296]);
  assign t[248] = (t[297] & ~t[298]);
  assign t[249] = (t[299] & ~t[300]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (t[301] & ~t[302]);
  assign t[251] = (t[303] & ~t[304]);
  assign t[252] = (t[305] & ~t[306]);
  assign t[253] = t[307] ^ x[4];
  assign t[254] = t[308] ^ x[3];
  assign t[255] = t[309] ^ x[9];
  assign t[256] = t[310] ^ x[8];
  assign t[257] = t[311] ^ x[12];
  assign t[258] = t[312] ^ x[11];
  assign t[259] = t[313] ^ x[15];
  assign t[25] = t[8] ? t[45] : t[173];
  assign t[260] = t[314] ^ x[14];
  assign t[261] = t[315] ^ x[18];
  assign t[262] = t[316] ^ x[17];
  assign t[263] = t[317] ^ x[21];
  assign t[264] = t[318] ^ x[20];
  assign t[265] = t[319] ^ x[24];
  assign t[266] = t[320] ^ x[23];
  assign t[267] = t[321] ^ x[27];
  assign t[268] = t[322] ^ x[26];
  assign t[269] = t[323] ^ x[30];
  assign t[26] = t[46] ^ t[47];
  assign t[270] = t[324] ^ x[29];
  assign t[271] = t[325] ^ x[33];
  assign t[272] = t[326] ^ x[32];
  assign t[273] = t[327] ^ x[36];
  assign t[274] = t[328] ^ x[35];
  assign t[275] = t[329] ^ x[39];
  assign t[276] = t[330] ^ x[38];
  assign t[277] = t[331] ^ x[42];
  assign t[278] = t[332] ^ x[41];
  assign t[279] = t[333] ^ x[45];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[44];
  assign t[281] = t[335] ^ x[50];
  assign t[282] = t[336] ^ x[49];
  assign t[283] = t[337] ^ x[53];
  assign t[284] = t[338] ^ x[52];
  assign t[285] = t[339] ^ x[58];
  assign t[286] = t[340] ^ x[57];
  assign t[287] = t[341] ^ x[61];
  assign t[288] = t[342] ^ x[60];
  assign t[289] = t[343] ^ x[64];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[63];
  assign t[291] = t[345] ^ x[67];
  assign t[292] = t[346] ^ x[66];
  assign t[293] = t[347] ^ x[70];
  assign t[294] = t[348] ^ x[69];
  assign t[295] = t[349] ^ x[81];
  assign t[296] = t[350] ^ x[80];
  assign t[297] = t[351] ^ x[84];
  assign t[298] = t[352] ^ x[83];
  assign t[299] = t[353] ^ x[89];
  assign t[29] = ~(t[174]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[88];
  assign t[301] = t[355] ^ x[92];
  assign t[302] = t[356] ^ x[91];
  assign t[303] = t[357] ^ x[97];
  assign t[304] = t[358] ^ x[96];
  assign t[305] = t[359] ^ x[104];
  assign t[306] = t[360] ^ x[103];
  assign t[307] = (x[2]);
  assign t[308] = (x[2]);
  assign t[309] = (x[7]);
  assign t[30] = ~(t[175]);
  assign t[310] = (x[7]);
  assign t[311] = (x[10]);
  assign t[312] = (x[10]);
  assign t[313] = (x[13]);
  assign t[314] = (x[13]);
  assign t[315] = (x[16]);
  assign t[316] = (x[16]);
  assign t[317] = (x[19]);
  assign t[318] = (x[19]);
  assign t[319] = (x[22]);
  assign t[31] = ~(t[176]);
  assign t[320] = (x[22]);
  assign t[321] = (x[25]);
  assign t[322] = (x[25]);
  assign t[323] = (x[28]);
  assign t[324] = (x[28]);
  assign t[325] = (x[31]);
  assign t[326] = (x[31]);
  assign t[327] = (x[34]);
  assign t[328] = (x[34]);
  assign t[329] = (x[37]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[37]);
  assign t[331] = (x[40]);
  assign t[332] = (x[40]);
  assign t[333] = (x[43]);
  assign t[334] = (x[43]);
  assign t[335] = (x[48]);
  assign t[336] = (x[48]);
  assign t[337] = (x[51]);
  assign t[338] = (x[51]);
  assign t[339] = (x[56]);
  assign t[33] = t[8] ? t[52] : t[177];
  assign t[340] = (x[56]);
  assign t[341] = (x[59]);
  assign t[342] = (x[59]);
  assign t[343] = (x[62]);
  assign t[344] = (x[62]);
  assign t[345] = (x[65]);
  assign t[346] = (x[65]);
  assign t[347] = (x[68]);
  assign t[348] = (x[68]);
  assign t[349] = (x[79]);
  assign t[34] = t[178] ^ t[53];
  assign t[350] = (x[79]);
  assign t[351] = (x[82]);
  assign t[352] = (x[82]);
  assign t[353] = (x[87]);
  assign t[354] = (x[87]);
  assign t[355] = (x[90]);
  assign t[356] = (x[90]);
  assign t[357] = (x[95]);
  assign t[358] = (x[95]);
  assign t[359] = (x[102]);
  assign t[35] = ~(t[54]);
  assign t[360] = (x[102]);
  assign t[36] = t[175] ^ t[55];
  assign t[37] = t[56];
  assign t[38] = ~t[57];
  assign t[39] = t[58] ^ t[59];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[60] & t[61];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] ^ t[25];
  assign t[44] = t[46] ^ t[67];
  assign t[45] = t[173] ^ t[68];
  assign t[46] = t[69] ^ t[70];
  assign t[47] = t[71] & t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[179] | t[75];
  assign t[4] = t[8] ? t[9] : t[172];
  assign t[50] = ~(t[180]);
  assign t[51] = ~(t[76] & t[178]);
  assign t[52] = t[177] ^ t[77];
  assign t[53] = t[8] ? t[78] : t[181];
  assign t[54] = t[174] ^ t[79];
  assign t[55] = t[8] ? t[80] : t[182];
  assign t[56] = t[27] ? t[81] : t[183];
  assign t[57] = t[27] ? t[82] : t[184];
  assign t[58] = t[83] & t[84];
  assign t[59] = t[85] & t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = ~(t[58] ^ t[87]);
  assign t[61] = t[88] ^ t[89];
  assign t[62] = t[90] ^ t[91];
  assign t[63] = t[38] ^ t[92];
  assign t[64] = t[93] ^ t[94];
  assign t[65] = t[95] & t[96];
  assign t[66] = t[8] ? t[97] : t[185];
  assign t[67] = t[98] & t[99];
  assign t[68] = t[100] ? x[47] : x[46];
  assign t[69] = t[101] & t[102];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[103] & t[104];
  assign t[71] = ~(t[105] ^ t[46]);
  assign t[72] = t[43] ^ t[104];
  assign t[73] = ~(t[75] & t[106]);
  assign t[74] = ~(t[186] ^ t[107]);
  assign t[75] = ~(t[108] & t[109]);
  assign t[76] = ~(t[187]);
  assign t[77] = t[28] ? x[55] : x[54];
  assign t[78] = t[181] ^ t[110];
  assign t[79] = t[27] ? t[111] : t[188];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[182] ^ t[112];
  assign t[81] = t[183] ^ t[113];
  assign t[82] = t[184] ^ t[114];
  assign t[83] = ~(t[89]);
  assign t[84] = ~(t[115]);
  assign t[85] = ~(t[37]);
  assign t[86] = t[116];
  assign t[87] = t[21] ^ t[115];
  assign t[88] = t[115] ^ t[38];
  assign t[89] = t[86] ^ t[37];
  assign t[8] = ~(t[15]);
  assign t[90] = t[54] ^ t[34];
  assign t[91] = t[117] ^ t[118];
  assign t[92] = t[39] ^ t[119];
  assign t[93] = t[120] ? t[121] : t[189];
  assign t[94] = t[120] ? t[122] : t[190];
  assign t[95] = ~(t[64] ^ t[123]);
  assign t[96] = t[124] ^ t[125];
  assign t[97] = t[185] ^ t[126];
  assign t[98] = ~(t[69] ^ t[127]);
  assign t[99] = t[128] ^ t[129];
  assign t[9] = t[172] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind81(x, y);
 input [116:0] x;
 output y;

 wire [360:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[130]);
  assign t[101] = ~(t[129]);
  assign t[102] = ~(t[131]);
  assign t[103] = ~(t[66]);
  assign t[104] = t[8] ? t[132] : t[191];
  assign t[105] = t[131] ^ t[66];
  assign t[106] = ~(t[133] & t[134]);
  assign t[107] = t[135] ^ t[192];
  assign t[108] = ~(t[186]);
  assign t[109] = t[136] & t[135];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[28] ? x[72] : x[71];
  assign t[111] = t[188] ^ t[137];
  assign t[112] = t[138] ? x[74] : x[73];
  assign t[113] = t[138] ? x[76] : x[75];
  assign t[114] = t[28] ? x[78] : x[77];
  assign t[115] = ~t[139];
  assign t[116] = t[27] ? t[140] : t[193];
  assign t[117] = t[141] ^ t[20];
  assign t[118] = t[142] & t[143];
  assign t[119] = t[144] & t[145];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = ~(t[15]);
  assign t[121] = t[189] ^ t[146];
  assign t[122] = t[190] ^ t[147];
  assign t[123] = t[148] ^ t[149];
  assign t[124] = t[94] ^ t[150];
  assign t[125] = t[120] ? t[151] : t[194];
  assign t[126] = t[100] ? x[86] : x[85];
  assign t[127] = t[43] ^ t[131];
  assign t[128] = t[131] ^ t[25];
  assign t[129] = t[104] ^ t[66];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = ~(t[28]);
  assign t[131] = t[8] ? t[152] : t[195];
  assign t[132] = t[191] ^ t[153];
  assign t[133] = ~(t[136] | t[135]);
  assign t[134] = ~(t[154] | t[108]);
  assign t[135] = ~(t[196]);
  assign t[136] = ~(t[192]);
  assign t[137] = t[138] ? x[94] : x[93];
  assign t[138] = ~(t[130]);
  assign t[139] = t[27] ? t[155] : t[197];
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[193] ^ t[156];
  assign t[141] = t[157] & t[158];
  assign t[142] = ~(t[141] ^ t[159]);
  assign t[143] = t[19] ^ t[160];
  assign t[144] = ~(t[161] ^ t[39]);
  assign t[145] = t[21] ^ t[86];
  assign t[146] = t[162] ? x[99] : x[98];
  assign t[147] = t[162] ? x[101] : x[100];
  assign t[148] = t[163] & t[164];
  assign t[149] = t[165] & t[125];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[120] ? t[166] : t[198];
  assign t[151] = t[194] ^ t[167];
  assign t[152] = t[195] ^ t[168];
  assign t[153] = t[100] ? x[106] : x[105];
  assign t[154] = ~(t[179]);
  assign t[155] = t[197] ^ t[169];
  assign t[156] = t[100] ? x[108] : x[107];
  assign t[157] = ~(t[160]);
  assign t[158] = ~(t[33]);
  assign t[159] = t[90] ^ t[33];
  assign t[15] = ~(t[27]);
  assign t[160] = t[36] ^ t[54];
  assign t[161] = t[115] ^ t[37];
  assign t[162] = ~(t[130]);
  assign t[163] = ~(t[170]);
  assign t[164] = ~(t[93]);
  assign t[165] = ~(t[94]);
  assign t[166] = t[198] ^ t[171];
  assign t[167] = t[162] ? x[110] : x[109];
  assign t[168] = t[100] ? x[112] : x[111];
  assign t[169] = t[28] ? x[114] : x[113];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[125] ^ t[94];
  assign t[171] = t[162] ? x[116] : x[115];
  assign t[172] = (t[199]);
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = t[226] ^ x[4];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[9];
  assign t[201] = t[228] ^ x[12];
  assign t[202] = t[229] ^ x[15];
  assign t[203] = t[230] ^ x[18];
  assign t[204] = t[231] ^ x[21];
  assign t[205] = t[232] ^ x[24];
  assign t[206] = t[233] ^ x[27];
  assign t[207] = t[234] ^ x[30];
  assign t[208] = t[235] ^ x[33];
  assign t[209] = t[236] ^ x[36];
  assign t[20] = t[35] & t[36];
  assign t[210] = t[237] ^ x[39];
  assign t[211] = t[238] ^ x[42];
  assign t[212] = t[239] ^ x[45];
  assign t[213] = t[240] ^ x[50];
  assign t[214] = t[241] ^ x[53];
  assign t[215] = t[242] ^ x[58];
  assign t[216] = t[243] ^ x[61];
  assign t[217] = t[244] ^ x[64];
  assign t[218] = t[245] ^ x[67];
  assign t[219] = t[246] ^ x[70];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[81];
  assign t[221] = t[248] ^ x[84];
  assign t[222] = t[249] ^ x[89];
  assign t[223] = t[250] ^ x[92];
  assign t[224] = t[251] ^ x[97];
  assign t[225] = t[252] ^ x[104];
  assign t[226] = (t[253] & ~t[254]);
  assign t[227] = (t[255] & ~t[256]);
  assign t[228] = (t[257] & ~t[258]);
  assign t[229] = (t[259] & ~t[260]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[261] & ~t[262]);
  assign t[231] = (t[263] & ~t[264]);
  assign t[232] = (t[265] & ~t[266]);
  assign t[233] = (t[267] & ~t[268]);
  assign t[234] = (t[269] & ~t[270]);
  assign t[235] = (t[271] & ~t[272]);
  assign t[236] = (t[273] & ~t[274]);
  assign t[237] = (t[275] & ~t[276]);
  assign t[238] = (t[277] & ~t[278]);
  assign t[239] = (t[279] & ~t[280]);
  assign t[23] = ~(t[41] ^ t[42]);
  assign t[240] = (t[281] & ~t[282]);
  assign t[241] = (t[283] & ~t[284]);
  assign t[242] = (t[285] & ~t[286]);
  assign t[243] = (t[287] & ~t[288]);
  assign t[244] = (t[289] & ~t[290]);
  assign t[245] = (t[291] & ~t[292]);
  assign t[246] = (t[293] & ~t[294]);
  assign t[247] = (t[295] & ~t[296]);
  assign t[248] = (t[297] & ~t[298]);
  assign t[249] = (t[299] & ~t[300]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (t[301] & ~t[302]);
  assign t[251] = (t[303] & ~t[304]);
  assign t[252] = (t[305] & ~t[306]);
  assign t[253] = t[307] ^ x[4];
  assign t[254] = t[308] ^ x[3];
  assign t[255] = t[309] ^ x[9];
  assign t[256] = t[310] ^ x[8];
  assign t[257] = t[311] ^ x[12];
  assign t[258] = t[312] ^ x[11];
  assign t[259] = t[313] ^ x[15];
  assign t[25] = t[8] ? t[45] : t[173];
  assign t[260] = t[314] ^ x[14];
  assign t[261] = t[315] ^ x[18];
  assign t[262] = t[316] ^ x[17];
  assign t[263] = t[317] ^ x[21];
  assign t[264] = t[318] ^ x[20];
  assign t[265] = t[319] ^ x[24];
  assign t[266] = t[320] ^ x[23];
  assign t[267] = t[321] ^ x[27];
  assign t[268] = t[322] ^ x[26];
  assign t[269] = t[323] ^ x[30];
  assign t[26] = t[46] ^ t[47];
  assign t[270] = t[324] ^ x[29];
  assign t[271] = t[325] ^ x[33];
  assign t[272] = t[326] ^ x[32];
  assign t[273] = t[327] ^ x[36];
  assign t[274] = t[328] ^ x[35];
  assign t[275] = t[329] ^ x[39];
  assign t[276] = t[330] ^ x[38];
  assign t[277] = t[331] ^ x[42];
  assign t[278] = t[332] ^ x[41];
  assign t[279] = t[333] ^ x[45];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[44];
  assign t[281] = t[335] ^ x[50];
  assign t[282] = t[336] ^ x[49];
  assign t[283] = t[337] ^ x[53];
  assign t[284] = t[338] ^ x[52];
  assign t[285] = t[339] ^ x[58];
  assign t[286] = t[340] ^ x[57];
  assign t[287] = t[341] ^ x[61];
  assign t[288] = t[342] ^ x[60];
  assign t[289] = t[343] ^ x[64];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[63];
  assign t[291] = t[345] ^ x[67];
  assign t[292] = t[346] ^ x[66];
  assign t[293] = t[347] ^ x[70];
  assign t[294] = t[348] ^ x[69];
  assign t[295] = t[349] ^ x[81];
  assign t[296] = t[350] ^ x[80];
  assign t[297] = t[351] ^ x[84];
  assign t[298] = t[352] ^ x[83];
  assign t[299] = t[353] ^ x[89];
  assign t[29] = ~(t[174]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[88];
  assign t[301] = t[355] ^ x[92];
  assign t[302] = t[356] ^ x[91];
  assign t[303] = t[357] ^ x[97];
  assign t[304] = t[358] ^ x[96];
  assign t[305] = t[359] ^ x[104];
  assign t[306] = t[360] ^ x[103];
  assign t[307] = (x[2]);
  assign t[308] = (x[2]);
  assign t[309] = (x[7]);
  assign t[30] = ~(t[175]);
  assign t[310] = (x[7]);
  assign t[311] = (x[10]);
  assign t[312] = (x[10]);
  assign t[313] = (x[13]);
  assign t[314] = (x[13]);
  assign t[315] = (x[16]);
  assign t[316] = (x[16]);
  assign t[317] = (x[19]);
  assign t[318] = (x[19]);
  assign t[319] = (x[22]);
  assign t[31] = ~(t[176]);
  assign t[320] = (x[22]);
  assign t[321] = (x[25]);
  assign t[322] = (x[25]);
  assign t[323] = (x[28]);
  assign t[324] = (x[28]);
  assign t[325] = (x[31]);
  assign t[326] = (x[31]);
  assign t[327] = (x[34]);
  assign t[328] = (x[34]);
  assign t[329] = (x[37]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[37]);
  assign t[331] = (x[40]);
  assign t[332] = (x[40]);
  assign t[333] = (x[43]);
  assign t[334] = (x[43]);
  assign t[335] = (x[48]);
  assign t[336] = (x[48]);
  assign t[337] = (x[51]);
  assign t[338] = (x[51]);
  assign t[339] = (x[56]);
  assign t[33] = t[8] ? t[52] : t[177];
  assign t[340] = (x[56]);
  assign t[341] = (x[59]);
  assign t[342] = (x[59]);
  assign t[343] = (x[62]);
  assign t[344] = (x[62]);
  assign t[345] = (x[65]);
  assign t[346] = (x[65]);
  assign t[347] = (x[68]);
  assign t[348] = (x[68]);
  assign t[349] = (x[79]);
  assign t[34] = t[178] ^ t[53];
  assign t[350] = (x[79]);
  assign t[351] = (x[82]);
  assign t[352] = (x[82]);
  assign t[353] = (x[87]);
  assign t[354] = (x[87]);
  assign t[355] = (x[90]);
  assign t[356] = (x[90]);
  assign t[357] = (x[95]);
  assign t[358] = (x[95]);
  assign t[359] = (x[102]);
  assign t[35] = ~(t[54]);
  assign t[360] = (x[102]);
  assign t[36] = t[175] ^ t[55];
  assign t[37] = t[56];
  assign t[38] = ~t[57];
  assign t[39] = t[58] ^ t[59];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[60] & t[61];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] ^ t[25];
  assign t[44] = t[46] ^ t[67];
  assign t[45] = t[173] ^ t[68];
  assign t[46] = t[69] ^ t[70];
  assign t[47] = t[71] & t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[179] | t[75];
  assign t[4] = t[8] ? t[9] : t[172];
  assign t[50] = ~(t[180]);
  assign t[51] = ~(t[76] & t[178]);
  assign t[52] = t[177] ^ t[77];
  assign t[53] = t[8] ? t[78] : t[181];
  assign t[54] = t[174] ^ t[79];
  assign t[55] = t[8] ? t[80] : t[182];
  assign t[56] = t[27] ? t[81] : t[183];
  assign t[57] = t[27] ? t[82] : t[184];
  assign t[58] = t[83] & t[84];
  assign t[59] = t[85] & t[86];
  assign t[5] = ~(t[10]);
  assign t[60] = ~(t[58] ^ t[87]);
  assign t[61] = t[88] ^ t[89];
  assign t[62] = t[90] ^ t[91];
  assign t[63] = t[38] ^ t[92];
  assign t[64] = t[93] ^ t[94];
  assign t[65] = t[95] & t[96];
  assign t[66] = t[8] ? t[97] : t[185];
  assign t[67] = t[98] & t[99];
  assign t[68] = t[100] ? x[47] : x[46];
  assign t[69] = t[101] & t[102];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[103] & t[104];
  assign t[71] = ~(t[105] ^ t[46]);
  assign t[72] = t[43] ^ t[104];
  assign t[73] = ~(t[75] & t[106]);
  assign t[74] = ~(t[186] ^ t[107]);
  assign t[75] = ~(t[108] & t[109]);
  assign t[76] = ~(t[187]);
  assign t[77] = t[28] ? x[55] : x[54];
  assign t[78] = t[181] ^ t[110];
  assign t[79] = t[27] ? t[111] : t[188];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[182] ^ t[112];
  assign t[81] = t[183] ^ t[113];
  assign t[82] = t[184] ^ t[114];
  assign t[83] = ~(t[89]);
  assign t[84] = ~(t[115]);
  assign t[85] = ~(t[37]);
  assign t[86] = t[116];
  assign t[87] = t[21] ^ t[115];
  assign t[88] = t[115] ^ t[38];
  assign t[89] = t[86] ^ t[37];
  assign t[8] = ~(t[15]);
  assign t[90] = t[54] ^ t[34];
  assign t[91] = t[117] ^ t[118];
  assign t[92] = t[39] ^ t[119];
  assign t[93] = t[120] ? t[121] : t[189];
  assign t[94] = t[120] ? t[122] : t[190];
  assign t[95] = ~(t[64] ^ t[123]);
  assign t[96] = t[124] ^ t[125];
  assign t[97] = t[185] ^ t[126];
  assign t[98] = ~(t[69] ^ t[127]);
  assign t[99] = t[128] ^ t[129];
  assign t[9] = t[172] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [116:0] x;
 output y;

 wire [381:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[127] ^ t[132];
  assign t[101] = t[133] ^ t[134];
  assign t[102] = t[135] ^ t[39];
  assign t[103] = t[202] ^ t[136];
  assign t[104] = t[122] ^ t[65];
  assign t[105] = ~(t[137] & t[138]);
  assign t[106] = t[139] ^ t[208];
  assign t[107] = ~(t[205]);
  assign t[108] = t[140] & t[139];
  assign t[109] = t[38] ^ t[57];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[78] ? x[59] : x[58];
  assign t[111] = t[76] ? x[61] : x[60];
  assign t[112] = ~(t[141]);
  assign t[113] = ~(t[135]);
  assign t[114] = ~(t[90]);
  assign t[115] = t[142];
  assign t[116] = t[135] ^ t[90];
  assign t[117] = t[27] ? t[143] : t[209];
  assign t[118] = ~(t[86] ^ t[144]);
  assign t[119] = t[102] ^ t[141];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[207] ^ t[145];
  assign t[121] = t[27] ? t[146] : t[210];
  assign t[122] = t[147] ^ t[148];
  assign t[123] = t[93] ^ t[103];
  assign t[124] = t[196] ^ t[149];
  assign t[125] = t[122] ^ t[150];
  assign t[126] = t[151] ? t[152] : t[211];
  assign t[127] = t[151] ? t[153] : t[212];
  assign t[128] = ~(t[97] ^ t[133]);
  assign t[129] = t[100] ^ t[154];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = ~(t[53] ^ t[155]);
  assign t[131] = t[21] ^ t[109];
  assign t[132] = t[151] ? t[156] : t[213];
  assign t[133] = t[157] ^ t[158];
  assign t[134] = t[159] & t[160];
  assign t[135] = ~t[161];
  assign t[136] = t[8] ? t[162] : t[214];
  assign t[137] = ~(t[140] | t[139]);
  assign t[138] = ~(t[163] | t[107]);
  assign t[139] = ~(t[215]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = ~(t[208]);
  assign t[141] = t[115] ^ t[90];
  assign t[142] = t[27] ? t[164] : t[216];
  assign t[143] = t[209] ^ t[165];
  assign t[144] = t[62] ^ t[135];
  assign t[145] = t[76] ? x[87] : x[86];
  assign t[146] = t[210] ^ t[166];
  assign t[147] = t[167] & t[168];
  assign t[148] = t[169] & t[124];
  assign t[149] = t[8] ? t[170] : t[217];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[171] & t[172];
  assign t[151] = ~(t[15]);
  assign t[152] = t[211] ^ t[173];
  assign t[153] = t[212] ^ t[174];
  assign t[154] = t[151] ? t[175] : t[218];
  assign t[155] = t[68] ^ t[36];
  assign t[156] = t[213] ^ t[176];
  assign t[157] = t[177] & t[178];
  assign t[158] = t[179] & t[154];
  assign t[159] = ~(t[157] ^ t[180]);
  assign t[15] = ~(t[27]);
  assign t[160] = t[181] ^ t[182];
  assign t[161] = t[27] ? t[183] : t[219];
  assign t[162] = t[214] ^ t[184];
  assign t[163] = ~(t[200]);
  assign t[164] = t[216] ^ t[185];
  assign t[165] = t[28] ? x[98] : x[97];
  assign t[166] = t[28] ? x[100] : x[99];
  assign t[167] = ~(t[186]);
  assign t[168] = ~(t[92]);
  assign t[169] = ~(t[93]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[217] ^ t[187];
  assign t[171] = ~(t[147] ^ t[188]);
  assign t[172] = t[189] ^ t[186];
  assign t[173] = t[190] ? x[102] : x[101];
  assign t[174] = t[190] ? x[104] : x[103];
  assign t[175] = t[218] ^ t[191];
  assign t[176] = t[190] ? x[106] : x[105];
  assign t[177] = ~(t[182]);
  assign t[178] = ~(t[126]);
  assign t[179] = ~(t[127]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[100] ^ t[126];
  assign t[181] = t[126] ^ t[132];
  assign t[182] = t[154] ^ t[127];
  assign t[183] = t[219] ^ t[192];
  assign t[184] = t[76] ? x[108] : x[107];
  assign t[185] = t[78] ? x[110] : x[109];
  assign t[186] = t[124] ^ t[93];
  assign t[187] = t[28] ? x[112] : x[111];
  assign t[188] = t[123] ^ t[92];
  assign t[189] = t[92] ^ t[103];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = ~(t[49]);
  assign t[191] = t[190] ? x[114] : x[113];
  assign t[192] = t[76] ? x[116] : x[115];
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[8] ? t[33] : t[194];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[34] ^ t[35];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[36] ^ t[19];
  assign t[220] = t[247] ^ x[4];
  assign t[221] = t[248] ^ x[9];
  assign t[222] = t[249] ^ x[12];
  assign t[223] = t[250] ^ x[15];
  assign t[224] = t[251] ^ x[18];
  assign t[225] = t[252] ^ x[21];
  assign t[226] = t[253] ^ x[24];
  assign t[227] = t[254] ^ x[27];
  assign t[228] = t[255] ^ x[30];
  assign t[229] = t[256] ^ x[33];
  assign t[22] = t[37] & t[38];
  assign t[230] = t[257] ^ x[38];
  assign t[231] = t[258] ^ x[41];
  assign t[232] = t[259] ^ x[44];
  assign t[233] = t[260] ^ x[47];
  assign t[234] = t[261] ^ x[54];
  assign t[235] = t[262] ^ x[57];
  assign t[236] = t[263] ^ x[64];
  assign t[237] = t[264] ^ x[67];
  assign t[238] = t[265] ^ x[70];
  assign t[239] = t[266] ^ x[73];
  assign t[23] = t[39] ^ t[40];
  assign t[240] = t[267] ^ x[76];
  assign t[241] = t[268] ^ x[79];
  assign t[242] = t[269] ^ x[82];
  assign t[243] = t[270] ^ x[85];
  assign t[244] = t[271] ^ x[90];
  assign t[245] = t[272] ^ x[93];
  assign t[246] = t[273] ^ x[96];
  assign t[247] = (t[274] & ~t[275]);
  assign t[248] = (t[276] & ~t[277]);
  assign t[249] = (t[278] & ~t[279]);
  assign t[24] = t[41] ^ t[42];
  assign t[250] = (t[280] & ~t[281]);
  assign t[251] = (t[282] & ~t[283]);
  assign t[252] = (t[284] & ~t[285]);
  assign t[253] = (t[286] & ~t[287]);
  assign t[254] = (t[288] & ~t[289]);
  assign t[255] = (t[290] & ~t[291]);
  assign t[256] = (t[292] & ~t[293]);
  assign t[257] = (t[294] & ~t[295]);
  assign t[258] = (t[296] & ~t[297]);
  assign t[259] = (t[298] & ~t[299]);
  assign t[25] = ~(t[43] ^ t[44]);
  assign t[260] = (t[300] & ~t[301]);
  assign t[261] = (t[302] & ~t[303]);
  assign t[262] = (t[304] & ~t[305]);
  assign t[263] = (t[306] & ~t[307]);
  assign t[264] = (t[308] & ~t[309]);
  assign t[265] = (t[310] & ~t[311]);
  assign t[266] = (t[312] & ~t[313]);
  assign t[267] = (t[314] & ~t[315]);
  assign t[268] = (t[316] & ~t[317]);
  assign t[269] = (t[318] & ~t[319]);
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[270] = (t[320] & ~t[321]);
  assign t[271] = (t[322] & ~t[323]);
  assign t[272] = (t[324] & ~t[325]);
  assign t[273] = (t[326] & ~t[327]);
  assign t[274] = t[328] ^ x[4];
  assign t[275] = t[329] ^ x[3];
  assign t[276] = t[330] ^ x[9];
  assign t[277] = t[331] ^ x[8];
  assign t[278] = t[332] ^ x[12];
  assign t[279] = t[333] ^ x[11];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[334] ^ x[15];
  assign t[281] = t[335] ^ x[14];
  assign t[282] = t[336] ^ x[18];
  assign t[283] = t[337] ^ x[17];
  assign t[284] = t[338] ^ x[21];
  assign t[285] = t[339] ^ x[20];
  assign t[286] = t[340] ^ x[24];
  assign t[287] = t[341] ^ x[23];
  assign t[288] = t[342] ^ x[27];
  assign t[289] = t[343] ^ x[26];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[30];
  assign t[291] = t[345] ^ x[29];
  assign t[292] = t[346] ^ x[33];
  assign t[293] = t[347] ^ x[32];
  assign t[294] = t[348] ^ x[38];
  assign t[295] = t[349] ^ x[37];
  assign t[296] = t[350] ^ x[41];
  assign t[297] = t[351] ^ x[40];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[43];
  assign t[29] = ~(t[195]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[47];
  assign t[301] = t[355] ^ x[46];
  assign t[302] = t[356] ^ x[54];
  assign t[303] = t[357] ^ x[53];
  assign t[304] = t[358] ^ x[57];
  assign t[305] = t[359] ^ x[56];
  assign t[306] = t[360] ^ x[64];
  assign t[307] = t[361] ^ x[63];
  assign t[308] = t[362] ^ x[67];
  assign t[309] = t[363] ^ x[66];
  assign t[30] = ~(t[196]);
  assign t[310] = t[364] ^ x[70];
  assign t[311] = t[365] ^ x[69];
  assign t[312] = t[366] ^ x[73];
  assign t[313] = t[367] ^ x[72];
  assign t[314] = t[368] ^ x[76];
  assign t[315] = t[369] ^ x[75];
  assign t[316] = t[370] ^ x[79];
  assign t[317] = t[371] ^ x[78];
  assign t[318] = t[372] ^ x[82];
  assign t[319] = t[373] ^ x[81];
  assign t[31] = ~(t[197]);
  assign t[320] = t[374] ^ x[85];
  assign t[321] = t[375] ^ x[84];
  assign t[322] = t[376] ^ x[90];
  assign t[323] = t[377] ^ x[89];
  assign t[324] = t[378] ^ x[93];
  assign t[325] = t[379] ^ x[92];
  assign t[326] = t[380] ^ x[96];
  assign t[327] = t[381] ^ x[95];
  assign t[328] = (x[2]);
  assign t[329] = (x[2]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[7]);
  assign t[331] = (x[7]);
  assign t[332] = (x[10]);
  assign t[333] = (x[10]);
  assign t[334] = (x[13]);
  assign t[335] = (x[13]);
  assign t[336] = (x[16]);
  assign t[337] = (x[16]);
  assign t[338] = (x[19]);
  assign t[339] = (x[19]);
  assign t[33] = t[194] ^ t[52];
  assign t[340] = (x[22]);
  assign t[341] = (x[22]);
  assign t[342] = (x[25]);
  assign t[343] = (x[25]);
  assign t[344] = (x[28]);
  assign t[345] = (x[28]);
  assign t[346] = (x[31]);
  assign t[347] = (x[31]);
  assign t[348] = (x[36]);
  assign t[349] = (x[36]);
  assign t[34] = t[53] ^ t[22];
  assign t[350] = (x[39]);
  assign t[351] = (x[39]);
  assign t[352] = (x[42]);
  assign t[353] = (x[42]);
  assign t[354] = (x[45]);
  assign t[355] = (x[45]);
  assign t[356] = (x[52]);
  assign t[357] = (x[52]);
  assign t[358] = (x[55]);
  assign t[359] = (x[55]);
  assign t[35] = t[54] & t[55];
  assign t[360] = (x[62]);
  assign t[361] = (x[62]);
  assign t[362] = (x[65]);
  assign t[363] = (x[65]);
  assign t[364] = (x[68]);
  assign t[365] = (x[68]);
  assign t[366] = (x[71]);
  assign t[367] = (x[71]);
  assign t[368] = (x[74]);
  assign t[369] = (x[74]);
  assign t[36] = t[8] ? t[56] : t[198];
  assign t[370] = (x[77]);
  assign t[371] = (x[77]);
  assign t[372] = (x[80]);
  assign t[373] = (x[80]);
  assign t[374] = (x[83]);
  assign t[375] = (x[83]);
  assign t[376] = (x[88]);
  assign t[377] = (x[88]);
  assign t[378] = (x[91]);
  assign t[379] = (x[91]);
  assign t[37] = ~(t[57]);
  assign t[380] = (x[94]);
  assign t[381] = (x[94]);
  assign t[38] = t[8] ? t[58] : t[199];
  assign t[39] = ~t[59];
  assign t[3] = t[6] ^ t[7];
  assign t[40] = t[60] ^ t[61];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[66] ^ t[67]);
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[11] ^ t[72]);
  assign t[47] = ~(t[73] & t[74]);
  assign t[48] = t[200] | t[75];
  assign t[49] = ~(t[76]);
  assign t[4] = t[8] ? t[9] : t[193];
  assign t[50] = ~(t[201]);
  assign t[51] = ~(t[77] & t[202]);
  assign t[52] = t[78] ? x[35] : x[34];
  assign t[53] = t[79] & t[80];
  assign t[54] = ~(t[81] ^ t[34]);
  assign t[55] = t[68] ^ t[38];
  assign t[56] = t[198] ^ t[82];
  assign t[57] = t[8] ? t[83] : t[203];
  assign t[58] = t[199] ^ t[84];
  assign t[59] = t[27] ? t[85] : t[204];
  assign t[5] = ~(t[10]);
  assign t[60] = t[86] ^ t[87];
  assign t[61] = t[88] & t[89];
  assign t[62] = t[90] ^ t[39];
  assign t[63] = t[60] ^ t[91];
  assign t[64] = t[92] ^ t[93];
  assign t[65] = t[94] & t[95];
  assign t[66] = t[96] ^ t[23];
  assign t[67] = t[97] ^ t[98];
  assign t[68] = t[57] ^ t[19];
  assign t[69] = t[34] ^ t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[100] ^ t[101];
  assign t[71] = t[102] ^ t[87];
  assign t[72] = t[103] ^ t[104];
  assign t[73] = ~(t[75] & t[105]);
  assign t[74] = ~(t[205] ^ t[106]);
  assign t[75] = ~(t[107] & t[108]);
  assign t[76] = ~(t[48]);
  assign t[77] = ~(t[206]);
  assign t[78] = ~(t[49]);
  assign t[79] = ~(t[109]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[36]);
  assign t[81] = t[36] ^ t[57];
  assign t[82] = t[78] ? x[49] : x[48];
  assign t[83] = t[203] ^ t[110];
  assign t[84] = t[78] ? x[51] : x[50];
  assign t[85] = t[204] ^ t[111];
  assign t[86] = t[112] & t[113];
  assign t[87] = t[114] & t[115];
  assign t[88] = ~(t[116] ^ t[60]);
  assign t[89] = t[62] ^ t[115];
  assign t[8] = ~(t[15]);
  assign t[90] = t[117];
  assign t[91] = t[118] & t[119];
  assign t[92] = t[8] ? t[120] : t[207];
  assign t[93] = t[195] ^ t[121];
  assign t[94] = ~(t[64] ^ t[122]);
  assign t[95] = t[123] ^ t[124];
  assign t[96] = t[123] ^ t[125];
  assign t[97] = t[126] ^ t[127];
  assign t[98] = t[128] & t[129];
  assign t[99] = t[130] & t[131];
  assign t[9] = t[193] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [116:0] x;
 output y;

 wire [381:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[127] ^ t[132];
  assign t[101] = t[133] ^ t[134];
  assign t[102] = t[135] ^ t[39];
  assign t[103] = t[202] ^ t[136];
  assign t[104] = t[122] ^ t[65];
  assign t[105] = ~(t[137] & t[138]);
  assign t[106] = t[139] ^ t[208];
  assign t[107] = ~(t[205]);
  assign t[108] = t[140] & t[139];
  assign t[109] = t[38] ^ t[57];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[78] ? x[59] : x[58];
  assign t[111] = t[76] ? x[61] : x[60];
  assign t[112] = ~(t[141]);
  assign t[113] = ~(t[135]);
  assign t[114] = ~(t[90]);
  assign t[115] = t[142];
  assign t[116] = t[135] ^ t[90];
  assign t[117] = t[27] ? t[143] : t[209];
  assign t[118] = ~(t[86] ^ t[144]);
  assign t[119] = t[102] ^ t[141];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[207] ^ t[145];
  assign t[121] = t[27] ? t[146] : t[210];
  assign t[122] = t[147] ^ t[148];
  assign t[123] = t[93] ^ t[103];
  assign t[124] = t[196] ^ t[149];
  assign t[125] = t[122] ^ t[150];
  assign t[126] = t[151] ? t[152] : t[211];
  assign t[127] = t[151] ? t[153] : t[212];
  assign t[128] = ~(t[97] ^ t[133]);
  assign t[129] = t[100] ^ t[154];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = ~(t[53] ^ t[155]);
  assign t[131] = t[21] ^ t[109];
  assign t[132] = t[151] ? t[156] : t[213];
  assign t[133] = t[157] ^ t[158];
  assign t[134] = t[159] & t[160];
  assign t[135] = ~t[161];
  assign t[136] = t[8] ? t[162] : t[214];
  assign t[137] = ~(t[140] | t[139]);
  assign t[138] = ~(t[163] | t[107]);
  assign t[139] = ~(t[215]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = ~(t[208]);
  assign t[141] = t[115] ^ t[90];
  assign t[142] = t[27] ? t[164] : t[216];
  assign t[143] = t[209] ^ t[165];
  assign t[144] = t[62] ^ t[135];
  assign t[145] = t[76] ? x[87] : x[86];
  assign t[146] = t[210] ^ t[166];
  assign t[147] = t[167] & t[168];
  assign t[148] = t[169] & t[124];
  assign t[149] = t[8] ? t[170] : t[217];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[171] & t[172];
  assign t[151] = ~(t[15]);
  assign t[152] = t[211] ^ t[173];
  assign t[153] = t[212] ^ t[174];
  assign t[154] = t[151] ? t[175] : t[218];
  assign t[155] = t[68] ^ t[36];
  assign t[156] = t[213] ^ t[176];
  assign t[157] = t[177] & t[178];
  assign t[158] = t[179] & t[154];
  assign t[159] = ~(t[157] ^ t[180]);
  assign t[15] = ~(t[27]);
  assign t[160] = t[181] ^ t[182];
  assign t[161] = t[27] ? t[183] : t[219];
  assign t[162] = t[214] ^ t[184];
  assign t[163] = ~(t[200]);
  assign t[164] = t[216] ^ t[185];
  assign t[165] = t[28] ? x[98] : x[97];
  assign t[166] = t[28] ? x[100] : x[99];
  assign t[167] = ~(t[186]);
  assign t[168] = ~(t[92]);
  assign t[169] = ~(t[93]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[217] ^ t[187];
  assign t[171] = ~(t[147] ^ t[188]);
  assign t[172] = t[189] ^ t[186];
  assign t[173] = t[190] ? x[102] : x[101];
  assign t[174] = t[190] ? x[104] : x[103];
  assign t[175] = t[218] ^ t[191];
  assign t[176] = t[190] ? x[106] : x[105];
  assign t[177] = ~(t[182]);
  assign t[178] = ~(t[126]);
  assign t[179] = ~(t[127]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[100] ^ t[126];
  assign t[181] = t[126] ^ t[132];
  assign t[182] = t[154] ^ t[127];
  assign t[183] = t[219] ^ t[192];
  assign t[184] = t[76] ? x[108] : x[107];
  assign t[185] = t[78] ? x[110] : x[109];
  assign t[186] = t[124] ^ t[93];
  assign t[187] = t[28] ? x[112] : x[111];
  assign t[188] = t[123] ^ t[92];
  assign t[189] = t[92] ^ t[103];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = ~(t[49]);
  assign t[191] = t[190] ? x[114] : x[113];
  assign t[192] = t[76] ? x[116] : x[115];
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[8] ? t[33] : t[194];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[34] ^ t[35];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[36] ^ t[19];
  assign t[220] = t[247] ^ x[4];
  assign t[221] = t[248] ^ x[9];
  assign t[222] = t[249] ^ x[12];
  assign t[223] = t[250] ^ x[15];
  assign t[224] = t[251] ^ x[18];
  assign t[225] = t[252] ^ x[21];
  assign t[226] = t[253] ^ x[24];
  assign t[227] = t[254] ^ x[27];
  assign t[228] = t[255] ^ x[30];
  assign t[229] = t[256] ^ x[33];
  assign t[22] = t[37] & t[38];
  assign t[230] = t[257] ^ x[38];
  assign t[231] = t[258] ^ x[41];
  assign t[232] = t[259] ^ x[44];
  assign t[233] = t[260] ^ x[47];
  assign t[234] = t[261] ^ x[54];
  assign t[235] = t[262] ^ x[57];
  assign t[236] = t[263] ^ x[64];
  assign t[237] = t[264] ^ x[67];
  assign t[238] = t[265] ^ x[70];
  assign t[239] = t[266] ^ x[73];
  assign t[23] = t[39] ^ t[40];
  assign t[240] = t[267] ^ x[76];
  assign t[241] = t[268] ^ x[79];
  assign t[242] = t[269] ^ x[82];
  assign t[243] = t[270] ^ x[85];
  assign t[244] = t[271] ^ x[90];
  assign t[245] = t[272] ^ x[93];
  assign t[246] = t[273] ^ x[96];
  assign t[247] = (t[274] & ~t[275]);
  assign t[248] = (t[276] & ~t[277]);
  assign t[249] = (t[278] & ~t[279]);
  assign t[24] = t[41] ^ t[42];
  assign t[250] = (t[280] & ~t[281]);
  assign t[251] = (t[282] & ~t[283]);
  assign t[252] = (t[284] & ~t[285]);
  assign t[253] = (t[286] & ~t[287]);
  assign t[254] = (t[288] & ~t[289]);
  assign t[255] = (t[290] & ~t[291]);
  assign t[256] = (t[292] & ~t[293]);
  assign t[257] = (t[294] & ~t[295]);
  assign t[258] = (t[296] & ~t[297]);
  assign t[259] = (t[298] & ~t[299]);
  assign t[25] = ~(t[43] ^ t[44]);
  assign t[260] = (t[300] & ~t[301]);
  assign t[261] = (t[302] & ~t[303]);
  assign t[262] = (t[304] & ~t[305]);
  assign t[263] = (t[306] & ~t[307]);
  assign t[264] = (t[308] & ~t[309]);
  assign t[265] = (t[310] & ~t[311]);
  assign t[266] = (t[312] & ~t[313]);
  assign t[267] = (t[314] & ~t[315]);
  assign t[268] = (t[316] & ~t[317]);
  assign t[269] = (t[318] & ~t[319]);
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[270] = (t[320] & ~t[321]);
  assign t[271] = (t[322] & ~t[323]);
  assign t[272] = (t[324] & ~t[325]);
  assign t[273] = (t[326] & ~t[327]);
  assign t[274] = t[328] ^ x[4];
  assign t[275] = t[329] ^ x[3];
  assign t[276] = t[330] ^ x[9];
  assign t[277] = t[331] ^ x[8];
  assign t[278] = t[332] ^ x[12];
  assign t[279] = t[333] ^ x[11];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[334] ^ x[15];
  assign t[281] = t[335] ^ x[14];
  assign t[282] = t[336] ^ x[18];
  assign t[283] = t[337] ^ x[17];
  assign t[284] = t[338] ^ x[21];
  assign t[285] = t[339] ^ x[20];
  assign t[286] = t[340] ^ x[24];
  assign t[287] = t[341] ^ x[23];
  assign t[288] = t[342] ^ x[27];
  assign t[289] = t[343] ^ x[26];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[30];
  assign t[291] = t[345] ^ x[29];
  assign t[292] = t[346] ^ x[33];
  assign t[293] = t[347] ^ x[32];
  assign t[294] = t[348] ^ x[38];
  assign t[295] = t[349] ^ x[37];
  assign t[296] = t[350] ^ x[41];
  assign t[297] = t[351] ^ x[40];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[43];
  assign t[29] = ~(t[195]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[47];
  assign t[301] = t[355] ^ x[46];
  assign t[302] = t[356] ^ x[54];
  assign t[303] = t[357] ^ x[53];
  assign t[304] = t[358] ^ x[57];
  assign t[305] = t[359] ^ x[56];
  assign t[306] = t[360] ^ x[64];
  assign t[307] = t[361] ^ x[63];
  assign t[308] = t[362] ^ x[67];
  assign t[309] = t[363] ^ x[66];
  assign t[30] = ~(t[196]);
  assign t[310] = t[364] ^ x[70];
  assign t[311] = t[365] ^ x[69];
  assign t[312] = t[366] ^ x[73];
  assign t[313] = t[367] ^ x[72];
  assign t[314] = t[368] ^ x[76];
  assign t[315] = t[369] ^ x[75];
  assign t[316] = t[370] ^ x[79];
  assign t[317] = t[371] ^ x[78];
  assign t[318] = t[372] ^ x[82];
  assign t[319] = t[373] ^ x[81];
  assign t[31] = ~(t[197]);
  assign t[320] = t[374] ^ x[85];
  assign t[321] = t[375] ^ x[84];
  assign t[322] = t[376] ^ x[90];
  assign t[323] = t[377] ^ x[89];
  assign t[324] = t[378] ^ x[93];
  assign t[325] = t[379] ^ x[92];
  assign t[326] = t[380] ^ x[96];
  assign t[327] = t[381] ^ x[95];
  assign t[328] = (x[2]);
  assign t[329] = (x[2]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[7]);
  assign t[331] = (x[7]);
  assign t[332] = (x[10]);
  assign t[333] = (x[10]);
  assign t[334] = (x[13]);
  assign t[335] = (x[13]);
  assign t[336] = (x[16]);
  assign t[337] = (x[16]);
  assign t[338] = (x[19]);
  assign t[339] = (x[19]);
  assign t[33] = t[194] ^ t[52];
  assign t[340] = (x[22]);
  assign t[341] = (x[22]);
  assign t[342] = (x[25]);
  assign t[343] = (x[25]);
  assign t[344] = (x[28]);
  assign t[345] = (x[28]);
  assign t[346] = (x[31]);
  assign t[347] = (x[31]);
  assign t[348] = (x[36]);
  assign t[349] = (x[36]);
  assign t[34] = t[53] ^ t[22];
  assign t[350] = (x[39]);
  assign t[351] = (x[39]);
  assign t[352] = (x[42]);
  assign t[353] = (x[42]);
  assign t[354] = (x[45]);
  assign t[355] = (x[45]);
  assign t[356] = (x[52]);
  assign t[357] = (x[52]);
  assign t[358] = (x[55]);
  assign t[359] = (x[55]);
  assign t[35] = t[54] & t[55];
  assign t[360] = (x[62]);
  assign t[361] = (x[62]);
  assign t[362] = (x[65]);
  assign t[363] = (x[65]);
  assign t[364] = (x[68]);
  assign t[365] = (x[68]);
  assign t[366] = (x[71]);
  assign t[367] = (x[71]);
  assign t[368] = (x[74]);
  assign t[369] = (x[74]);
  assign t[36] = t[8] ? t[56] : t[198];
  assign t[370] = (x[77]);
  assign t[371] = (x[77]);
  assign t[372] = (x[80]);
  assign t[373] = (x[80]);
  assign t[374] = (x[83]);
  assign t[375] = (x[83]);
  assign t[376] = (x[88]);
  assign t[377] = (x[88]);
  assign t[378] = (x[91]);
  assign t[379] = (x[91]);
  assign t[37] = ~(t[57]);
  assign t[380] = (x[94]);
  assign t[381] = (x[94]);
  assign t[38] = t[8] ? t[58] : t[199];
  assign t[39] = ~t[59];
  assign t[3] = t[6] ^ t[7];
  assign t[40] = t[60] ^ t[61];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[66] ^ t[67]);
  assign t[44] = t[68] ^ t[69];
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[11] ^ t[72]);
  assign t[47] = ~(t[73] & t[74]);
  assign t[48] = t[200] | t[75];
  assign t[49] = ~(t[76]);
  assign t[4] = t[8] ? t[9] : t[193];
  assign t[50] = ~(t[201]);
  assign t[51] = ~(t[77] & t[202]);
  assign t[52] = t[78] ? x[35] : x[34];
  assign t[53] = t[79] & t[80];
  assign t[54] = ~(t[81] ^ t[34]);
  assign t[55] = t[68] ^ t[38];
  assign t[56] = t[198] ^ t[82];
  assign t[57] = t[8] ? t[83] : t[203];
  assign t[58] = t[199] ^ t[84];
  assign t[59] = t[27] ? t[85] : t[204];
  assign t[5] = ~(t[10]);
  assign t[60] = t[86] ^ t[87];
  assign t[61] = t[88] & t[89];
  assign t[62] = t[90] ^ t[39];
  assign t[63] = t[60] ^ t[91];
  assign t[64] = t[92] ^ t[93];
  assign t[65] = t[94] & t[95];
  assign t[66] = t[96] ^ t[23];
  assign t[67] = t[97] ^ t[98];
  assign t[68] = t[57] ^ t[19];
  assign t[69] = t[34] ^ t[99];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[100] ^ t[101];
  assign t[71] = t[102] ^ t[87];
  assign t[72] = t[103] ^ t[104];
  assign t[73] = ~(t[75] & t[105]);
  assign t[74] = ~(t[205] ^ t[106]);
  assign t[75] = ~(t[107] & t[108]);
  assign t[76] = ~(t[48]);
  assign t[77] = ~(t[206]);
  assign t[78] = ~(t[49]);
  assign t[79] = ~(t[109]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[36]);
  assign t[81] = t[36] ^ t[57];
  assign t[82] = t[78] ? x[49] : x[48];
  assign t[83] = t[203] ^ t[110];
  assign t[84] = t[78] ? x[51] : x[50];
  assign t[85] = t[204] ^ t[111];
  assign t[86] = t[112] & t[113];
  assign t[87] = t[114] & t[115];
  assign t[88] = ~(t[116] ^ t[60]);
  assign t[89] = t[62] ^ t[115];
  assign t[8] = ~(t[15]);
  assign t[90] = t[117];
  assign t[91] = t[118] & t[119];
  assign t[92] = t[8] ? t[120] : t[207];
  assign t[93] = t[195] ^ t[121];
  assign t[94] = ~(t[64] ^ t[122]);
  assign t[95] = t[123] ^ t[124];
  assign t[96] = t[123] ^ t[125];
  assign t[97] = t[126] ^ t[127];
  assign t[98] = t[128] & t[129];
  assign t[99] = t[130] & t[131];
  assign t[9] = t[193] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [116:0] x;
 output y;

 wire [370:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[57] ^ t[133];
  assign t[101] = t[134] & t[135];
  assign t[102] = ~(t[114] ^ t[68]);
  assign t[103] = t[136] ^ t[40];
  assign t[104] = t[137] ? x[65] : x[64];
  assign t[105] = t[137] ? x[67] : x[66];
  assign t[106] = t[138] & t[139];
  assign t[107] = t[194] ^ t[140];
  assign t[108] = ~(t[141] & t[142]);
  assign t[109] = t[143] ^ t[202];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[195]);
  assign t[111] = t[144] & t[143];
  assign t[112] = t[197] ^ t[145];
  assign t[113] = ~(t[45]);
  assign t[114] = t[37] ^ t[63];
  assign t[115] = t[146] ? t[147] : t[203];
  assign t[116] = t[118] ^ t[148];
  assign t[117] = t[146] ? t[149] : t[204];
  assign t[118] = t[150] ^ t[151];
  assign t[119] = t[152] & t[153];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[198] ^ t[154];
  assign t[121] = t[8] ? t[155] : t[205];
  assign t[122] = t[199] ^ t[156];
  assign t[123] = ~(t[157] ^ t[66]);
  assign t[124] = t[41] ^ t[90];
  assign t[125] = t[78] ? x[81] : x[80];
  assign t[126] = t[78] ? x[83] : x[82];
  assign t[127] = t[200] ^ t[158];
  assign t[128] = t[137] ? x[85] : x[84];
  assign t[129] = t[201] ^ t[159];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = ~(t[133]);
  assign t[131] = ~(t[88]);
  assign t[132] = t[41] ^ t[88];
  assign t[133] = t[90] ^ t[65];
  assign t[134] = ~(t[160]);
  assign t[135] = ~(t[37]);
  assign t[136] = t[63] ^ t[38];
  assign t[137] = ~(t[50]);
  assign t[138] = ~(t[161]);
  assign t[139] = ~(t[44]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[137] ? x[87] : x[86];
  assign t[141] = ~(t[144] | t[143]);
  assign t[142] = ~(t[162] | t[110]);
  assign t[143] = ~(t[206]);
  assign t[144] = ~(t[202]);
  assign t[145] = t[137] ? x[92] : x[91];
  assign t[146] = ~(t[15]);
  assign t[147] = t[203] ^ t[163];
  assign t[148] = t[164] & t[165];
  assign t[149] = t[204] ^ t[166];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[167] & t[168];
  assign t[151] = t[169] & t[170];
  assign t[152] = ~(t[150] ^ t[171]);
  assign t[153] = t[172] ^ t[173];
  assign t[154] = t[78] ? x[94] : x[93];
  assign t[155] = t[205] ^ t[174];
  assign t[156] = t[78] ? x[96] : x[95];
  assign t[157] = t[88] ^ t[65];
  assign t[158] = t[28] ? x[98] : x[97];
  assign t[159] = t[28] ? x[100] : x[99];
  assign t[15] = ~(t[27]);
  assign t[160] = t[40] ^ t[63];
  assign t[161] = t[74] ^ t[45];
  assign t[162] = ~(t[188]);
  assign t[163] = t[175] ? x[102] : x[101];
  assign t[164] = ~(t[176] ^ t[118]);
  assign t[165] = t[86] ^ t[170];
  assign t[166] = t[175] ? x[104] : x[103];
  assign t[167] = ~(t[173]);
  assign t[168] = ~(t[177]);
  assign t[169] = ~(t[117]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[146] ? t[178] : t[207];
  assign t[171] = t[86] ^ t[177];
  assign t[172] = t[177] ^ t[115];
  assign t[173] = t[170] ^ t[117];
  assign t[174] = t[28] ? x[109] : x[108];
  assign t[175] = ~(t[50]);
  assign t[176] = t[177] ^ t[117];
  assign t[177] = t[146] ? t[179] : t[208];
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[208] ^ t[181];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[175] ? x[114] : x[113];
  assign t[181] = t[175] ? x[116] : x[115];
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = t[236] ^ x[4];
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = t[237] ^ x[9];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[60];
  assign t[228] = t[255] ^ x[63];
  assign t[229] = t[256] ^ x[70];
  assign t[22] = t[39] & t[40];
  assign t[230] = t[257] ^ x[73];
  assign t[231] = t[258] ^ x[76];
  assign t[232] = t[259] ^ x[79];
  assign t[233] = t[260] ^ x[90];
  assign t[234] = t[261] ^ x[107];
  assign t[235] = t[262] ^ x[112];
  assign t[236] = (t[263] & ~t[264]);
  assign t[237] = (t[265] & ~t[266]);
  assign t[238] = (t[267] & ~t[268]);
  assign t[239] = (t[269] & ~t[270]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (t[271] & ~t[272]);
  assign t[241] = (t[273] & ~t[274]);
  assign t[242] = (t[275] & ~t[276]);
  assign t[243] = (t[277] & ~t[278]);
  assign t[244] = (t[279] & ~t[280]);
  assign t[245] = (t[281] & ~t[282]);
  assign t[246] = (t[283] & ~t[284]);
  assign t[247] = (t[285] & ~t[286]);
  assign t[248] = (t[287] & ~t[288]);
  assign t[249] = (t[289] & ~t[290]);
  assign t[24] = t[38] ^ t[43];
  assign t[250] = (t[291] & ~t[292]);
  assign t[251] = (t[293] & ~t[294]);
  assign t[252] = (t[295] & ~t[296]);
  assign t[253] = (t[297] & ~t[298]);
  assign t[254] = (t[299] & ~t[300]);
  assign t[255] = (t[301] & ~t[302]);
  assign t[256] = (t[303] & ~t[304]);
  assign t[257] = (t[305] & ~t[306]);
  assign t[258] = (t[307] & ~t[308]);
  assign t[259] = (t[309] & ~t[310]);
  assign t[25] = t[44] ^ t[45];
  assign t[260] = (t[311] & ~t[312]);
  assign t[261] = (t[313] & ~t[314]);
  assign t[262] = (t[315] & ~t[316]);
  assign t[263] = t[317] ^ x[4];
  assign t[264] = t[318] ^ x[3];
  assign t[265] = t[319] ^ x[9];
  assign t[266] = t[320] ^ x[8];
  assign t[267] = t[321] ^ x[12];
  assign t[268] = t[322] ^ x[11];
  assign t[269] = t[323] ^ x[15];
  assign t[26] = t[46] & t[47];
  assign t[270] = t[324] ^ x[14];
  assign t[271] = t[325] ^ x[18];
  assign t[272] = t[326] ^ x[17];
  assign t[273] = t[327] ^ x[21];
  assign t[274] = t[328] ^ x[20];
  assign t[275] = t[329] ^ x[24];
  assign t[276] = t[330] ^ x[23];
  assign t[277] = t[331] ^ x[27];
  assign t[278] = t[332] ^ x[26];
  assign t[279] = t[333] ^ x[30];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[29];
  assign t[281] = t[335] ^ x[33];
  assign t[282] = t[336] ^ x[32];
  assign t[283] = t[337] ^ x[36];
  assign t[284] = t[338] ^ x[35];
  assign t[285] = t[339] ^ x[39];
  assign t[286] = t[340] ^ x[38];
  assign t[287] = t[341] ^ x[42];
  assign t[288] = t[342] ^ x[41];
  assign t[289] = t[343] ^ x[45];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[44];
  assign t[291] = t[345] ^ x[48];
  assign t[292] = t[346] ^ x[47];
  assign t[293] = t[347] ^ x[51];
  assign t[294] = t[348] ^ x[50];
  assign t[295] = t[349] ^ x[54];
  assign t[296] = t[350] ^ x[53];
  assign t[297] = t[351] ^ x[57];
  assign t[298] = t[352] ^ x[56];
  assign t[299] = t[353] ^ x[60];
  assign t[29] = ~(t[183]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[59];
  assign t[301] = t[355] ^ x[63];
  assign t[302] = t[356] ^ x[62];
  assign t[303] = t[357] ^ x[70];
  assign t[304] = t[358] ^ x[69];
  assign t[305] = t[359] ^ x[73];
  assign t[306] = t[360] ^ x[72];
  assign t[307] = t[361] ^ x[76];
  assign t[308] = t[362] ^ x[75];
  assign t[309] = t[363] ^ x[79];
  assign t[30] = ~(t[184]);
  assign t[310] = t[364] ^ x[78];
  assign t[311] = t[365] ^ x[90];
  assign t[312] = t[366] ^ x[89];
  assign t[313] = t[367] ^ x[107];
  assign t[314] = t[368] ^ x[106];
  assign t[315] = t[369] ^ x[112];
  assign t[316] = t[370] ^ x[111];
  assign t[317] = (x[2]);
  assign t[318] = (x[2]);
  assign t[319] = (x[7]);
  assign t[31] = ~(t[185]);
  assign t[320] = (x[7]);
  assign t[321] = (x[10]);
  assign t[322] = (x[10]);
  assign t[323] = (x[13]);
  assign t[324] = (x[13]);
  assign t[325] = (x[16]);
  assign t[326] = (x[16]);
  assign t[327] = (x[19]);
  assign t[328] = (x[19]);
  assign t[329] = (x[22]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[22]);
  assign t[331] = (x[25]);
  assign t[332] = (x[25]);
  assign t[333] = (x[28]);
  assign t[334] = (x[28]);
  assign t[335] = (x[31]);
  assign t[336] = (x[31]);
  assign t[337] = (x[34]);
  assign t[338] = (x[34]);
  assign t[339] = (x[37]);
  assign t[33] = t[53] ^ t[54];
  assign t[340] = (x[37]);
  assign t[341] = (x[40]);
  assign t[342] = (x[40]);
  assign t[343] = (x[43]);
  assign t[344] = (x[43]);
  assign t[345] = (x[46]);
  assign t[346] = (x[46]);
  assign t[347] = (x[49]);
  assign t[348] = (x[49]);
  assign t[349] = (x[52]);
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[350] = (x[52]);
  assign t[351] = (x[55]);
  assign t[352] = (x[55]);
  assign t[353] = (x[58]);
  assign t[354] = (x[58]);
  assign t[355] = (x[61]);
  assign t[356] = (x[61]);
  assign t[357] = (x[68]);
  assign t[358] = (x[68]);
  assign t[359] = (x[71]);
  assign t[35] = t[57] ^ t[58];
  assign t[360] = (x[71]);
  assign t[361] = (x[74]);
  assign t[362] = (x[74]);
  assign t[363] = (x[77]);
  assign t[364] = (x[77]);
  assign t[365] = (x[88]);
  assign t[366] = (x[88]);
  assign t[367] = (x[105]);
  assign t[368] = (x[105]);
  assign t[369] = (x[110]);
  assign t[36] = t[59] ^ t[60];
  assign t[370] = (x[110]);
  assign t[37] = ~t[61];
  assign t[38] = ~t[62];
  assign t[39] = ~(t[63]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64];
  assign t[41] = t[65] ^ t[59];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[8] ? t[70] : t[186];
  assign t[45] = t[8] ? t[71] : t[187];
  assign t[46] = ~(t[25] ^ t[72]);
  assign t[47] = t[73] ^ t[74];
  assign t[48] = ~(t[75] & t[76]);
  assign t[49] = t[188] | t[77];
  assign t[4] = t[8] ? t[9] : t[182];
  assign t[50] = ~(t[78]);
  assign t[51] = ~(t[189]);
  assign t[52] = ~(t[79] & t[190]);
  assign t[53] = t[80] ^ t[81];
  assign t[54] = t[82] ^ t[83];
  assign t[55] = ~(t[84] ^ t[85]);
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ^ t[59];
  assign t[58] = t[89] & t[90];
  assign t[59] = t[190] ^ t[91];
  assign t[5] = ~(t[10]);
  assign t[60] = t[66] ^ t[92];
  assign t[61] = t[27] ? t[93] : t[191];
  assign t[62] = t[27] ? t[94] : t[192];
  assign t[63] = t[95];
  assign t[64] = t[27] ? t[96] : t[193];
  assign t[65] = t[183] ^ t[97];
  assign t[66] = t[98] ^ t[58];
  assign t[67] = t[99] & t[100];
  assign t[68] = t[101] ^ t[22];
  assign t[69] = t[102] & t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[186] ^ t[104];
  assign t[71] = t[187] ^ t[105];
  assign t[72] = t[106] ^ t[83];
  assign t[73] = t[45] ^ t[80];
  assign t[74] = t[8] ? t[107] : t[194];
  assign t[75] = ~(t[77] & t[108]);
  assign t[76] = ~(t[195] ^ t[109]);
  assign t[77] = ~(t[110] & t[111]);
  assign t[78] = ~(t[49]);
  assign t[79] = ~(t[196]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[112] : t[197];
  assign t[81] = t[72] ^ t[26];
  assign t[82] = t[44] ^ t[80];
  assign t[83] = t[113] & t[74];
  assign t[84] = t[114] ^ t[69];
  assign t[85] = t[115] ^ t[116];
  assign t[86] = t[117] ^ t[115];
  assign t[87] = t[118] ^ t[119];
  assign t[88] = t[8] ? t[120] : t[198];
  assign t[89] = ~(t[65]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[184] ^ t[121];
  assign t[91] = t[8] ? t[122] : t[199];
  assign t[92] = t[123] & t[124];
  assign t[93] = t[191] ^ t[125];
  assign t[94] = t[192] ^ t[126];
  assign t[95] = t[27] ? t[127] : t[200];
  assign t[96] = t[193] ^ t[128];
  assign t[97] = t[27] ? t[129] : t[201];
  assign t[98] = t[130] & t[131];
  assign t[99] = ~(t[98] ^ t[132]);
  assign t[9] = t[182] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [116:0] x;
 output y;

 wire [370:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[57] ^ t[133];
  assign t[101] = t[134] & t[135];
  assign t[102] = ~(t[114] ^ t[68]);
  assign t[103] = t[136] ^ t[40];
  assign t[104] = t[137] ? x[65] : x[64];
  assign t[105] = t[137] ? x[67] : x[66];
  assign t[106] = t[138] & t[139];
  assign t[107] = t[194] ^ t[140];
  assign t[108] = ~(t[141] & t[142]);
  assign t[109] = t[143] ^ t[202];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[195]);
  assign t[111] = t[144] & t[143];
  assign t[112] = t[197] ^ t[145];
  assign t[113] = ~(t[45]);
  assign t[114] = t[37] ^ t[63];
  assign t[115] = t[146] ? t[147] : t[203];
  assign t[116] = t[118] ^ t[148];
  assign t[117] = t[146] ? t[149] : t[204];
  assign t[118] = t[150] ^ t[151];
  assign t[119] = t[152] & t[153];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[198] ^ t[154];
  assign t[121] = t[8] ? t[155] : t[205];
  assign t[122] = t[199] ^ t[156];
  assign t[123] = ~(t[157] ^ t[66]);
  assign t[124] = t[41] ^ t[90];
  assign t[125] = t[78] ? x[81] : x[80];
  assign t[126] = t[78] ? x[83] : x[82];
  assign t[127] = t[200] ^ t[158];
  assign t[128] = t[137] ? x[85] : x[84];
  assign t[129] = t[201] ^ t[159];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = ~(t[133]);
  assign t[131] = ~(t[88]);
  assign t[132] = t[41] ^ t[88];
  assign t[133] = t[90] ^ t[65];
  assign t[134] = ~(t[160]);
  assign t[135] = ~(t[37]);
  assign t[136] = t[63] ^ t[38];
  assign t[137] = ~(t[50]);
  assign t[138] = ~(t[161]);
  assign t[139] = ~(t[44]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[137] ? x[87] : x[86];
  assign t[141] = ~(t[144] | t[143]);
  assign t[142] = ~(t[162] | t[110]);
  assign t[143] = ~(t[206]);
  assign t[144] = ~(t[202]);
  assign t[145] = t[137] ? x[92] : x[91];
  assign t[146] = ~(t[15]);
  assign t[147] = t[203] ^ t[163];
  assign t[148] = t[164] & t[165];
  assign t[149] = t[204] ^ t[166];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[167] & t[168];
  assign t[151] = t[169] & t[170];
  assign t[152] = ~(t[150] ^ t[171]);
  assign t[153] = t[172] ^ t[173];
  assign t[154] = t[78] ? x[94] : x[93];
  assign t[155] = t[205] ^ t[174];
  assign t[156] = t[78] ? x[96] : x[95];
  assign t[157] = t[88] ^ t[65];
  assign t[158] = t[28] ? x[98] : x[97];
  assign t[159] = t[28] ? x[100] : x[99];
  assign t[15] = ~(t[27]);
  assign t[160] = t[40] ^ t[63];
  assign t[161] = t[74] ^ t[45];
  assign t[162] = ~(t[188]);
  assign t[163] = t[175] ? x[102] : x[101];
  assign t[164] = ~(t[176] ^ t[118]);
  assign t[165] = t[86] ^ t[170];
  assign t[166] = t[175] ? x[104] : x[103];
  assign t[167] = ~(t[173]);
  assign t[168] = ~(t[177]);
  assign t[169] = ~(t[117]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[146] ? t[178] : t[207];
  assign t[171] = t[86] ^ t[177];
  assign t[172] = t[177] ^ t[115];
  assign t[173] = t[170] ^ t[117];
  assign t[174] = t[28] ? x[109] : x[108];
  assign t[175] = ~(t[50]);
  assign t[176] = t[177] ^ t[117];
  assign t[177] = t[146] ? t[179] : t[208];
  assign t[178] = t[207] ^ t[180];
  assign t[179] = t[208] ^ t[181];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[175] ? x[114] : x[113];
  assign t[181] = t[175] ? x[116] : x[115];
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = t[236] ^ x[4];
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = t[237] ^ x[9];
  assign t[211] = t[238] ^ x[12];
  assign t[212] = t[239] ^ x[15];
  assign t[213] = t[240] ^ x[18];
  assign t[214] = t[241] ^ x[21];
  assign t[215] = t[242] ^ x[24];
  assign t[216] = t[243] ^ x[27];
  assign t[217] = t[244] ^ x[30];
  assign t[218] = t[245] ^ x[33];
  assign t[219] = t[246] ^ x[36];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[39];
  assign t[221] = t[248] ^ x[42];
  assign t[222] = t[249] ^ x[45];
  assign t[223] = t[250] ^ x[48];
  assign t[224] = t[251] ^ x[51];
  assign t[225] = t[252] ^ x[54];
  assign t[226] = t[253] ^ x[57];
  assign t[227] = t[254] ^ x[60];
  assign t[228] = t[255] ^ x[63];
  assign t[229] = t[256] ^ x[70];
  assign t[22] = t[39] & t[40];
  assign t[230] = t[257] ^ x[73];
  assign t[231] = t[258] ^ x[76];
  assign t[232] = t[259] ^ x[79];
  assign t[233] = t[260] ^ x[90];
  assign t[234] = t[261] ^ x[107];
  assign t[235] = t[262] ^ x[112];
  assign t[236] = (t[263] & ~t[264]);
  assign t[237] = (t[265] & ~t[266]);
  assign t[238] = (t[267] & ~t[268]);
  assign t[239] = (t[269] & ~t[270]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (t[271] & ~t[272]);
  assign t[241] = (t[273] & ~t[274]);
  assign t[242] = (t[275] & ~t[276]);
  assign t[243] = (t[277] & ~t[278]);
  assign t[244] = (t[279] & ~t[280]);
  assign t[245] = (t[281] & ~t[282]);
  assign t[246] = (t[283] & ~t[284]);
  assign t[247] = (t[285] & ~t[286]);
  assign t[248] = (t[287] & ~t[288]);
  assign t[249] = (t[289] & ~t[290]);
  assign t[24] = t[38] ^ t[43];
  assign t[250] = (t[291] & ~t[292]);
  assign t[251] = (t[293] & ~t[294]);
  assign t[252] = (t[295] & ~t[296]);
  assign t[253] = (t[297] & ~t[298]);
  assign t[254] = (t[299] & ~t[300]);
  assign t[255] = (t[301] & ~t[302]);
  assign t[256] = (t[303] & ~t[304]);
  assign t[257] = (t[305] & ~t[306]);
  assign t[258] = (t[307] & ~t[308]);
  assign t[259] = (t[309] & ~t[310]);
  assign t[25] = t[44] ^ t[45];
  assign t[260] = (t[311] & ~t[312]);
  assign t[261] = (t[313] & ~t[314]);
  assign t[262] = (t[315] & ~t[316]);
  assign t[263] = t[317] ^ x[4];
  assign t[264] = t[318] ^ x[3];
  assign t[265] = t[319] ^ x[9];
  assign t[266] = t[320] ^ x[8];
  assign t[267] = t[321] ^ x[12];
  assign t[268] = t[322] ^ x[11];
  assign t[269] = t[323] ^ x[15];
  assign t[26] = t[46] & t[47];
  assign t[270] = t[324] ^ x[14];
  assign t[271] = t[325] ^ x[18];
  assign t[272] = t[326] ^ x[17];
  assign t[273] = t[327] ^ x[21];
  assign t[274] = t[328] ^ x[20];
  assign t[275] = t[329] ^ x[24];
  assign t[276] = t[330] ^ x[23];
  assign t[277] = t[331] ^ x[27];
  assign t[278] = t[332] ^ x[26];
  assign t[279] = t[333] ^ x[30];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[29];
  assign t[281] = t[335] ^ x[33];
  assign t[282] = t[336] ^ x[32];
  assign t[283] = t[337] ^ x[36];
  assign t[284] = t[338] ^ x[35];
  assign t[285] = t[339] ^ x[39];
  assign t[286] = t[340] ^ x[38];
  assign t[287] = t[341] ^ x[42];
  assign t[288] = t[342] ^ x[41];
  assign t[289] = t[343] ^ x[45];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[44];
  assign t[291] = t[345] ^ x[48];
  assign t[292] = t[346] ^ x[47];
  assign t[293] = t[347] ^ x[51];
  assign t[294] = t[348] ^ x[50];
  assign t[295] = t[349] ^ x[54];
  assign t[296] = t[350] ^ x[53];
  assign t[297] = t[351] ^ x[57];
  assign t[298] = t[352] ^ x[56];
  assign t[299] = t[353] ^ x[60];
  assign t[29] = ~(t[183]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[59];
  assign t[301] = t[355] ^ x[63];
  assign t[302] = t[356] ^ x[62];
  assign t[303] = t[357] ^ x[70];
  assign t[304] = t[358] ^ x[69];
  assign t[305] = t[359] ^ x[73];
  assign t[306] = t[360] ^ x[72];
  assign t[307] = t[361] ^ x[76];
  assign t[308] = t[362] ^ x[75];
  assign t[309] = t[363] ^ x[79];
  assign t[30] = ~(t[184]);
  assign t[310] = t[364] ^ x[78];
  assign t[311] = t[365] ^ x[90];
  assign t[312] = t[366] ^ x[89];
  assign t[313] = t[367] ^ x[107];
  assign t[314] = t[368] ^ x[106];
  assign t[315] = t[369] ^ x[112];
  assign t[316] = t[370] ^ x[111];
  assign t[317] = (x[2]);
  assign t[318] = (x[2]);
  assign t[319] = (x[7]);
  assign t[31] = ~(t[185]);
  assign t[320] = (x[7]);
  assign t[321] = (x[10]);
  assign t[322] = (x[10]);
  assign t[323] = (x[13]);
  assign t[324] = (x[13]);
  assign t[325] = (x[16]);
  assign t[326] = (x[16]);
  assign t[327] = (x[19]);
  assign t[328] = (x[19]);
  assign t[329] = (x[22]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[22]);
  assign t[331] = (x[25]);
  assign t[332] = (x[25]);
  assign t[333] = (x[28]);
  assign t[334] = (x[28]);
  assign t[335] = (x[31]);
  assign t[336] = (x[31]);
  assign t[337] = (x[34]);
  assign t[338] = (x[34]);
  assign t[339] = (x[37]);
  assign t[33] = t[53] ^ t[54];
  assign t[340] = (x[37]);
  assign t[341] = (x[40]);
  assign t[342] = (x[40]);
  assign t[343] = (x[43]);
  assign t[344] = (x[43]);
  assign t[345] = (x[46]);
  assign t[346] = (x[46]);
  assign t[347] = (x[49]);
  assign t[348] = (x[49]);
  assign t[349] = (x[52]);
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[350] = (x[52]);
  assign t[351] = (x[55]);
  assign t[352] = (x[55]);
  assign t[353] = (x[58]);
  assign t[354] = (x[58]);
  assign t[355] = (x[61]);
  assign t[356] = (x[61]);
  assign t[357] = (x[68]);
  assign t[358] = (x[68]);
  assign t[359] = (x[71]);
  assign t[35] = t[57] ^ t[58];
  assign t[360] = (x[71]);
  assign t[361] = (x[74]);
  assign t[362] = (x[74]);
  assign t[363] = (x[77]);
  assign t[364] = (x[77]);
  assign t[365] = (x[88]);
  assign t[366] = (x[88]);
  assign t[367] = (x[105]);
  assign t[368] = (x[105]);
  assign t[369] = (x[110]);
  assign t[36] = t[59] ^ t[60];
  assign t[370] = (x[110]);
  assign t[37] = ~t[61];
  assign t[38] = ~t[62];
  assign t[39] = ~(t[63]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64];
  assign t[41] = t[65] ^ t[59];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[8] ? t[70] : t[186];
  assign t[45] = t[8] ? t[71] : t[187];
  assign t[46] = ~(t[25] ^ t[72]);
  assign t[47] = t[73] ^ t[74];
  assign t[48] = ~(t[75] & t[76]);
  assign t[49] = t[188] | t[77];
  assign t[4] = t[8] ? t[9] : t[182];
  assign t[50] = ~(t[78]);
  assign t[51] = ~(t[189]);
  assign t[52] = ~(t[79] & t[190]);
  assign t[53] = t[80] ^ t[81];
  assign t[54] = t[82] ^ t[83];
  assign t[55] = ~(t[84] ^ t[85]);
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ^ t[59];
  assign t[58] = t[89] & t[90];
  assign t[59] = t[190] ^ t[91];
  assign t[5] = ~(t[10]);
  assign t[60] = t[66] ^ t[92];
  assign t[61] = t[27] ? t[93] : t[191];
  assign t[62] = t[27] ? t[94] : t[192];
  assign t[63] = t[95];
  assign t[64] = t[27] ? t[96] : t[193];
  assign t[65] = t[183] ^ t[97];
  assign t[66] = t[98] ^ t[58];
  assign t[67] = t[99] & t[100];
  assign t[68] = t[101] ^ t[22];
  assign t[69] = t[102] & t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[186] ^ t[104];
  assign t[71] = t[187] ^ t[105];
  assign t[72] = t[106] ^ t[83];
  assign t[73] = t[45] ^ t[80];
  assign t[74] = t[8] ? t[107] : t[194];
  assign t[75] = ~(t[77] & t[108]);
  assign t[76] = ~(t[195] ^ t[109]);
  assign t[77] = ~(t[110] & t[111]);
  assign t[78] = ~(t[49]);
  assign t[79] = ~(t[196]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[112] : t[197];
  assign t[81] = t[72] ^ t[26];
  assign t[82] = t[44] ^ t[80];
  assign t[83] = t[113] & t[74];
  assign t[84] = t[114] ^ t[69];
  assign t[85] = t[115] ^ t[116];
  assign t[86] = t[117] ^ t[115];
  assign t[87] = t[118] ^ t[119];
  assign t[88] = t[8] ? t[120] : t[198];
  assign t[89] = ~(t[65]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[184] ^ t[121];
  assign t[91] = t[8] ? t[122] : t[199];
  assign t[92] = t[123] & t[124];
  assign t[93] = t[191] ^ t[125];
  assign t[94] = t[192] ^ t[126];
  assign t[95] = t[27] ? t[127] : t[200];
  assign t[96] = t[193] ^ t[128];
  assign t[97] = t[27] ? t[129] : t[201];
  assign t[98] = t[130] & t[131];
  assign t[99] = ~(t[98] ^ t[132]);
  assign t[9] = t[182] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind86(x, y);
 input [116:0] x;
 output y;

 wire [361:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[137] ? x[62] : x[61];
  assign t[101] = t[137] ? x[64] : x[63];
  assign t[102] = ~(t[108]);
  assign t[103] = ~(t[85]);
  assign t[104] = ~(t[41]);
  assign t[105] = t[8] ? t[138] : t[192];
  assign t[106] = t[23] ^ t[85];
  assign t[107] = t[85] ^ t[42];
  assign t[108] = t[105] ^ t[41];
  assign t[109] = t[80] ? x[69] : x[68];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[139]);
  assign t[111] = ~(t[124]);
  assign t[112] = ~(t[125]);
  assign t[113] = t[176] ^ t[140];
  assign t[114] = t[125] ^ t[25];
  assign t[115] = ~(t[141] & t[142]);
  assign t[116] = t[143] ^ t[193];
  assign t[117] = ~(t[186]);
  assign t[118] = t[144] & t[143];
  assign t[119] = t[188] ^ t[145];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[90] ? t[146] : t[194];
  assign t[121] = t[189] ^ t[147];
  assign t[122] = t[190] ^ t[148];
  assign t[123] = t[149] & t[150];
  assign t[124] = t[8] ? t[151] : t[195];
  assign t[125] = t[175] ^ t[152];
  assign t[126] = t[153] ? x[80] : x[79];
  assign t[127] = t[154] & t[155];
  assign t[128] = ~(t[156] ^ t[92]);
  assign t[129] = t[157] ^ t[84];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[80] ? x[82] : x[81];
  assign t[131] = t[28] ? x[84] : x[83];
  assign t[132] = ~(t[158]);
  assign t[133] = ~(t[37]);
  assign t[134] = ~(t[38]);
  assign t[135] = t[27] ? t[159] : t[196];
  assign t[136] = t[191] ^ t[160];
  assign t[137] = ~(t[50]);
  assign t[138] = t[192] ^ t[161];
  assign t[139] = t[113] ^ t[125];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[8] ? t[162] : t[197];
  assign t[141] = ~(t[144] | t[143]);
  assign t[142] = ~(t[163] | t[117]);
  assign t[143] = ~(t[198]);
  assign t[144] = ~(t[193]);
  assign t[145] = t[153] ? x[95] : x[94];
  assign t[146] = t[194] ^ t[164];
  assign t[147] = t[153] ? x[97] : x[96];
  assign t[148] = t[137] ? x[99] : x[98];
  assign t[149] = ~(t[96] ^ t[165]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[166] ^ t[158];
  assign t[151] = t[195] ^ t[167];
  assign t[152] = t[27] ? t[168] : t[199];
  assign t[153] = ~(t[50]);
  assign t[154] = ~(t[169]);
  assign t[155] = ~(t[82]);
  assign t[156] = t[82] ^ t[120];
  assign t[157] = t[120] ^ t[59];
  assign t[158] = t[65] ^ t[38];
  assign t[159] = t[196] ^ t[170];
  assign t[15] = ~(t[27]);
  assign t[160] = t[137] ? x[104] : x[103];
  assign t[161] = t[137] ? x[106] : x[105];
  assign t[162] = t[197] ^ t[171];
  assign t[163] = ~(t[181]);
  assign t[164] = t[153] ? x[108] : x[107];
  assign t[165] = t[64] ^ t[37];
  assign t[166] = t[37] ^ t[98];
  assign t[167] = t[80] ? x[110] : x[109];
  assign t[168] = t[199] ^ t[172];
  assign t[169] = t[84] ^ t[120];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[80] ? x[112] : x[111];
  assign t[171] = t[28] ? x[114] : x[113];
  assign t[172] = t[28] ? x[116] : x[115];
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[4];
  assign t[201] = t[228] ^ x[9];
  assign t[202] = t[229] ^ x[12];
  assign t[203] = t[230] ^ x[15];
  assign t[204] = t[231] ^ x[18];
  assign t[205] = t[232] ^ x[21];
  assign t[206] = t[233] ^ x[24];
  assign t[207] = t[234] ^ x[27];
  assign t[208] = t[235] ^ x[30];
  assign t[209] = t[236] ^ x[33];
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = t[237] ^ x[36];
  assign t[211] = t[238] ^ x[39];
  assign t[212] = t[239] ^ x[42];
  assign t[213] = t[240] ^ x[45];
  assign t[214] = t[241] ^ x[48];
  assign t[215] = t[242] ^ x[51];
  assign t[216] = t[243] ^ x[54];
  assign t[217] = t[244] ^ x[57];
  assign t[218] = t[245] ^ x[60];
  assign t[219] = t[246] ^ x[67];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[72];
  assign t[221] = t[248] ^ x[75];
  assign t[222] = t[249] ^ x[78];
  assign t[223] = t[250] ^ x[87];
  assign t[224] = t[251] ^ x[90];
  assign t[225] = t[252] ^ x[93];
  assign t[226] = t[253] ^ x[102];
  assign t[227] = (t[254] & ~t[255]);
  assign t[228] = (t[256] & ~t[257]);
  assign t[229] = (t[258] & ~t[259]);
  assign t[22] = t[39] & t[40];
  assign t[230] = (t[260] & ~t[261]);
  assign t[231] = (t[262] & ~t[263]);
  assign t[232] = (t[264] & ~t[265]);
  assign t[233] = (t[266] & ~t[267]);
  assign t[234] = (t[268] & ~t[269]);
  assign t[235] = (t[270] & ~t[271]);
  assign t[236] = (t[272] & ~t[273]);
  assign t[237] = (t[274] & ~t[275]);
  assign t[238] = (t[276] & ~t[277]);
  assign t[239] = (t[278] & ~t[279]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (t[280] & ~t[281]);
  assign t[241] = (t[282] & ~t[283]);
  assign t[242] = (t[284] & ~t[285]);
  assign t[243] = (t[286] & ~t[287]);
  assign t[244] = (t[288] & ~t[289]);
  assign t[245] = (t[290] & ~t[291]);
  assign t[246] = (t[292] & ~t[293]);
  assign t[247] = (t[294] & ~t[295]);
  assign t[248] = (t[296] & ~t[297]);
  assign t[249] = (t[298] & ~t[299]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (t[300] & ~t[301]);
  assign t[251] = (t[302] & ~t[303]);
  assign t[252] = (t[304] & ~t[305]);
  assign t[253] = (t[306] & ~t[307]);
  assign t[254] = t[308] ^ x[4];
  assign t[255] = t[309] ^ x[3];
  assign t[256] = t[310] ^ x[9];
  assign t[257] = t[311] ^ x[8];
  assign t[258] = t[312] ^ x[12];
  assign t[259] = t[313] ^ x[11];
  assign t[25] = t[174] ^ t[45];
  assign t[260] = t[314] ^ x[15];
  assign t[261] = t[315] ^ x[14];
  assign t[262] = t[316] ^ x[18];
  assign t[263] = t[317] ^ x[17];
  assign t[264] = t[318] ^ x[21];
  assign t[265] = t[319] ^ x[20];
  assign t[266] = t[320] ^ x[24];
  assign t[267] = t[321] ^ x[23];
  assign t[268] = t[322] ^ x[27];
  assign t[269] = t[323] ^ x[26];
  assign t[26] = t[46] ^ t[47];
  assign t[270] = t[324] ^ x[30];
  assign t[271] = t[325] ^ x[29];
  assign t[272] = t[326] ^ x[33];
  assign t[273] = t[327] ^ x[32];
  assign t[274] = t[328] ^ x[36];
  assign t[275] = t[329] ^ x[35];
  assign t[276] = t[330] ^ x[39];
  assign t[277] = t[331] ^ x[38];
  assign t[278] = t[332] ^ x[42];
  assign t[279] = t[333] ^ x[41];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[45];
  assign t[281] = t[335] ^ x[44];
  assign t[282] = t[336] ^ x[48];
  assign t[283] = t[337] ^ x[47];
  assign t[284] = t[338] ^ x[51];
  assign t[285] = t[339] ^ x[50];
  assign t[286] = t[340] ^ x[54];
  assign t[287] = t[341] ^ x[53];
  assign t[288] = t[342] ^ x[57];
  assign t[289] = t[343] ^ x[56];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[60];
  assign t[291] = t[345] ^ x[59];
  assign t[292] = t[346] ^ x[67];
  assign t[293] = t[347] ^ x[66];
  assign t[294] = t[348] ^ x[72];
  assign t[295] = t[349] ^ x[71];
  assign t[296] = t[350] ^ x[75];
  assign t[297] = t[351] ^ x[74];
  assign t[298] = t[352] ^ x[78];
  assign t[299] = t[353] ^ x[77];
  assign t[29] = ~(t[175]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[87];
  assign t[301] = t[355] ^ x[86];
  assign t[302] = t[356] ^ x[90];
  assign t[303] = t[357] ^ x[89];
  assign t[304] = t[358] ^ x[93];
  assign t[305] = t[359] ^ x[92];
  assign t[306] = t[360] ^ x[102];
  assign t[307] = t[361] ^ x[101];
  assign t[308] = (x[2]);
  assign t[309] = (x[2]);
  assign t[30] = ~(t[176]);
  assign t[310] = (x[7]);
  assign t[311] = (x[7]);
  assign t[312] = (x[10]);
  assign t[313] = (x[10]);
  assign t[314] = (x[13]);
  assign t[315] = (x[13]);
  assign t[316] = (x[16]);
  assign t[317] = (x[16]);
  assign t[318] = (x[19]);
  assign t[319] = (x[19]);
  assign t[31] = ~(t[177]);
  assign t[320] = (x[22]);
  assign t[321] = (x[22]);
  assign t[322] = (x[25]);
  assign t[323] = (x[25]);
  assign t[324] = (x[28]);
  assign t[325] = (x[28]);
  assign t[326] = (x[31]);
  assign t[327] = (x[31]);
  assign t[328] = (x[34]);
  assign t[329] = (x[34]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[37]);
  assign t[331] = (x[37]);
  assign t[332] = (x[40]);
  assign t[333] = (x[40]);
  assign t[334] = (x[43]);
  assign t[335] = (x[43]);
  assign t[336] = (x[46]);
  assign t[337] = (x[46]);
  assign t[338] = (x[49]);
  assign t[339] = (x[49]);
  assign t[33] = t[53] ^ t[54];
  assign t[340] = (x[52]);
  assign t[341] = (x[52]);
  assign t[342] = (x[55]);
  assign t[343] = (x[55]);
  assign t[344] = (x[58]);
  assign t[345] = (x[58]);
  assign t[346] = (x[65]);
  assign t[347] = (x[65]);
  assign t[348] = (x[70]);
  assign t[349] = (x[70]);
  assign t[34] = t[55] ^ t[56];
  assign t[350] = (x[73]);
  assign t[351] = (x[73]);
  assign t[352] = (x[76]);
  assign t[353] = (x[76]);
  assign t[354] = (x[85]);
  assign t[355] = (x[85]);
  assign t[356] = (x[88]);
  assign t[357] = (x[88]);
  assign t[358] = (x[91]);
  assign t[359] = (x[91]);
  assign t[35] = t[57] ^ t[58];
  assign t[360] = (x[100]);
  assign t[361] = (x[100]);
  assign t[36] = t[59] ^ t[60];
  assign t[37] = ~t[61];
  assign t[38] = t[62];
  assign t[39] = ~(t[21] ^ t[63]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[8] ? t[66] : t[178];
  assign t[42] = t[8] ? t[67] : t[179];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[70] & t[71];
  assign t[45] = t[8] ? t[72] : t[180];
  assign t[46] = t[73] ^ t[74];
  assign t[47] = t[75] & t[76];
  assign t[48] = ~(t[77] & t[78]);
  assign t[49] = t[181] | t[79];
  assign t[4] = t[8] ? t[9] : t[173];
  assign t[50] = ~(t[80]);
  assign t[51] = ~(t[182]);
  assign t[52] = ~(t[81] & t[174]);
  assign t[53] = t[82] ^ t[59];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[85] ^ t[41];
  assign t[56] = t[86] & t[87];
  assign t[57] = t[64] ^ t[88];
  assign t[58] = t[89] ^ t[47];
  assign t[59] = t[90] ? t[91] : t[183];
  assign t[5] = ~(t[10]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[27] ? t[94] : t[184];
  assign t[62] = t[27] ? t[95] : t[185];
  assign t[63] = t[96] ^ t[97];
  assign t[64] = t[38] ^ t[98];
  assign t[65] = t[99];
  assign t[66] = t[178] ^ t[100];
  assign t[67] = t[179] ^ t[101];
  assign t[68] = t[102] & t[103];
  assign t[69] = t[104] & t[105];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[68] ^ t[106]);
  assign t[71] = t[107] ^ t[108];
  assign t[72] = t[180] ^ t[109];
  assign t[73] = t[110] & t[111];
  assign t[74] = t[112] & t[113];
  assign t[75] = ~(t[89] ^ t[46]);
  assign t[76] = t[114] ^ t[113];
  assign t[77] = ~(t[79] & t[115]);
  assign t[78] = ~(t[186] ^ t[116]);
  assign t[79] = ~(t[117] & t[118]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[49]);
  assign t[81] = ~(t[187]);
  assign t[82] = t[90] ? t[119] : t[188];
  assign t[83] = ~(t[120]);
  assign t[84] = t[90] ? t[121] : t[189];
  assign t[85] = t[8] ? t[122] : t[190];
  assign t[86] = ~(t[55] ^ t[43]);
  assign t[87] = t[23] ^ t[105];
  assign t[88] = t[63] ^ t[123];
  assign t[89] = t[124] ^ t[125];
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[15]);
  assign t[91] = t[183] ^ t[126];
  assign t[92] = t[127] ^ t[54];
  assign t[93] = t[128] & t[129];
  assign t[94] = t[184] ^ t[130];
  assign t[95] = t[185] ^ t[131];
  assign t[96] = t[132] & t[133];
  assign t[97] = t[134] & t[65];
  assign t[98] = ~t[135];
  assign t[99] = t[27] ? t[136] : t[191];
  assign t[9] = t[173] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [116:0] x;
 output y;

 wire [361:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[137] ? x[62] : x[61];
  assign t[101] = t[137] ? x[64] : x[63];
  assign t[102] = ~(t[108]);
  assign t[103] = ~(t[85]);
  assign t[104] = ~(t[41]);
  assign t[105] = t[8] ? t[138] : t[192];
  assign t[106] = t[23] ^ t[85];
  assign t[107] = t[85] ^ t[42];
  assign t[108] = t[105] ^ t[41];
  assign t[109] = t[80] ? x[69] : x[68];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[139]);
  assign t[111] = ~(t[124]);
  assign t[112] = ~(t[125]);
  assign t[113] = t[176] ^ t[140];
  assign t[114] = t[125] ^ t[25];
  assign t[115] = ~(t[141] & t[142]);
  assign t[116] = t[143] ^ t[193];
  assign t[117] = ~(t[186]);
  assign t[118] = t[144] & t[143];
  assign t[119] = t[188] ^ t[145];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[90] ? t[146] : t[194];
  assign t[121] = t[189] ^ t[147];
  assign t[122] = t[190] ^ t[148];
  assign t[123] = t[149] & t[150];
  assign t[124] = t[8] ? t[151] : t[195];
  assign t[125] = t[175] ^ t[152];
  assign t[126] = t[153] ? x[80] : x[79];
  assign t[127] = t[154] & t[155];
  assign t[128] = ~(t[156] ^ t[92]);
  assign t[129] = t[157] ^ t[84];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[80] ? x[82] : x[81];
  assign t[131] = t[28] ? x[84] : x[83];
  assign t[132] = ~(t[158]);
  assign t[133] = ~(t[37]);
  assign t[134] = ~(t[38]);
  assign t[135] = t[27] ? t[159] : t[196];
  assign t[136] = t[191] ^ t[160];
  assign t[137] = ~(t[50]);
  assign t[138] = t[192] ^ t[161];
  assign t[139] = t[113] ^ t[125];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[8] ? t[162] : t[197];
  assign t[141] = ~(t[144] | t[143]);
  assign t[142] = ~(t[163] | t[117]);
  assign t[143] = ~(t[198]);
  assign t[144] = ~(t[193]);
  assign t[145] = t[153] ? x[95] : x[94];
  assign t[146] = t[194] ^ t[164];
  assign t[147] = t[153] ? x[97] : x[96];
  assign t[148] = t[137] ? x[99] : x[98];
  assign t[149] = ~(t[96] ^ t[165]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[166] ^ t[158];
  assign t[151] = t[195] ^ t[167];
  assign t[152] = t[27] ? t[168] : t[199];
  assign t[153] = ~(t[50]);
  assign t[154] = ~(t[169]);
  assign t[155] = ~(t[82]);
  assign t[156] = t[82] ^ t[120];
  assign t[157] = t[120] ^ t[59];
  assign t[158] = t[65] ^ t[38];
  assign t[159] = t[196] ^ t[170];
  assign t[15] = ~(t[27]);
  assign t[160] = t[137] ? x[104] : x[103];
  assign t[161] = t[137] ? x[106] : x[105];
  assign t[162] = t[197] ^ t[171];
  assign t[163] = ~(t[181]);
  assign t[164] = t[153] ? x[108] : x[107];
  assign t[165] = t[64] ^ t[37];
  assign t[166] = t[37] ^ t[98];
  assign t[167] = t[80] ? x[110] : x[109];
  assign t[168] = t[199] ^ t[172];
  assign t[169] = t[84] ^ t[120];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[80] ? x[112] : x[111];
  assign t[171] = t[28] ? x[114] : x[113];
  assign t[172] = t[28] ? x[116] : x[115];
  assign t[173] = (t[200]);
  assign t[174] = (t[201]);
  assign t[175] = (t[202]);
  assign t[176] = (t[203]);
  assign t[177] = (t[204]);
  assign t[178] = (t[205]);
  assign t[179] = (t[206]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = (t[207]);
  assign t[181] = (t[208]);
  assign t[182] = (t[209]);
  assign t[183] = (t[210]);
  assign t[184] = (t[211]);
  assign t[185] = (t[212]);
  assign t[186] = (t[213]);
  assign t[187] = (t[214]);
  assign t[188] = (t[215]);
  assign t[189] = (t[216]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[227] ^ x[4];
  assign t[201] = t[228] ^ x[9];
  assign t[202] = t[229] ^ x[12];
  assign t[203] = t[230] ^ x[15];
  assign t[204] = t[231] ^ x[18];
  assign t[205] = t[232] ^ x[21];
  assign t[206] = t[233] ^ x[24];
  assign t[207] = t[234] ^ x[27];
  assign t[208] = t[235] ^ x[30];
  assign t[209] = t[236] ^ x[33];
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = t[237] ^ x[36];
  assign t[211] = t[238] ^ x[39];
  assign t[212] = t[239] ^ x[42];
  assign t[213] = t[240] ^ x[45];
  assign t[214] = t[241] ^ x[48];
  assign t[215] = t[242] ^ x[51];
  assign t[216] = t[243] ^ x[54];
  assign t[217] = t[244] ^ x[57];
  assign t[218] = t[245] ^ x[60];
  assign t[219] = t[246] ^ x[67];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[72];
  assign t[221] = t[248] ^ x[75];
  assign t[222] = t[249] ^ x[78];
  assign t[223] = t[250] ^ x[87];
  assign t[224] = t[251] ^ x[90];
  assign t[225] = t[252] ^ x[93];
  assign t[226] = t[253] ^ x[102];
  assign t[227] = (t[254] & ~t[255]);
  assign t[228] = (t[256] & ~t[257]);
  assign t[229] = (t[258] & ~t[259]);
  assign t[22] = t[39] & t[40];
  assign t[230] = (t[260] & ~t[261]);
  assign t[231] = (t[262] & ~t[263]);
  assign t[232] = (t[264] & ~t[265]);
  assign t[233] = (t[266] & ~t[267]);
  assign t[234] = (t[268] & ~t[269]);
  assign t[235] = (t[270] & ~t[271]);
  assign t[236] = (t[272] & ~t[273]);
  assign t[237] = (t[274] & ~t[275]);
  assign t[238] = (t[276] & ~t[277]);
  assign t[239] = (t[278] & ~t[279]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (t[280] & ~t[281]);
  assign t[241] = (t[282] & ~t[283]);
  assign t[242] = (t[284] & ~t[285]);
  assign t[243] = (t[286] & ~t[287]);
  assign t[244] = (t[288] & ~t[289]);
  assign t[245] = (t[290] & ~t[291]);
  assign t[246] = (t[292] & ~t[293]);
  assign t[247] = (t[294] & ~t[295]);
  assign t[248] = (t[296] & ~t[297]);
  assign t[249] = (t[298] & ~t[299]);
  assign t[24] = t[43] ^ t[44];
  assign t[250] = (t[300] & ~t[301]);
  assign t[251] = (t[302] & ~t[303]);
  assign t[252] = (t[304] & ~t[305]);
  assign t[253] = (t[306] & ~t[307]);
  assign t[254] = t[308] ^ x[4];
  assign t[255] = t[309] ^ x[3];
  assign t[256] = t[310] ^ x[9];
  assign t[257] = t[311] ^ x[8];
  assign t[258] = t[312] ^ x[12];
  assign t[259] = t[313] ^ x[11];
  assign t[25] = t[174] ^ t[45];
  assign t[260] = t[314] ^ x[15];
  assign t[261] = t[315] ^ x[14];
  assign t[262] = t[316] ^ x[18];
  assign t[263] = t[317] ^ x[17];
  assign t[264] = t[318] ^ x[21];
  assign t[265] = t[319] ^ x[20];
  assign t[266] = t[320] ^ x[24];
  assign t[267] = t[321] ^ x[23];
  assign t[268] = t[322] ^ x[27];
  assign t[269] = t[323] ^ x[26];
  assign t[26] = t[46] ^ t[47];
  assign t[270] = t[324] ^ x[30];
  assign t[271] = t[325] ^ x[29];
  assign t[272] = t[326] ^ x[33];
  assign t[273] = t[327] ^ x[32];
  assign t[274] = t[328] ^ x[36];
  assign t[275] = t[329] ^ x[35];
  assign t[276] = t[330] ^ x[39];
  assign t[277] = t[331] ^ x[38];
  assign t[278] = t[332] ^ x[42];
  assign t[279] = t[333] ^ x[41];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[45];
  assign t[281] = t[335] ^ x[44];
  assign t[282] = t[336] ^ x[48];
  assign t[283] = t[337] ^ x[47];
  assign t[284] = t[338] ^ x[51];
  assign t[285] = t[339] ^ x[50];
  assign t[286] = t[340] ^ x[54];
  assign t[287] = t[341] ^ x[53];
  assign t[288] = t[342] ^ x[57];
  assign t[289] = t[343] ^ x[56];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[60];
  assign t[291] = t[345] ^ x[59];
  assign t[292] = t[346] ^ x[67];
  assign t[293] = t[347] ^ x[66];
  assign t[294] = t[348] ^ x[72];
  assign t[295] = t[349] ^ x[71];
  assign t[296] = t[350] ^ x[75];
  assign t[297] = t[351] ^ x[74];
  assign t[298] = t[352] ^ x[78];
  assign t[299] = t[353] ^ x[77];
  assign t[29] = ~(t[175]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[87];
  assign t[301] = t[355] ^ x[86];
  assign t[302] = t[356] ^ x[90];
  assign t[303] = t[357] ^ x[89];
  assign t[304] = t[358] ^ x[93];
  assign t[305] = t[359] ^ x[92];
  assign t[306] = t[360] ^ x[102];
  assign t[307] = t[361] ^ x[101];
  assign t[308] = (x[2]);
  assign t[309] = (x[2]);
  assign t[30] = ~(t[176]);
  assign t[310] = (x[7]);
  assign t[311] = (x[7]);
  assign t[312] = (x[10]);
  assign t[313] = (x[10]);
  assign t[314] = (x[13]);
  assign t[315] = (x[13]);
  assign t[316] = (x[16]);
  assign t[317] = (x[16]);
  assign t[318] = (x[19]);
  assign t[319] = (x[19]);
  assign t[31] = ~(t[177]);
  assign t[320] = (x[22]);
  assign t[321] = (x[22]);
  assign t[322] = (x[25]);
  assign t[323] = (x[25]);
  assign t[324] = (x[28]);
  assign t[325] = (x[28]);
  assign t[326] = (x[31]);
  assign t[327] = (x[31]);
  assign t[328] = (x[34]);
  assign t[329] = (x[34]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[37]);
  assign t[331] = (x[37]);
  assign t[332] = (x[40]);
  assign t[333] = (x[40]);
  assign t[334] = (x[43]);
  assign t[335] = (x[43]);
  assign t[336] = (x[46]);
  assign t[337] = (x[46]);
  assign t[338] = (x[49]);
  assign t[339] = (x[49]);
  assign t[33] = t[53] ^ t[54];
  assign t[340] = (x[52]);
  assign t[341] = (x[52]);
  assign t[342] = (x[55]);
  assign t[343] = (x[55]);
  assign t[344] = (x[58]);
  assign t[345] = (x[58]);
  assign t[346] = (x[65]);
  assign t[347] = (x[65]);
  assign t[348] = (x[70]);
  assign t[349] = (x[70]);
  assign t[34] = t[55] ^ t[56];
  assign t[350] = (x[73]);
  assign t[351] = (x[73]);
  assign t[352] = (x[76]);
  assign t[353] = (x[76]);
  assign t[354] = (x[85]);
  assign t[355] = (x[85]);
  assign t[356] = (x[88]);
  assign t[357] = (x[88]);
  assign t[358] = (x[91]);
  assign t[359] = (x[91]);
  assign t[35] = t[57] ^ t[58];
  assign t[360] = (x[100]);
  assign t[361] = (x[100]);
  assign t[36] = t[59] ^ t[60];
  assign t[37] = ~t[61];
  assign t[38] = t[62];
  assign t[39] = ~(t[21] ^ t[63]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[8] ? t[66] : t[178];
  assign t[42] = t[8] ? t[67] : t[179];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[70] & t[71];
  assign t[45] = t[8] ? t[72] : t[180];
  assign t[46] = t[73] ^ t[74];
  assign t[47] = t[75] & t[76];
  assign t[48] = ~(t[77] & t[78]);
  assign t[49] = t[181] | t[79];
  assign t[4] = t[8] ? t[9] : t[173];
  assign t[50] = ~(t[80]);
  assign t[51] = ~(t[182]);
  assign t[52] = ~(t[81] & t[174]);
  assign t[53] = t[82] ^ t[59];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[85] ^ t[41];
  assign t[56] = t[86] & t[87];
  assign t[57] = t[64] ^ t[88];
  assign t[58] = t[89] ^ t[47];
  assign t[59] = t[90] ? t[91] : t[183];
  assign t[5] = ~(t[10]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[27] ? t[94] : t[184];
  assign t[62] = t[27] ? t[95] : t[185];
  assign t[63] = t[96] ^ t[97];
  assign t[64] = t[38] ^ t[98];
  assign t[65] = t[99];
  assign t[66] = t[178] ^ t[100];
  assign t[67] = t[179] ^ t[101];
  assign t[68] = t[102] & t[103];
  assign t[69] = t[104] & t[105];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[68] ^ t[106]);
  assign t[71] = t[107] ^ t[108];
  assign t[72] = t[180] ^ t[109];
  assign t[73] = t[110] & t[111];
  assign t[74] = t[112] & t[113];
  assign t[75] = ~(t[89] ^ t[46]);
  assign t[76] = t[114] ^ t[113];
  assign t[77] = ~(t[79] & t[115]);
  assign t[78] = ~(t[186] ^ t[116]);
  assign t[79] = ~(t[117] & t[118]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[49]);
  assign t[81] = ~(t[187]);
  assign t[82] = t[90] ? t[119] : t[188];
  assign t[83] = ~(t[120]);
  assign t[84] = t[90] ? t[121] : t[189];
  assign t[85] = t[8] ? t[122] : t[190];
  assign t[86] = ~(t[55] ^ t[43]);
  assign t[87] = t[23] ^ t[105];
  assign t[88] = t[63] ^ t[123];
  assign t[89] = t[124] ^ t[125];
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[15]);
  assign t[91] = t[183] ^ t[126];
  assign t[92] = t[127] ^ t[54];
  assign t[93] = t[128] & t[129];
  assign t[94] = t[184] ^ t[130];
  assign t[95] = t[185] ^ t[131];
  assign t[96] = t[132] & t[133];
  assign t[97] = t[134] & t[65];
  assign t[98] = ~t[135];
  assign t[99] = t[27] ? t[136] : t[191];
  assign t[9] = t[173] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [116:0] x;
 output y;

 wire [378:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~t[132];
  assign t[101] = t[133];
  assign t[102] = ~(t[68] ^ t[134]);
  assign t[103] = t[135] ^ t[136];
  assign t[104] = t[137] & t[138];
  assign t[105] = ~(t[104] ^ t[139]);
  assign t[106] = t[19] ^ t[140];
  assign t[107] = ~(t[141] & t[142]);
  assign t[108] = t[143] ^ t[207];
  assign t[109] = ~(t[203]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[144] & t[143];
  assign t[111] = ~(t[145]);
  assign t[112] = t[111] ? x[69] : x[68];
  assign t[113] = t[100] ^ t[119];
  assign t[114] = t[146] & t[136];
  assign t[115] = t[33] ^ t[54];
  assign t[116] = t[147] & t[148];
  assign t[117] = t[124] ^ t[149];
  assign t[118] = t[150] ^ t[88];
  assign t[119] = t[151];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[134] ^ t[69];
  assign t[121] = t[205] ^ t[152];
  assign t[122] = t[27] ? t[153] : t[208];
  assign t[123] = t[154] ^ t[155];
  assign t[124] = t[85] ^ t[98];
  assign t[125] = t[204] ^ t[156];
  assign t[126] = ~(t[150] ^ t[42]);
  assign t[127] = t[23] ^ t[94];
  assign t[128] = ~(t[145]);
  assign t[129] = t[8] ? t[157] : t[209];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[206] ^ t[158];
  assign t[131] = t[159] ? t[160] : t[210];
  assign t[132] = t[27] ? t[161] : t[211];
  assign t[133] = t[27] ? t[162] : t[212];
  assign t[134] = t[163] ^ t[114];
  assign t[135] = t[101] ^ t[119];
  assign t[136] = t[164];
  assign t[137] = ~(t[140]);
  assign t[138] = ~(t[33]);
  assign t[139] = t[46] ^ t[33];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[36] ^ t[54];
  assign t[141] = ~(t[144] | t[143]);
  assign t[142] = ~(t[165] | t[109]);
  assign t[143] = ~(t[213]);
  assign t[144] = ~(t[207]);
  assign t[145] = ~(t[28]);
  assign t[146] = ~(t[101]);
  assign t[147] = ~(t[115] ^ t[70]);
  assign t[148] = t[46] ^ t[36];
  assign t[149] = t[123] ^ t[166];
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[129] ^ t[40];
  assign t[151] = t[27] ? t[167] : t[214];
  assign t[152] = t[111] ? x[92] : x[91];
  assign t[153] = t[208] ^ t[168];
  assign t[154] = t[169] & t[170];
  assign t[155] = t[171] & t[125];
  assign t[156] = t[27] ? t[172] : t[215];
  assign t[157] = t[209] ^ t[173];
  assign t[158] = t[128] ? x[97] : x[96];
  assign t[159] = ~(t[15]);
  assign t[15] = ~(t[27]);
  assign t[160] = t[210] ^ t[174];
  assign t[161] = t[211] ^ t[175];
  assign t[162] = t[212] ^ t[176];
  assign t[163] = t[177] & t[178];
  assign t[164] = t[27] ? t[179] : t[216];
  assign t[165] = ~(t[199]);
  assign t[166] = t[180] & t[181];
  assign t[167] = t[214] ^ t[182];
  assign t[168] = t[111] ? x[102] : x[101];
  assign t[169] = ~(t[183]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[84]);
  assign t[171] = ~(t[85]);
  assign t[172] = t[215] ^ t[184];
  assign t[173] = t[128] ? x[104] : x[103];
  assign t[174] = t[185] ? x[106] : x[105];
  assign t[175] = t[28] ? x[108] : x[107];
  assign t[176] = t[185] ? x[110] : x[109];
  assign t[177] = ~(t[186]);
  assign t[178] = ~(t[100]);
  assign t[179] = t[216] ^ t[187];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[154] ^ t[188]);
  assign t[181] = t[189] ^ t[183];
  assign t[182] = t[28] ? x[112] : x[111];
  assign t[183] = t[125] ^ t[85];
  assign t[184] = t[28] ? x[114] : x[113];
  assign t[185] = ~(t[145]);
  assign t[186] = t[136] ^ t[101];
  assign t[187] = t[185] ? x[116] : x[115];
  assign t[188] = t[124] ^ t[84];
  assign t[189] = t[84] ^ t[98];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] & t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = t[244] ^ x[4];
  assign t[218] = t[245] ^ x[9];
  assign t[219] = t[246] ^ x[12];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[15];
  assign t[221] = t[248] ^ x[18];
  assign t[222] = t[249] ^ x[21];
  assign t[223] = t[250] ^ x[24];
  assign t[224] = t[251] ^ x[27];
  assign t[225] = t[252] ^ x[30];
  assign t[226] = t[253] ^ x[33];
  assign t[227] = t[254] ^ x[36];
  assign t[228] = t[255] ^ x[39];
  assign t[229] = t[256] ^ x[42];
  assign t[22] = ~(t[26] ^ t[39]);
  assign t[230] = t[257] ^ x[45];
  assign t[231] = t[258] ^ x[48];
  assign t[232] = t[259] ^ x[57];
  assign t[233] = t[260] ^ x[64];
  assign t[234] = t[261] ^ x[67];
  assign t[235] = t[262] ^ x[72];
  assign t[236] = t[263] ^ x[75];
  assign t[237] = t[264] ^ x[78];
  assign t[238] = t[265] ^ x[81];
  assign t[239] = t[266] ^ x[84];
  assign t[23] = t[40] ^ t[41];
  assign t[240] = t[267] ^ x[87];
  assign t[241] = t[268] ^ x[90];
  assign t[242] = t[269] ^ x[95];
  assign t[243] = t[270] ^ x[100];
  assign t[244] = (t[271] & ~t[272]);
  assign t[245] = (t[273] & ~t[274]);
  assign t[246] = (t[275] & ~t[276]);
  assign t[247] = (t[277] & ~t[278]);
  assign t[248] = (t[279] & ~t[280]);
  assign t[249] = (t[281] & ~t[282]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[283] & ~t[284]);
  assign t[251] = (t[285] & ~t[286]);
  assign t[252] = (t[287] & ~t[288]);
  assign t[253] = (t[289] & ~t[290]);
  assign t[254] = (t[291] & ~t[292]);
  assign t[255] = (t[293] & ~t[294]);
  assign t[256] = (t[295] & ~t[296]);
  assign t[257] = (t[297] & ~t[298]);
  assign t[258] = (t[299] & ~t[300]);
  assign t[259] = (t[301] & ~t[302]);
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[260] = (t[303] & ~t[304]);
  assign t[261] = (t[305] & ~t[306]);
  assign t[262] = (t[307] & ~t[308]);
  assign t[263] = (t[309] & ~t[310]);
  assign t[264] = (t[311] & ~t[312]);
  assign t[265] = (t[313] & ~t[314]);
  assign t[266] = (t[315] & ~t[316]);
  assign t[267] = (t[317] & ~t[318]);
  assign t[268] = (t[319] & ~t[320]);
  assign t[269] = (t[321] & ~t[322]);
  assign t[26] = t[46] ^ t[47];
  assign t[270] = (t[323] & ~t[324]);
  assign t[271] = t[325] ^ x[4];
  assign t[272] = t[326] ^ x[3];
  assign t[273] = t[327] ^ x[9];
  assign t[274] = t[328] ^ x[8];
  assign t[275] = t[329] ^ x[12];
  assign t[276] = t[330] ^ x[11];
  assign t[277] = t[331] ^ x[15];
  assign t[278] = t[332] ^ x[14];
  assign t[279] = t[333] ^ x[18];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[17];
  assign t[281] = t[335] ^ x[21];
  assign t[282] = t[336] ^ x[20];
  assign t[283] = t[337] ^ x[24];
  assign t[284] = t[338] ^ x[23];
  assign t[285] = t[339] ^ x[27];
  assign t[286] = t[340] ^ x[26];
  assign t[287] = t[341] ^ x[30];
  assign t[288] = t[342] ^ x[29];
  assign t[289] = t[343] ^ x[33];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[32];
  assign t[291] = t[345] ^ x[36];
  assign t[292] = t[346] ^ x[35];
  assign t[293] = t[347] ^ x[39];
  assign t[294] = t[348] ^ x[38];
  assign t[295] = t[349] ^ x[42];
  assign t[296] = t[350] ^ x[41];
  assign t[297] = t[351] ^ x[45];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[48];
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[47];
  assign t[301] = t[355] ^ x[57];
  assign t[302] = t[356] ^ x[56];
  assign t[303] = t[357] ^ x[64];
  assign t[304] = t[358] ^ x[63];
  assign t[305] = t[359] ^ x[67];
  assign t[306] = t[360] ^ x[66];
  assign t[307] = t[361] ^ x[72];
  assign t[308] = t[362] ^ x[71];
  assign t[309] = t[363] ^ x[75];
  assign t[30] = ~(t[192]);
  assign t[310] = t[364] ^ x[74];
  assign t[311] = t[365] ^ x[78];
  assign t[312] = t[366] ^ x[77];
  assign t[313] = t[367] ^ x[81];
  assign t[314] = t[368] ^ x[80];
  assign t[315] = t[369] ^ x[84];
  assign t[316] = t[370] ^ x[83];
  assign t[317] = t[371] ^ x[87];
  assign t[318] = t[372] ^ x[86];
  assign t[319] = t[373] ^ x[90];
  assign t[31] = ~(t[193]);
  assign t[320] = t[374] ^ x[89];
  assign t[321] = t[375] ^ x[95];
  assign t[322] = t[376] ^ x[94];
  assign t[323] = t[377] ^ x[100];
  assign t[324] = t[378] ^ x[99];
  assign t[325] = (x[2]);
  assign t[326] = (x[2]);
  assign t[327] = (x[7]);
  assign t[328] = (x[7]);
  assign t[329] = (x[10]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[10]);
  assign t[331] = (x[13]);
  assign t[332] = (x[13]);
  assign t[333] = (x[16]);
  assign t[334] = (x[16]);
  assign t[335] = (x[19]);
  assign t[336] = (x[19]);
  assign t[337] = (x[22]);
  assign t[338] = (x[22]);
  assign t[339] = (x[25]);
  assign t[33] = t[8] ? t[52] : t[194];
  assign t[340] = (x[25]);
  assign t[341] = (x[28]);
  assign t[342] = (x[28]);
  assign t[343] = (x[31]);
  assign t[344] = (x[31]);
  assign t[345] = (x[34]);
  assign t[346] = (x[34]);
  assign t[347] = (x[37]);
  assign t[348] = (x[37]);
  assign t[349] = (x[40]);
  assign t[34] = t[8] ? t[53] : t[195];
  assign t[350] = (x[40]);
  assign t[351] = (x[43]);
  assign t[352] = (x[43]);
  assign t[353] = (x[46]);
  assign t[354] = (x[46]);
  assign t[355] = (x[55]);
  assign t[356] = (x[55]);
  assign t[357] = (x[62]);
  assign t[358] = (x[62]);
  assign t[359] = (x[65]);
  assign t[35] = ~(t[54]);
  assign t[360] = (x[65]);
  assign t[361] = (x[70]);
  assign t[362] = (x[70]);
  assign t[363] = (x[73]);
  assign t[364] = (x[73]);
  assign t[365] = (x[76]);
  assign t[366] = (x[76]);
  assign t[367] = (x[79]);
  assign t[368] = (x[79]);
  assign t[369] = (x[82]);
  assign t[36] = t[8] ? t[55] : t[196];
  assign t[370] = (x[82]);
  assign t[371] = (x[85]);
  assign t[372] = (x[85]);
  assign t[373] = (x[88]);
  assign t[374] = (x[88]);
  assign t[375] = (x[93]);
  assign t[376] = (x[93]);
  assign t[377] = (x[98]);
  assign t[378] = (x[98]);
  assign t[37] = ~(t[56] ^ t[57]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[41] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[61] : t[197];
  assign t[41] = t[8] ? t[62] : t[198];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[65] & t[66];
  assign t[44] = t[13] ^ t[67];
  assign t[45] = t[68] ^ t[69];
  assign t[46] = t[54] ^ t[34];
  assign t[47] = t[70] ^ t[71];
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = t[199] | t[74];
  assign t[4] = t[8] ? t[9] : t[190];
  assign t[50] = ~(t[200]);
  assign t[51] = ~(t[75] & t[201]);
  assign t[52] = t[194] ^ t[76];
  assign t[53] = t[195] ^ t[77];
  assign t[54] = t[8] ? t[78] : t[202];
  assign t[55] = t[196] ^ t[79];
  assign t[56] = t[80] ^ t[81];
  assign t[57] = ~(t[82] ^ t[83]);
  assign t[58] = t[84] ^ t[85];
  assign t[59] = t[86] & t[87];
  assign t[5] = ~(t[10]);
  assign t[60] = t[42] ^ t[88];
  assign t[61] = t[197] ^ t[89];
  assign t[62] = t[198] ^ t[90];
  assign t[63] = t[91] & t[92];
  assign t[64] = t[93] & t[94];
  assign t[65] = ~(t[63] ^ t[95]);
  assign t[66] = t[96] ^ t[97];
  assign t[67] = t[98] ^ t[99];
  assign t[68] = t[100] ^ t[101];
  assign t[69] = t[102] & t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[104] ^ t[20];
  assign t[71] = t[105] & t[106];
  assign t[72] = ~(t[74] & t[107]);
  assign t[73] = ~(t[203] ^ t[108]);
  assign t[74] = ~(t[109] & t[110]);
  assign t[75] = ~(t[204]);
  assign t[76] = t[111] ? x[50] : x[49];
  assign t[77] = t[111] ? x[52] : x[51];
  assign t[78] = t[202] ^ t[112];
  assign t[79] = t[111] ? x[54] : x[53];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[113] ^ t[114];
  assign t[81] = t[115] ^ t[116];
  assign t[82] = t[117] ^ t[118];
  assign t[83] = t[119] ^ t[120];
  assign t[84] = t[27] ? t[121] : t[205];
  assign t[85] = t[193] ^ t[122];
  assign t[86] = ~(t[58] ^ t[123]);
  assign t[87] = t[124] ^ t[125];
  assign t[88] = t[126] & t[127];
  assign t[89] = t[128] ? x[59] : x[58];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] ? x[61] : x[60];
  assign t[91] = ~(t[97]);
  assign t[92] = ~(t[129]);
  assign t[93] = ~(t[40]);
  assign t[94] = t[8] ? t[130] : t[206];
  assign t[95] = t[23] ^ t[129];
  assign t[96] = t[129] ^ t[41];
  assign t[97] = t[94] ^ t[40];
  assign t[98] = t[200] ^ t[131];
  assign t[99] = t[123] ^ t[59];
  assign t[9] = t[190] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [116:0] x;
 output y;

 wire [378:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~t[132];
  assign t[101] = t[133];
  assign t[102] = ~(t[68] ^ t[134]);
  assign t[103] = t[135] ^ t[136];
  assign t[104] = t[137] & t[138];
  assign t[105] = ~(t[104] ^ t[139]);
  assign t[106] = t[19] ^ t[140];
  assign t[107] = ~(t[141] & t[142]);
  assign t[108] = t[143] ^ t[207];
  assign t[109] = ~(t[203]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[144] & t[143];
  assign t[111] = ~(t[145]);
  assign t[112] = t[111] ? x[69] : x[68];
  assign t[113] = t[100] ^ t[119];
  assign t[114] = t[146] & t[136];
  assign t[115] = t[33] ^ t[54];
  assign t[116] = t[147] & t[148];
  assign t[117] = t[124] ^ t[149];
  assign t[118] = t[150] ^ t[88];
  assign t[119] = t[151];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[134] ^ t[69];
  assign t[121] = t[205] ^ t[152];
  assign t[122] = t[27] ? t[153] : t[208];
  assign t[123] = t[154] ^ t[155];
  assign t[124] = t[85] ^ t[98];
  assign t[125] = t[204] ^ t[156];
  assign t[126] = ~(t[150] ^ t[42]);
  assign t[127] = t[23] ^ t[94];
  assign t[128] = ~(t[145]);
  assign t[129] = t[8] ? t[157] : t[209];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[206] ^ t[158];
  assign t[131] = t[159] ? t[160] : t[210];
  assign t[132] = t[27] ? t[161] : t[211];
  assign t[133] = t[27] ? t[162] : t[212];
  assign t[134] = t[163] ^ t[114];
  assign t[135] = t[101] ^ t[119];
  assign t[136] = t[164];
  assign t[137] = ~(t[140]);
  assign t[138] = ~(t[33]);
  assign t[139] = t[46] ^ t[33];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[36] ^ t[54];
  assign t[141] = ~(t[144] | t[143]);
  assign t[142] = ~(t[165] | t[109]);
  assign t[143] = ~(t[213]);
  assign t[144] = ~(t[207]);
  assign t[145] = ~(t[28]);
  assign t[146] = ~(t[101]);
  assign t[147] = ~(t[115] ^ t[70]);
  assign t[148] = t[46] ^ t[36];
  assign t[149] = t[123] ^ t[166];
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[129] ^ t[40];
  assign t[151] = t[27] ? t[167] : t[214];
  assign t[152] = t[111] ? x[92] : x[91];
  assign t[153] = t[208] ^ t[168];
  assign t[154] = t[169] & t[170];
  assign t[155] = t[171] & t[125];
  assign t[156] = t[27] ? t[172] : t[215];
  assign t[157] = t[209] ^ t[173];
  assign t[158] = t[128] ? x[97] : x[96];
  assign t[159] = ~(t[15]);
  assign t[15] = ~(t[27]);
  assign t[160] = t[210] ^ t[174];
  assign t[161] = t[211] ^ t[175];
  assign t[162] = t[212] ^ t[176];
  assign t[163] = t[177] & t[178];
  assign t[164] = t[27] ? t[179] : t[216];
  assign t[165] = ~(t[199]);
  assign t[166] = t[180] & t[181];
  assign t[167] = t[214] ^ t[182];
  assign t[168] = t[111] ? x[102] : x[101];
  assign t[169] = ~(t[183]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[84]);
  assign t[171] = ~(t[85]);
  assign t[172] = t[215] ^ t[184];
  assign t[173] = t[128] ? x[104] : x[103];
  assign t[174] = t[185] ? x[106] : x[105];
  assign t[175] = t[28] ? x[108] : x[107];
  assign t[176] = t[185] ? x[110] : x[109];
  assign t[177] = ~(t[186]);
  assign t[178] = ~(t[100]);
  assign t[179] = t[216] ^ t[187];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[154] ^ t[188]);
  assign t[181] = t[189] ^ t[183];
  assign t[182] = t[28] ? x[112] : x[111];
  assign t[183] = t[125] ^ t[85];
  assign t[184] = t[28] ? x[114] : x[113];
  assign t[185] = ~(t[145]);
  assign t[186] = t[136] ^ t[101];
  assign t[187] = t[185] ? x[116] : x[115];
  assign t[188] = t[124] ^ t[84];
  assign t[189] = t[84] ^ t[98];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] & t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = t[244] ^ x[4];
  assign t[218] = t[245] ^ x[9];
  assign t[219] = t[246] ^ x[12];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[15];
  assign t[221] = t[248] ^ x[18];
  assign t[222] = t[249] ^ x[21];
  assign t[223] = t[250] ^ x[24];
  assign t[224] = t[251] ^ x[27];
  assign t[225] = t[252] ^ x[30];
  assign t[226] = t[253] ^ x[33];
  assign t[227] = t[254] ^ x[36];
  assign t[228] = t[255] ^ x[39];
  assign t[229] = t[256] ^ x[42];
  assign t[22] = ~(t[26] ^ t[39]);
  assign t[230] = t[257] ^ x[45];
  assign t[231] = t[258] ^ x[48];
  assign t[232] = t[259] ^ x[57];
  assign t[233] = t[260] ^ x[64];
  assign t[234] = t[261] ^ x[67];
  assign t[235] = t[262] ^ x[72];
  assign t[236] = t[263] ^ x[75];
  assign t[237] = t[264] ^ x[78];
  assign t[238] = t[265] ^ x[81];
  assign t[239] = t[266] ^ x[84];
  assign t[23] = t[40] ^ t[41];
  assign t[240] = t[267] ^ x[87];
  assign t[241] = t[268] ^ x[90];
  assign t[242] = t[269] ^ x[95];
  assign t[243] = t[270] ^ x[100];
  assign t[244] = (t[271] & ~t[272]);
  assign t[245] = (t[273] & ~t[274]);
  assign t[246] = (t[275] & ~t[276]);
  assign t[247] = (t[277] & ~t[278]);
  assign t[248] = (t[279] & ~t[280]);
  assign t[249] = (t[281] & ~t[282]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[283] & ~t[284]);
  assign t[251] = (t[285] & ~t[286]);
  assign t[252] = (t[287] & ~t[288]);
  assign t[253] = (t[289] & ~t[290]);
  assign t[254] = (t[291] & ~t[292]);
  assign t[255] = (t[293] & ~t[294]);
  assign t[256] = (t[295] & ~t[296]);
  assign t[257] = (t[297] & ~t[298]);
  assign t[258] = (t[299] & ~t[300]);
  assign t[259] = (t[301] & ~t[302]);
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[260] = (t[303] & ~t[304]);
  assign t[261] = (t[305] & ~t[306]);
  assign t[262] = (t[307] & ~t[308]);
  assign t[263] = (t[309] & ~t[310]);
  assign t[264] = (t[311] & ~t[312]);
  assign t[265] = (t[313] & ~t[314]);
  assign t[266] = (t[315] & ~t[316]);
  assign t[267] = (t[317] & ~t[318]);
  assign t[268] = (t[319] & ~t[320]);
  assign t[269] = (t[321] & ~t[322]);
  assign t[26] = t[46] ^ t[47];
  assign t[270] = (t[323] & ~t[324]);
  assign t[271] = t[325] ^ x[4];
  assign t[272] = t[326] ^ x[3];
  assign t[273] = t[327] ^ x[9];
  assign t[274] = t[328] ^ x[8];
  assign t[275] = t[329] ^ x[12];
  assign t[276] = t[330] ^ x[11];
  assign t[277] = t[331] ^ x[15];
  assign t[278] = t[332] ^ x[14];
  assign t[279] = t[333] ^ x[18];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[17];
  assign t[281] = t[335] ^ x[21];
  assign t[282] = t[336] ^ x[20];
  assign t[283] = t[337] ^ x[24];
  assign t[284] = t[338] ^ x[23];
  assign t[285] = t[339] ^ x[27];
  assign t[286] = t[340] ^ x[26];
  assign t[287] = t[341] ^ x[30];
  assign t[288] = t[342] ^ x[29];
  assign t[289] = t[343] ^ x[33];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[32];
  assign t[291] = t[345] ^ x[36];
  assign t[292] = t[346] ^ x[35];
  assign t[293] = t[347] ^ x[39];
  assign t[294] = t[348] ^ x[38];
  assign t[295] = t[349] ^ x[42];
  assign t[296] = t[350] ^ x[41];
  assign t[297] = t[351] ^ x[45];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[48];
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[47];
  assign t[301] = t[355] ^ x[57];
  assign t[302] = t[356] ^ x[56];
  assign t[303] = t[357] ^ x[64];
  assign t[304] = t[358] ^ x[63];
  assign t[305] = t[359] ^ x[67];
  assign t[306] = t[360] ^ x[66];
  assign t[307] = t[361] ^ x[72];
  assign t[308] = t[362] ^ x[71];
  assign t[309] = t[363] ^ x[75];
  assign t[30] = ~(t[192]);
  assign t[310] = t[364] ^ x[74];
  assign t[311] = t[365] ^ x[78];
  assign t[312] = t[366] ^ x[77];
  assign t[313] = t[367] ^ x[81];
  assign t[314] = t[368] ^ x[80];
  assign t[315] = t[369] ^ x[84];
  assign t[316] = t[370] ^ x[83];
  assign t[317] = t[371] ^ x[87];
  assign t[318] = t[372] ^ x[86];
  assign t[319] = t[373] ^ x[90];
  assign t[31] = ~(t[193]);
  assign t[320] = t[374] ^ x[89];
  assign t[321] = t[375] ^ x[95];
  assign t[322] = t[376] ^ x[94];
  assign t[323] = t[377] ^ x[100];
  assign t[324] = t[378] ^ x[99];
  assign t[325] = (x[2]);
  assign t[326] = (x[2]);
  assign t[327] = (x[7]);
  assign t[328] = (x[7]);
  assign t[329] = (x[10]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[10]);
  assign t[331] = (x[13]);
  assign t[332] = (x[13]);
  assign t[333] = (x[16]);
  assign t[334] = (x[16]);
  assign t[335] = (x[19]);
  assign t[336] = (x[19]);
  assign t[337] = (x[22]);
  assign t[338] = (x[22]);
  assign t[339] = (x[25]);
  assign t[33] = t[8] ? t[52] : t[194];
  assign t[340] = (x[25]);
  assign t[341] = (x[28]);
  assign t[342] = (x[28]);
  assign t[343] = (x[31]);
  assign t[344] = (x[31]);
  assign t[345] = (x[34]);
  assign t[346] = (x[34]);
  assign t[347] = (x[37]);
  assign t[348] = (x[37]);
  assign t[349] = (x[40]);
  assign t[34] = t[8] ? t[53] : t[195];
  assign t[350] = (x[40]);
  assign t[351] = (x[43]);
  assign t[352] = (x[43]);
  assign t[353] = (x[46]);
  assign t[354] = (x[46]);
  assign t[355] = (x[55]);
  assign t[356] = (x[55]);
  assign t[357] = (x[62]);
  assign t[358] = (x[62]);
  assign t[359] = (x[65]);
  assign t[35] = ~(t[54]);
  assign t[360] = (x[65]);
  assign t[361] = (x[70]);
  assign t[362] = (x[70]);
  assign t[363] = (x[73]);
  assign t[364] = (x[73]);
  assign t[365] = (x[76]);
  assign t[366] = (x[76]);
  assign t[367] = (x[79]);
  assign t[368] = (x[79]);
  assign t[369] = (x[82]);
  assign t[36] = t[8] ? t[55] : t[196];
  assign t[370] = (x[82]);
  assign t[371] = (x[85]);
  assign t[372] = (x[85]);
  assign t[373] = (x[88]);
  assign t[374] = (x[88]);
  assign t[375] = (x[93]);
  assign t[376] = (x[93]);
  assign t[377] = (x[98]);
  assign t[378] = (x[98]);
  assign t[37] = ~(t[56] ^ t[57]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[41] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[61] : t[197];
  assign t[41] = t[8] ? t[62] : t[198];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[65] & t[66];
  assign t[44] = t[13] ^ t[67];
  assign t[45] = t[68] ^ t[69];
  assign t[46] = t[54] ^ t[34];
  assign t[47] = t[70] ^ t[71];
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = t[199] | t[74];
  assign t[4] = t[8] ? t[9] : t[190];
  assign t[50] = ~(t[200]);
  assign t[51] = ~(t[75] & t[201]);
  assign t[52] = t[194] ^ t[76];
  assign t[53] = t[195] ^ t[77];
  assign t[54] = t[8] ? t[78] : t[202];
  assign t[55] = t[196] ^ t[79];
  assign t[56] = t[80] ^ t[81];
  assign t[57] = ~(t[82] ^ t[83]);
  assign t[58] = t[84] ^ t[85];
  assign t[59] = t[86] & t[87];
  assign t[5] = ~(t[10]);
  assign t[60] = t[42] ^ t[88];
  assign t[61] = t[197] ^ t[89];
  assign t[62] = t[198] ^ t[90];
  assign t[63] = t[91] & t[92];
  assign t[64] = t[93] & t[94];
  assign t[65] = ~(t[63] ^ t[95]);
  assign t[66] = t[96] ^ t[97];
  assign t[67] = t[98] ^ t[99];
  assign t[68] = t[100] ^ t[101];
  assign t[69] = t[102] & t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[104] ^ t[20];
  assign t[71] = t[105] & t[106];
  assign t[72] = ~(t[74] & t[107]);
  assign t[73] = ~(t[203] ^ t[108]);
  assign t[74] = ~(t[109] & t[110]);
  assign t[75] = ~(t[204]);
  assign t[76] = t[111] ? x[50] : x[49];
  assign t[77] = t[111] ? x[52] : x[51];
  assign t[78] = t[202] ^ t[112];
  assign t[79] = t[111] ? x[54] : x[53];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[113] ^ t[114];
  assign t[81] = t[115] ^ t[116];
  assign t[82] = t[117] ^ t[118];
  assign t[83] = t[119] ^ t[120];
  assign t[84] = t[27] ? t[121] : t[205];
  assign t[85] = t[193] ^ t[122];
  assign t[86] = ~(t[58] ^ t[123]);
  assign t[87] = t[124] ^ t[125];
  assign t[88] = t[126] & t[127];
  assign t[89] = t[128] ? x[59] : x[58];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] ? x[61] : x[60];
  assign t[91] = ~(t[97]);
  assign t[92] = ~(t[129]);
  assign t[93] = ~(t[40]);
  assign t[94] = t[8] ? t[130] : t[206];
  assign t[95] = t[23] ^ t[129];
  assign t[96] = t[129] ^ t[41];
  assign t[97] = t[94] ^ t[40];
  assign t[98] = t[200] ^ t[131];
  assign t[99] = t[123] ^ t[59];
  assign t[9] = t[190] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [116:0] x;
 output y;

 wire [396:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[214] ^ t[137];
  assign t[101] = t[138] ^ t[121];
  assign t[102] = t[139] & t[140];
  assign t[103] = t[219] ^ t[141];
  assign t[104] = t[142] ^ t[143];
  assign t[105] = t[42] ^ t[144];
  assign t[106] = t[145] ^ t[146];
  assign t[107] = t[27] ? t[147] : t[225];
  assign t[108] = ~(t[72] ^ t[101]);
  assign t[109] = t[66] ^ t[148];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[149] & t[150];
  assign t[111] = ~(t[151] & t[152]);
  assign t[112] = t[153] ^ t[226];
  assign t[113] = ~(t[220]);
  assign t[114] = t[154] & t[153];
  assign t[115] = t[100] ^ t[155];
  assign t[116] = t[156] ^ t[157];
  assign t[117] = t[158] & t[159];
  assign t[118] = t[157] ^ t[145];
  assign t[119] = t[160] ^ t[161];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[107] ^ t[100];
  assign t[121] = t[162] & t[148];
  assign t[122] = t[28] ? x[64] : x[63];
  assign t[123] = t[28] ? x[66] : x[65];
  assign t[124] = t[163] & t[164];
  assign t[125] = t[165] & t[88];
  assign t[126] = t[222] ^ t[166];
  assign t[127] = t[132] ? x[68] : x[67];
  assign t[128] = ~(t[131]);
  assign t[129] = ~(t[96]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[37] ^ t[96];
  assign t[131] = t[98] ^ t[59];
  assign t[132] = ~(t[49]);
  assign t[133] = t[96] ^ t[59];
  assign t[134] = t[223] ^ t[167];
  assign t[135] = t[224] ^ t[168];
  assign t[136] = t[27] ? t[169] : t[227];
  assign t[137] = t[170] ? t[171] : t[228];
  assign t[138] = t[172] & t[173];
  assign t[139] = ~(t[138] ^ t[174]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[120] ^ t[175];
  assign t[141] = t[28] ? x[76] : x[75];
  assign t[142] = t[156] ^ t[145];
  assign t[143] = t[176] & t[177];
  assign t[144] = t[133] ^ t[63];
  assign t[145] = t[178];
  assign t[146] = t[160] ^ t[117];
  assign t[147] = t[225] ^ t[179];
  assign t[148] = t[221] ^ t[180];
  assign t[149] = ~(t[124] ^ t[181]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[182] ^ t[183];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[184] | t[113]);
  assign t[153] = ~(t[229]);
  assign t[154] = ~(t[226]);
  assign t[155] = t[101] ^ t[73];
  assign t[156] = ~t[185];
  assign t[157] = t[186];
  assign t[158] = ~(t[116] ^ t[160]);
  assign t[159] = t[118] ^ t[177];
  assign t[15] = ~(t[27]);
  assign t[160] = t[187] ^ t[143];
  assign t[161] = t[188] & t[189];
  assign t[162] = ~(t[99]);
  assign t[163] = ~(t[183]);
  assign t[164] = ~(t[55]);
  assign t[165] = ~(t[56]);
  assign t[166] = t[28] ? x[81] : x[80];
  assign t[167] = t[132] ? x[83] : x[82];
  assign t[168] = t[132] ? x[85] : x[84];
  assign t[169] = t[227] ^ t[190];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[15]);
  assign t[171] = t[228] ^ t[191];
  assign t[172] = ~(t[175]);
  assign t[173] = ~(t[107]);
  assign t[174] = t[66] ^ t[107];
  assign t[175] = t[148] ^ t[99];
  assign t[176] = ~(t[157]);
  assign t[177] = t[192];
  assign t[178] = t[27] ? t[193] : t[230];
  assign t[179] = t[28] ? x[90] : x[89];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[27] ? t[194] : t[231];
  assign t[181] = t[74] ^ t[55];
  assign t[182] = t[55] ^ t[68];
  assign t[183] = t[88] ^ t[56];
  assign t[184] = ~(t[213]);
  assign t[185] = t[27] ? t[195] : t[232];
  assign t[186] = t[27] ? t[196] : t[233];
  assign t[187] = t[197] & t[198];
  assign t[188] = ~(t[187] ^ t[199]);
  assign t[189] = t[142] ^ t[200];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[28] ? x[101] : x[100];
  assign t[191] = t[201] ? x[103] : x[102];
  assign t[192] = t[27] ? t[202] : t[234];
  assign t[193] = t[230] ^ t[203];
  assign t[194] = t[231] ^ t[204];
  assign t[195] = t[232] ^ t[205];
  assign t[196] = t[233] ^ t[206];
  assign t[197] = ~(t[200]);
  assign t[198] = ~(t[156]);
  assign t[199] = t[118] ^ t[156];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[177] ^ t[157];
  assign t[201] = ~(t[49]);
  assign t[202] = t[234] ^ t[207];
  assign t[203] = t[79] ? x[108] : x[107];
  assign t[204] = t[79] ? x[110] : x[109];
  assign t[205] = t[79] ? x[112] : x[111];
  assign t[206] = t[201] ? x[114] : x[113];
  assign t[207] = t[201] ? x[116] : x[115];
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = t[262] ^ x[4];
  assign t[236] = t[263] ^ x[9];
  assign t[237] = t[264] ^ x[12];
  assign t[238] = t[265] ^ x[15];
  assign t[239] = t[266] ^ x[18];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[21];
  assign t[241] = t[268] ^ x[24];
  assign t[242] = t[269] ^ x[27];
  assign t[243] = t[270] ^ x[30];
  assign t[244] = t[271] ^ x[33];
  assign t[245] = t[272] ^ x[36];
  assign t[246] = t[273] ^ x[39];
  assign t[247] = t[274] ^ x[42];
  assign t[248] = t[275] ^ x[45];
  assign t[249] = t[276] ^ x[48];
  assign t[24] = ~(t[33] ^ t[43]);
  assign t[250] = t[277] ^ x[53];
  assign t[251] = t[278] ^ x[56];
  assign t[252] = t[279] ^ x[59];
  assign t[253] = t[280] ^ x[62];
  assign t[254] = t[281] ^ x[71];
  assign t[255] = t[282] ^ x[74];
  assign t[256] = t[283] ^ x[79];
  assign t[257] = t[284] ^ x[88];
  assign t[258] = t[285] ^ x[93];
  assign t[259] = t[286] ^ x[96];
  assign t[25] = t[44] ^ t[45];
  assign t[260] = t[287] ^ x[99];
  assign t[261] = t[288] ^ x[106];
  assign t[262] = (t[289] & ~t[290]);
  assign t[263] = (t[291] & ~t[292]);
  assign t[264] = (t[293] & ~t[294]);
  assign t[265] = (t[295] & ~t[296]);
  assign t[266] = (t[297] & ~t[298]);
  assign t[267] = (t[299] & ~t[300]);
  assign t[268] = (t[301] & ~t[302]);
  assign t[269] = (t[303] & ~t[304]);
  assign t[26] = ~(t[46] ^ t[22]);
  assign t[270] = (t[305] & ~t[306]);
  assign t[271] = (t[307] & ~t[308]);
  assign t[272] = (t[309] & ~t[310]);
  assign t[273] = (t[311] & ~t[312]);
  assign t[274] = (t[313] & ~t[314]);
  assign t[275] = (t[315] & ~t[316]);
  assign t[276] = (t[317] & ~t[318]);
  assign t[277] = (t[319] & ~t[320]);
  assign t[278] = (t[321] & ~t[322]);
  assign t[279] = (t[323] & ~t[324]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[325] & ~t[326]);
  assign t[281] = (t[327] & ~t[328]);
  assign t[282] = (t[329] & ~t[330]);
  assign t[283] = (t[331] & ~t[332]);
  assign t[284] = (t[333] & ~t[334]);
  assign t[285] = (t[335] & ~t[336]);
  assign t[286] = (t[337] & ~t[338]);
  assign t[287] = (t[339] & ~t[340]);
  assign t[288] = (t[341] & ~t[342]);
  assign t[289] = t[343] ^ x[4];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[3];
  assign t[291] = t[345] ^ x[9];
  assign t[292] = t[346] ^ x[8];
  assign t[293] = t[347] ^ x[12];
  assign t[294] = t[348] ^ x[11];
  assign t[295] = t[349] ^ x[15];
  assign t[296] = t[350] ^ x[14];
  assign t[297] = t[351] ^ x[18];
  assign t[298] = t[352] ^ x[17];
  assign t[299] = t[353] ^ x[21];
  assign t[29] = ~(t[209]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[20];
  assign t[301] = t[355] ^ x[24];
  assign t[302] = t[356] ^ x[23];
  assign t[303] = t[357] ^ x[27];
  assign t[304] = t[358] ^ x[26];
  assign t[305] = t[359] ^ x[30];
  assign t[306] = t[360] ^ x[29];
  assign t[307] = t[361] ^ x[33];
  assign t[308] = t[362] ^ x[32];
  assign t[309] = t[363] ^ x[36];
  assign t[30] = ~(t[210]);
  assign t[310] = t[364] ^ x[35];
  assign t[311] = t[365] ^ x[39];
  assign t[312] = t[366] ^ x[38];
  assign t[313] = t[367] ^ x[42];
  assign t[314] = t[368] ^ x[41];
  assign t[315] = t[369] ^ x[45];
  assign t[316] = t[370] ^ x[44];
  assign t[317] = t[371] ^ x[48];
  assign t[318] = t[372] ^ x[47];
  assign t[319] = t[373] ^ x[53];
  assign t[31] = ~(t[211]);
  assign t[320] = t[374] ^ x[52];
  assign t[321] = t[375] ^ x[56];
  assign t[322] = t[376] ^ x[55];
  assign t[323] = t[377] ^ x[59];
  assign t[324] = t[378] ^ x[58];
  assign t[325] = t[379] ^ x[62];
  assign t[326] = t[380] ^ x[61];
  assign t[327] = t[381] ^ x[71];
  assign t[328] = t[382] ^ x[70];
  assign t[329] = t[383] ^ x[74];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[73];
  assign t[331] = t[385] ^ x[79];
  assign t[332] = t[386] ^ x[78];
  assign t[333] = t[387] ^ x[88];
  assign t[334] = t[388] ^ x[87];
  assign t[335] = t[389] ^ x[93];
  assign t[336] = t[390] ^ x[92];
  assign t[337] = t[391] ^ x[96];
  assign t[338] = t[392] ^ x[95];
  assign t[339] = t[393] ^ x[99];
  assign t[33] = ~(t[52] ^ t[46]);
  assign t[340] = t[394] ^ x[98];
  assign t[341] = t[395] ^ x[106];
  assign t[342] = t[396] ^ x[105];
  assign t[343] = (x[2]);
  assign t[344] = (x[2]);
  assign t[345] = (x[7]);
  assign t[346] = (x[7]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[51]);
  assign t[374] = (x[51]);
  assign t[375] = (x[54]);
  assign t[376] = (x[54]);
  assign t[377] = (x[57]);
  assign t[378] = (x[57]);
  assign t[379] = (x[60]);
  assign t[37] = t[59] ^ t[39];
  assign t[380] = (x[60]);
  assign t[381] = (x[69]);
  assign t[382] = (x[69]);
  assign t[383] = (x[72]);
  assign t[384] = (x[72]);
  assign t[385] = (x[77]);
  assign t[386] = (x[77]);
  assign t[387] = (x[86]);
  assign t[388] = (x[86]);
  assign t[389] = (x[91]);
  assign t[38] = t[60] ^ t[61];
  assign t[390] = (x[91]);
  assign t[391] = (x[94]);
  assign t[392] = (x[94]);
  assign t[393] = (x[97]);
  assign t[394] = (x[97]);
  assign t[395] = (x[104]);
  assign t[396] = (x[104]);
  assign t[39] = t[8] ? t[62] : t[212];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[60] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = ~(t[70] ^ t[71]);
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = t[213] | t[78];
  assign t[49] = ~(t[79]);
  assign t[4] = t[8] ? t[9] : t[208];
  assign t[50] = ~(t[214]);
  assign t[51] = ~(t[80] & t[215]);
  assign t[52] = ~(t[81] ^ t[82]);
  assign t[53] = t[83] ^ t[84];
  assign t[54] = ~(t[43] ^ t[22]);
  assign t[55] = t[8] ? t[85] : t[216];
  assign t[56] = t[8] ? t[86] : t[217];
  assign t[57] = ~(t[35] ^ t[87]);
  assign t[58] = t[74] ^ t[88];
  assign t[59] = t[8] ? t[89] : t[218];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[65];
  assign t[61] = t[91] & t[92];
  assign t[62] = t[212] ^ t[93];
  assign t[63] = t[94] & t[95];
  assign t[64] = t[96] ^ t[39];
  assign t[65] = t[97] & t[98];
  assign t[66] = t[99] ^ t[100];
  assign t[67] = t[101] ^ t[102];
  assign t[68] = t[8] ? t[103] : t[219];
  assign t[69] = t[87] ^ t[36];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[104] ^ t[20];
  assign t[71] = ~(t[105] ^ t[106]);
  assign t[72] = t[107] ^ t[99];
  assign t[73] = t[108] & t[109];
  assign t[74] = t[56] ^ t[68];
  assign t[75] = t[87] ^ t[110];
  assign t[76] = ~(t[78] & t[111]);
  assign t[77] = ~(t[220] ^ t[112]);
  assign t[78] = ~(t[113] & t[114]);
  assign t[79] = ~(t[48]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[221]);
  assign t[81] = t[21] ^ t[115];
  assign t[82] = t[116] ^ t[117];
  assign t[83] = t[118] ^ t[119];
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[216] ^ t[122];
  assign t[86] = t[217] ^ t[123];
  assign t[87] = t[124] ^ t[125];
  assign t[88] = t[8] ? t[126] : t[222];
  assign t[89] = t[218] ^ t[127];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] & t[129];
  assign t[91] = ~(t[90] ^ t[130]);
  assign t[92] = t[64] ^ t[131];
  assign t[93] = t[132] ? x[50] : x[49];
  assign t[94] = ~(t[133] ^ t[60]);
  assign t[95] = t[37] ^ t[98];
  assign t[96] = t[8] ? t[134] : t[223];
  assign t[97] = ~(t[59]);
  assign t[98] = t[8] ? t[135] : t[224];
  assign t[99] = t[211] ^ t[136];
  assign t[9] = t[208] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind91(x, y);
 input [116:0] x;
 output y;

 wire [396:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[214] ^ t[137];
  assign t[101] = t[138] ^ t[121];
  assign t[102] = t[139] & t[140];
  assign t[103] = t[219] ^ t[141];
  assign t[104] = t[142] ^ t[143];
  assign t[105] = t[42] ^ t[144];
  assign t[106] = t[145] ^ t[146];
  assign t[107] = t[27] ? t[147] : t[225];
  assign t[108] = ~(t[72] ^ t[101]);
  assign t[109] = t[66] ^ t[148];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[149] & t[150];
  assign t[111] = ~(t[151] & t[152]);
  assign t[112] = t[153] ^ t[226];
  assign t[113] = ~(t[220]);
  assign t[114] = t[154] & t[153];
  assign t[115] = t[100] ^ t[155];
  assign t[116] = t[156] ^ t[157];
  assign t[117] = t[158] & t[159];
  assign t[118] = t[157] ^ t[145];
  assign t[119] = t[160] ^ t[161];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[107] ^ t[100];
  assign t[121] = t[162] & t[148];
  assign t[122] = t[28] ? x[64] : x[63];
  assign t[123] = t[28] ? x[66] : x[65];
  assign t[124] = t[163] & t[164];
  assign t[125] = t[165] & t[88];
  assign t[126] = t[222] ^ t[166];
  assign t[127] = t[132] ? x[68] : x[67];
  assign t[128] = ~(t[131]);
  assign t[129] = ~(t[96]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[37] ^ t[96];
  assign t[131] = t[98] ^ t[59];
  assign t[132] = ~(t[49]);
  assign t[133] = t[96] ^ t[59];
  assign t[134] = t[223] ^ t[167];
  assign t[135] = t[224] ^ t[168];
  assign t[136] = t[27] ? t[169] : t[227];
  assign t[137] = t[170] ? t[171] : t[228];
  assign t[138] = t[172] & t[173];
  assign t[139] = ~(t[138] ^ t[174]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[120] ^ t[175];
  assign t[141] = t[28] ? x[76] : x[75];
  assign t[142] = t[156] ^ t[145];
  assign t[143] = t[176] & t[177];
  assign t[144] = t[133] ^ t[63];
  assign t[145] = t[178];
  assign t[146] = t[160] ^ t[117];
  assign t[147] = t[225] ^ t[179];
  assign t[148] = t[221] ^ t[180];
  assign t[149] = ~(t[124] ^ t[181]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[182] ^ t[183];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[184] | t[113]);
  assign t[153] = ~(t[229]);
  assign t[154] = ~(t[226]);
  assign t[155] = t[101] ^ t[73];
  assign t[156] = ~t[185];
  assign t[157] = t[186];
  assign t[158] = ~(t[116] ^ t[160]);
  assign t[159] = t[118] ^ t[177];
  assign t[15] = ~(t[27]);
  assign t[160] = t[187] ^ t[143];
  assign t[161] = t[188] & t[189];
  assign t[162] = ~(t[99]);
  assign t[163] = ~(t[183]);
  assign t[164] = ~(t[55]);
  assign t[165] = ~(t[56]);
  assign t[166] = t[28] ? x[81] : x[80];
  assign t[167] = t[132] ? x[83] : x[82];
  assign t[168] = t[132] ? x[85] : x[84];
  assign t[169] = t[227] ^ t[190];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[15]);
  assign t[171] = t[228] ^ t[191];
  assign t[172] = ~(t[175]);
  assign t[173] = ~(t[107]);
  assign t[174] = t[66] ^ t[107];
  assign t[175] = t[148] ^ t[99];
  assign t[176] = ~(t[157]);
  assign t[177] = t[192];
  assign t[178] = t[27] ? t[193] : t[230];
  assign t[179] = t[28] ? x[90] : x[89];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[27] ? t[194] : t[231];
  assign t[181] = t[74] ^ t[55];
  assign t[182] = t[55] ^ t[68];
  assign t[183] = t[88] ^ t[56];
  assign t[184] = ~(t[213]);
  assign t[185] = t[27] ? t[195] : t[232];
  assign t[186] = t[27] ? t[196] : t[233];
  assign t[187] = t[197] & t[198];
  assign t[188] = ~(t[187] ^ t[199]);
  assign t[189] = t[142] ^ t[200];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[28] ? x[101] : x[100];
  assign t[191] = t[201] ? x[103] : x[102];
  assign t[192] = t[27] ? t[202] : t[234];
  assign t[193] = t[230] ^ t[203];
  assign t[194] = t[231] ^ t[204];
  assign t[195] = t[232] ^ t[205];
  assign t[196] = t[233] ^ t[206];
  assign t[197] = ~(t[200]);
  assign t[198] = ~(t[156]);
  assign t[199] = t[118] ^ t[156];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[177] ^ t[157];
  assign t[201] = ~(t[49]);
  assign t[202] = t[234] ^ t[207];
  assign t[203] = t[79] ? x[108] : x[107];
  assign t[204] = t[79] ? x[110] : x[109];
  assign t[205] = t[79] ? x[112] : x[111];
  assign t[206] = t[201] ? x[114] : x[113];
  assign t[207] = t[201] ? x[116] : x[115];
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = t[262] ^ x[4];
  assign t[236] = t[263] ^ x[9];
  assign t[237] = t[264] ^ x[12];
  assign t[238] = t[265] ^ x[15];
  assign t[239] = t[266] ^ x[18];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[21];
  assign t[241] = t[268] ^ x[24];
  assign t[242] = t[269] ^ x[27];
  assign t[243] = t[270] ^ x[30];
  assign t[244] = t[271] ^ x[33];
  assign t[245] = t[272] ^ x[36];
  assign t[246] = t[273] ^ x[39];
  assign t[247] = t[274] ^ x[42];
  assign t[248] = t[275] ^ x[45];
  assign t[249] = t[276] ^ x[48];
  assign t[24] = ~(t[33] ^ t[43]);
  assign t[250] = t[277] ^ x[53];
  assign t[251] = t[278] ^ x[56];
  assign t[252] = t[279] ^ x[59];
  assign t[253] = t[280] ^ x[62];
  assign t[254] = t[281] ^ x[71];
  assign t[255] = t[282] ^ x[74];
  assign t[256] = t[283] ^ x[79];
  assign t[257] = t[284] ^ x[88];
  assign t[258] = t[285] ^ x[93];
  assign t[259] = t[286] ^ x[96];
  assign t[25] = t[44] ^ t[45];
  assign t[260] = t[287] ^ x[99];
  assign t[261] = t[288] ^ x[106];
  assign t[262] = (t[289] & ~t[290]);
  assign t[263] = (t[291] & ~t[292]);
  assign t[264] = (t[293] & ~t[294]);
  assign t[265] = (t[295] & ~t[296]);
  assign t[266] = (t[297] & ~t[298]);
  assign t[267] = (t[299] & ~t[300]);
  assign t[268] = (t[301] & ~t[302]);
  assign t[269] = (t[303] & ~t[304]);
  assign t[26] = ~(t[46] ^ t[22]);
  assign t[270] = (t[305] & ~t[306]);
  assign t[271] = (t[307] & ~t[308]);
  assign t[272] = (t[309] & ~t[310]);
  assign t[273] = (t[311] & ~t[312]);
  assign t[274] = (t[313] & ~t[314]);
  assign t[275] = (t[315] & ~t[316]);
  assign t[276] = (t[317] & ~t[318]);
  assign t[277] = (t[319] & ~t[320]);
  assign t[278] = (t[321] & ~t[322]);
  assign t[279] = (t[323] & ~t[324]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[325] & ~t[326]);
  assign t[281] = (t[327] & ~t[328]);
  assign t[282] = (t[329] & ~t[330]);
  assign t[283] = (t[331] & ~t[332]);
  assign t[284] = (t[333] & ~t[334]);
  assign t[285] = (t[335] & ~t[336]);
  assign t[286] = (t[337] & ~t[338]);
  assign t[287] = (t[339] & ~t[340]);
  assign t[288] = (t[341] & ~t[342]);
  assign t[289] = t[343] ^ x[4];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[3];
  assign t[291] = t[345] ^ x[9];
  assign t[292] = t[346] ^ x[8];
  assign t[293] = t[347] ^ x[12];
  assign t[294] = t[348] ^ x[11];
  assign t[295] = t[349] ^ x[15];
  assign t[296] = t[350] ^ x[14];
  assign t[297] = t[351] ^ x[18];
  assign t[298] = t[352] ^ x[17];
  assign t[299] = t[353] ^ x[21];
  assign t[29] = ~(t[209]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[20];
  assign t[301] = t[355] ^ x[24];
  assign t[302] = t[356] ^ x[23];
  assign t[303] = t[357] ^ x[27];
  assign t[304] = t[358] ^ x[26];
  assign t[305] = t[359] ^ x[30];
  assign t[306] = t[360] ^ x[29];
  assign t[307] = t[361] ^ x[33];
  assign t[308] = t[362] ^ x[32];
  assign t[309] = t[363] ^ x[36];
  assign t[30] = ~(t[210]);
  assign t[310] = t[364] ^ x[35];
  assign t[311] = t[365] ^ x[39];
  assign t[312] = t[366] ^ x[38];
  assign t[313] = t[367] ^ x[42];
  assign t[314] = t[368] ^ x[41];
  assign t[315] = t[369] ^ x[45];
  assign t[316] = t[370] ^ x[44];
  assign t[317] = t[371] ^ x[48];
  assign t[318] = t[372] ^ x[47];
  assign t[319] = t[373] ^ x[53];
  assign t[31] = ~(t[211]);
  assign t[320] = t[374] ^ x[52];
  assign t[321] = t[375] ^ x[56];
  assign t[322] = t[376] ^ x[55];
  assign t[323] = t[377] ^ x[59];
  assign t[324] = t[378] ^ x[58];
  assign t[325] = t[379] ^ x[62];
  assign t[326] = t[380] ^ x[61];
  assign t[327] = t[381] ^ x[71];
  assign t[328] = t[382] ^ x[70];
  assign t[329] = t[383] ^ x[74];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[73];
  assign t[331] = t[385] ^ x[79];
  assign t[332] = t[386] ^ x[78];
  assign t[333] = t[387] ^ x[88];
  assign t[334] = t[388] ^ x[87];
  assign t[335] = t[389] ^ x[93];
  assign t[336] = t[390] ^ x[92];
  assign t[337] = t[391] ^ x[96];
  assign t[338] = t[392] ^ x[95];
  assign t[339] = t[393] ^ x[99];
  assign t[33] = ~(t[52] ^ t[46]);
  assign t[340] = t[394] ^ x[98];
  assign t[341] = t[395] ^ x[106];
  assign t[342] = t[396] ^ x[105];
  assign t[343] = (x[2]);
  assign t[344] = (x[2]);
  assign t[345] = (x[7]);
  assign t[346] = (x[7]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[51]);
  assign t[374] = (x[51]);
  assign t[375] = (x[54]);
  assign t[376] = (x[54]);
  assign t[377] = (x[57]);
  assign t[378] = (x[57]);
  assign t[379] = (x[60]);
  assign t[37] = t[59] ^ t[39];
  assign t[380] = (x[60]);
  assign t[381] = (x[69]);
  assign t[382] = (x[69]);
  assign t[383] = (x[72]);
  assign t[384] = (x[72]);
  assign t[385] = (x[77]);
  assign t[386] = (x[77]);
  assign t[387] = (x[86]);
  assign t[388] = (x[86]);
  assign t[389] = (x[91]);
  assign t[38] = t[60] ^ t[61];
  assign t[390] = (x[91]);
  assign t[391] = (x[94]);
  assign t[392] = (x[94]);
  assign t[393] = (x[97]);
  assign t[394] = (x[97]);
  assign t[395] = (x[104]);
  assign t[396] = (x[104]);
  assign t[39] = t[8] ? t[62] : t[212];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[60] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = ~(t[70] ^ t[71]);
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = t[213] | t[78];
  assign t[49] = ~(t[79]);
  assign t[4] = t[8] ? t[9] : t[208];
  assign t[50] = ~(t[214]);
  assign t[51] = ~(t[80] & t[215]);
  assign t[52] = ~(t[81] ^ t[82]);
  assign t[53] = t[83] ^ t[84];
  assign t[54] = ~(t[43] ^ t[22]);
  assign t[55] = t[8] ? t[85] : t[216];
  assign t[56] = t[8] ? t[86] : t[217];
  assign t[57] = ~(t[35] ^ t[87]);
  assign t[58] = t[74] ^ t[88];
  assign t[59] = t[8] ? t[89] : t[218];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[65];
  assign t[61] = t[91] & t[92];
  assign t[62] = t[212] ^ t[93];
  assign t[63] = t[94] & t[95];
  assign t[64] = t[96] ^ t[39];
  assign t[65] = t[97] & t[98];
  assign t[66] = t[99] ^ t[100];
  assign t[67] = t[101] ^ t[102];
  assign t[68] = t[8] ? t[103] : t[219];
  assign t[69] = t[87] ^ t[36];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[104] ^ t[20];
  assign t[71] = ~(t[105] ^ t[106]);
  assign t[72] = t[107] ^ t[99];
  assign t[73] = t[108] & t[109];
  assign t[74] = t[56] ^ t[68];
  assign t[75] = t[87] ^ t[110];
  assign t[76] = ~(t[78] & t[111]);
  assign t[77] = ~(t[220] ^ t[112]);
  assign t[78] = ~(t[113] & t[114]);
  assign t[79] = ~(t[48]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[221]);
  assign t[81] = t[21] ^ t[115];
  assign t[82] = t[116] ^ t[117];
  assign t[83] = t[118] ^ t[119];
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[216] ^ t[122];
  assign t[86] = t[217] ^ t[123];
  assign t[87] = t[124] ^ t[125];
  assign t[88] = t[8] ? t[126] : t[222];
  assign t[89] = t[218] ^ t[127];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] & t[129];
  assign t[91] = ~(t[90] ^ t[130]);
  assign t[92] = t[64] ^ t[131];
  assign t[93] = t[132] ? x[50] : x[49];
  assign t[94] = ~(t[133] ^ t[60]);
  assign t[95] = t[37] ^ t[98];
  assign t[96] = t[8] ? t[134] : t[223];
  assign t[97] = ~(t[59]);
  assign t[98] = t[8] ? t[135] : t[224];
  assign t[99] = t[211] ^ t[136];
  assign t[9] = t[208] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[15]);
  assign t[101] = t[206] ^ t[136];
  assign t[102] = t[137] & t[138];
  assign t[103] = t[139] & t[124];
  assign t[104] = t[140] & t[141];
  assign t[105] = t[8] ? t[142] : t[213];
  assign t[106] = t[8] ? t[143] : t[214];
  assign t[107] = ~(t[69] ^ t[144]);
  assign t[108] = t[145] ^ t[146];
  assign t[109] = t[145] ^ t[147];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[148] ^ t[62];
  assign t[111] = t[89] ^ t[41];
  assign t[112] = t[35] ^ t[149];
  assign t[113] = t[8] ? t[150] : t[215];
  assign t[114] = t[144] ^ t[70];
  assign t[115] = ~(t[151] & t[152]);
  assign t[116] = t[153] ^ t[216];
  assign t[117] = ~(t[207]);
  assign t[118] = t[154] & t[153];
  assign t[119] = ~(t[155]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[8] ? t[156] : t[217];
  assign t[121] = t[209] ^ t[157];
  assign t[122] = t[210] ^ t[158];
  assign t[123] = t[27] ? t[159] : t[218];
  assign t[124] = t[208] ^ t[160];
  assign t[125] = t[211] ^ t[161];
  assign t[126] = ~(t[110] ^ t[63]);
  assign t[127] = t[39] ^ t[132];
  assign t[128] = t[212] ^ t[162];
  assign t[129] = ~(t[135]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = ~(t[148]);
  assign t[131] = ~(t[62]);
  assign t[132] = t[163];
  assign t[133] = t[39] ^ t[148];
  assign t[134] = t[148] ^ t[60];
  assign t[135] = t[132] ^ t[62];
  assign t[136] = t[164] ? x[75] : x[74];
  assign t[137] = ~(t[165]);
  assign t[138] = ~(t[89]);
  assign t[139] = ~(t[90]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = ~(t[102] ^ t[166]);
  assign t[141] = t[111] ^ t[165];
  assign t[142] = t[213] ^ t[167];
  assign t[143] = t[214] ^ t[168];
  assign t[144] = t[169] ^ t[170];
  assign t[145] = t[106] ^ t[113];
  assign t[146] = t[8] ? t[171] : t[219];
  assign t[147] = t[144] ^ t[172];
  assign t[148] = ~t[173];
  assign t[149] = t[174] & t[175];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[215] ^ t[176];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[177] | t[117]);
  assign t[153] = ~(t[220]);
  assign t[154] = ~(t[216]);
  assign t[155] = ~(t[28]);
  assign t[156] = t[217] ^ t[178];
  assign t[157] = t[119] ? x[83] : x[82];
  assign t[158] = t[119] ? x[85] : x[84];
  assign t[159] = t[218] ^ t[179];
  assign t[15] = ~(t[27]);
  assign t[160] = t[27] ? t[180] : t[221];
  assign t[161] = t[28] ? x[90] : x[89];
  assign t[162] = t[164] ? x[92] : x[91];
  assign t[163] = t[27] ? t[181] : t[222];
  assign t[164] = ~(t[155]);
  assign t[165] = t[124] ^ t[90];
  assign t[166] = t[67] ^ t[89];
  assign t[167] = t[182] ? x[97] : x[96];
  assign t[168] = t[182] ? x[99] : x[98];
  assign t[169] = t[183] & t[184];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[185] & t[146];
  assign t[171] = t[219] ^ t[186];
  assign t[172] = t[187] & t[188];
  assign t[173] = t[27] ? t[189] : t[223];
  assign t[174] = ~(t[190] ^ t[35]);
  assign t[175] = t[19] ^ t[85];
  assign t[176] = t[182] ? x[104] : x[103];
  assign t[177] = ~(t[204]);
  assign t[178] = t[119] ? x[106] : x[105];
  assign t[179] = t[119] ? x[108] : x[107];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[221] ^ t[191];
  assign t[181] = t[222] ^ t[192];
  assign t[182] = ~(t[155]);
  assign t[183] = ~(t[193]);
  assign t[184] = ~(t[105]);
  assign t[185] = ~(t[106]);
  assign t[186] = t[182] ? x[110] : x[109];
  assign t[187] = ~(t[169] ^ t[194]);
  assign t[188] = t[195] ^ t[193];
  assign t[189] = t[223] ^ t[196];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[120] ^ t[33];
  assign t[191] = t[28] ? x[112] : x[111];
  assign t[192] = t[164] ? x[114] : x[113];
  assign t[193] = t[146] ^ t[106];
  assign t[194] = t[145] ^ t[105];
  assign t[195] = t[105] ^ t[113];
  assign t[196] = t[28] ? x[116] : x[115];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = t[39] ^ t[40];
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[36];
  assign t[235] = t[262] ^ x[39];
  assign t[236] = t[263] ^ x[46];
  assign t[237] = t[264] ^ x[49];
  assign t[238] = t[265] ^ x[52];
  assign t[239] = t[266] ^ x[55];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[58];
  assign t[241] = t[268] ^ x[61];
  assign t[242] = t[269] ^ x[64];
  assign t[243] = t[270] ^ x[67];
  assign t[244] = t[271] ^ x[70];
  assign t[245] = t[272] ^ x[73];
  assign t[246] = t[273] ^ x[78];
  assign t[247] = t[274] ^ x[81];
  assign t[248] = t[275] ^ x[88];
  assign t[249] = t[276] ^ x[95];
  assign t[24] = t[43] ^ t[44];
  assign t[250] = t[277] ^ x[102];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = ~(t[45] ^ t[11]);
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[36];
  assign t[299] = t[353] ^ x[35];
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[39];
  assign t[301] = t[355] ^ x[38];
  assign t[302] = t[356] ^ x[46];
  assign t[303] = t[357] ^ x[45];
  assign t[304] = t[358] ^ x[49];
  assign t[305] = t[359] ^ x[48];
  assign t[306] = t[360] ^ x[52];
  assign t[307] = t[361] ^ x[51];
  assign t[308] = t[362] ^ x[55];
  assign t[309] = t[363] ^ x[54];
  assign t[30] = ~(t[199]);
  assign t[310] = t[364] ^ x[58];
  assign t[311] = t[365] ^ x[57];
  assign t[312] = t[366] ^ x[61];
  assign t[313] = t[367] ^ x[60];
  assign t[314] = t[368] ^ x[64];
  assign t[315] = t[369] ^ x[63];
  assign t[316] = t[370] ^ x[67];
  assign t[317] = t[371] ^ x[66];
  assign t[318] = t[372] ^ x[70];
  assign t[319] = t[373] ^ x[69];
  assign t[31] = ~(t[200]);
  assign t[320] = t[374] ^ x[73];
  assign t[321] = t[375] ^ x[72];
  assign t[322] = t[376] ^ x[78];
  assign t[323] = t[377] ^ x[77];
  assign t[324] = t[378] ^ x[81];
  assign t[325] = t[379] ^ x[80];
  assign t[326] = t[380] ^ x[88];
  assign t[327] = t[381] ^ x[87];
  assign t[328] = t[382] ^ x[95];
  assign t[329] = t[383] ^ x[94];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[102];
  assign t[331] = t[385] ^ x[101];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = t[8] ? t[52] : t[201];
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = t[8] ? t[53] : t[202];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[34]);
  assign t[353] = (x[34]);
  assign t[354] = (x[37]);
  assign t[355] = (x[37]);
  assign t[356] = (x[44]);
  assign t[357] = (x[44]);
  assign t[358] = (x[47]);
  assign t[359] = (x[47]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[50]);
  assign t[361] = (x[50]);
  assign t[362] = (x[53]);
  assign t[363] = (x[53]);
  assign t[364] = (x[56]);
  assign t[365] = (x[56]);
  assign t[366] = (x[59]);
  assign t[367] = (x[59]);
  assign t[368] = (x[62]);
  assign t[369] = (x[62]);
  assign t[36] = t[56] & t[57];
  assign t[370] = (x[65]);
  assign t[371] = (x[65]);
  assign t[372] = (x[68]);
  assign t[373] = (x[68]);
  assign t[374] = (x[71]);
  assign t[375] = (x[71]);
  assign t[376] = (x[76]);
  assign t[377] = (x[76]);
  assign t[378] = (x[79]);
  assign t[379] = (x[79]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[86]);
  assign t[381] = (x[86]);
  assign t[382] = (x[93]);
  assign t[383] = (x[93]);
  assign t[384] = (x[100]);
  assign t[385] = (x[100]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[62] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[203] ^ t[65];
  assign t[42] = t[66] ^ t[59];
  assign t[43] = t[67] ^ t[68];
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[71] ^ t[72]);
  assign t[46] = t[22] ^ t[73];
  assign t[47] = ~(t[74] ^ t[75]);
  assign t[48] = ~(t[76] & t[77]);
  assign t[49] = t[204] | t[78];
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[203]);
  assign t[51] = ~(t[79] & t[205]);
  assign t[52] = t[201] ^ t[80];
  assign t[53] = t[202] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = t[84] & t[85];
  assign t[56] = ~(t[54] ^ t[86]);
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] ^ t[90];
  assign t[59] = t[91] & t[92];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93];
  assign t[61] = t[63] ^ t[94];
  assign t[62] = t[95];
  assign t[63] = t[96] ^ t[97];
  assign t[64] = t[98] & t[99];
  assign t[65] = t[100] ? t[101] : t[206];
  assign t[66] = t[102] ^ t[103];
  assign t[67] = t[90] ^ t[41];
  assign t[68] = t[66] ^ t[104];
  assign t[69] = t[105] ^ t[106];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[107] & t[108];
  assign t[71] = t[109] ^ t[23];
  assign t[72] = t[110] ^ t[94];
  assign t[73] = t[111] ^ t[103];
  assign t[74] = t[34] ^ t[112];
  assign t[75] = t[113] ^ t[114];
  assign t[76] = ~(t[78] & t[115]);
  assign t[77] = ~(t[207] ^ t[116]);
  assign t[78] = ~(t[117] & t[118]);
  assign t[79] = ~(t[208]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[119] ? x[41] : x[40];
  assign t[81] = t[119] ? x[43] : x[42];
  assign t[82] = ~(t[88]);
  assign t[83] = ~(t[120]);
  assign t[84] = ~(t[33]);
  assign t[85] = t[8] ? t[121] : t[209];
  assign t[86] = t[19] ^ t[120];
  assign t[87] = t[120] ^ t[34];
  assign t[88] = t[85] ^ t[33];
  assign t[89] = t[27] ? t[122] : t[210];
  assign t[8] = ~(t[15]);
  assign t[90] = t[200] ^ t[123];
  assign t[91] = ~(t[58] ^ t[66]);
  assign t[92] = t[67] ^ t[124];
  assign t[93] = t[27] ? t[125] : t[211];
  assign t[94] = t[126] & t[127];
  assign t[95] = t[27] ? t[128] : t[212];
  assign t[96] = t[129] & t[130];
  assign t[97] = t[131] & t[132];
  assign t[98] = ~(t[96] ^ t[133]);
  assign t[99] = t[134] ^ t[135];
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[15]);
  assign t[101] = t[206] ^ t[136];
  assign t[102] = t[137] & t[138];
  assign t[103] = t[139] & t[124];
  assign t[104] = t[140] & t[141];
  assign t[105] = t[8] ? t[142] : t[213];
  assign t[106] = t[8] ? t[143] : t[214];
  assign t[107] = ~(t[69] ^ t[144]);
  assign t[108] = t[145] ^ t[146];
  assign t[109] = t[145] ^ t[147];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[148] ^ t[62];
  assign t[111] = t[89] ^ t[41];
  assign t[112] = t[35] ^ t[149];
  assign t[113] = t[8] ? t[150] : t[215];
  assign t[114] = t[144] ^ t[70];
  assign t[115] = ~(t[151] & t[152]);
  assign t[116] = t[153] ^ t[216];
  assign t[117] = ~(t[207]);
  assign t[118] = t[154] & t[153];
  assign t[119] = ~(t[155]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[8] ? t[156] : t[217];
  assign t[121] = t[209] ^ t[157];
  assign t[122] = t[210] ^ t[158];
  assign t[123] = t[27] ? t[159] : t[218];
  assign t[124] = t[208] ^ t[160];
  assign t[125] = t[211] ^ t[161];
  assign t[126] = ~(t[110] ^ t[63]);
  assign t[127] = t[39] ^ t[132];
  assign t[128] = t[212] ^ t[162];
  assign t[129] = ~(t[135]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = ~(t[148]);
  assign t[131] = ~(t[62]);
  assign t[132] = t[163];
  assign t[133] = t[39] ^ t[148];
  assign t[134] = t[148] ^ t[60];
  assign t[135] = t[132] ^ t[62];
  assign t[136] = t[164] ? x[75] : x[74];
  assign t[137] = ~(t[165]);
  assign t[138] = ~(t[89]);
  assign t[139] = ~(t[90]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = ~(t[102] ^ t[166]);
  assign t[141] = t[111] ^ t[165];
  assign t[142] = t[213] ^ t[167];
  assign t[143] = t[214] ^ t[168];
  assign t[144] = t[169] ^ t[170];
  assign t[145] = t[106] ^ t[113];
  assign t[146] = t[8] ? t[171] : t[219];
  assign t[147] = t[144] ^ t[172];
  assign t[148] = ~t[173];
  assign t[149] = t[174] & t[175];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[215] ^ t[176];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[177] | t[117]);
  assign t[153] = ~(t[220]);
  assign t[154] = ~(t[216]);
  assign t[155] = ~(t[28]);
  assign t[156] = t[217] ^ t[178];
  assign t[157] = t[119] ? x[83] : x[82];
  assign t[158] = t[119] ? x[85] : x[84];
  assign t[159] = t[218] ^ t[179];
  assign t[15] = ~(t[27]);
  assign t[160] = t[27] ? t[180] : t[221];
  assign t[161] = t[28] ? x[90] : x[89];
  assign t[162] = t[164] ? x[92] : x[91];
  assign t[163] = t[27] ? t[181] : t[222];
  assign t[164] = ~(t[155]);
  assign t[165] = t[124] ^ t[90];
  assign t[166] = t[67] ^ t[89];
  assign t[167] = t[182] ? x[97] : x[96];
  assign t[168] = t[182] ? x[99] : x[98];
  assign t[169] = t[183] & t[184];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[185] & t[146];
  assign t[171] = t[219] ^ t[186];
  assign t[172] = t[187] & t[188];
  assign t[173] = t[27] ? t[189] : t[223];
  assign t[174] = ~(t[190] ^ t[35]);
  assign t[175] = t[19] ^ t[85];
  assign t[176] = t[182] ? x[104] : x[103];
  assign t[177] = ~(t[204]);
  assign t[178] = t[119] ? x[106] : x[105];
  assign t[179] = t[119] ? x[108] : x[107];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[221] ^ t[191];
  assign t[181] = t[222] ^ t[192];
  assign t[182] = ~(t[155]);
  assign t[183] = ~(t[193]);
  assign t[184] = ~(t[105]);
  assign t[185] = ~(t[106]);
  assign t[186] = t[182] ? x[110] : x[109];
  assign t[187] = ~(t[169] ^ t[194]);
  assign t[188] = t[195] ^ t[193];
  assign t[189] = t[223] ^ t[196];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[120] ^ t[33];
  assign t[191] = t[28] ? x[112] : x[111];
  assign t[192] = t[164] ? x[114] : x[113];
  assign t[193] = t[146] ^ t[106];
  assign t[194] = t[145] ^ t[105];
  assign t[195] = t[105] ^ t[113];
  assign t[196] = t[28] ? x[116] : x[115];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = t[39] ^ t[40];
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[36];
  assign t[235] = t[262] ^ x[39];
  assign t[236] = t[263] ^ x[46];
  assign t[237] = t[264] ^ x[49];
  assign t[238] = t[265] ^ x[52];
  assign t[239] = t[266] ^ x[55];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[58];
  assign t[241] = t[268] ^ x[61];
  assign t[242] = t[269] ^ x[64];
  assign t[243] = t[270] ^ x[67];
  assign t[244] = t[271] ^ x[70];
  assign t[245] = t[272] ^ x[73];
  assign t[246] = t[273] ^ x[78];
  assign t[247] = t[274] ^ x[81];
  assign t[248] = t[275] ^ x[88];
  assign t[249] = t[276] ^ x[95];
  assign t[24] = t[43] ^ t[44];
  assign t[250] = t[277] ^ x[102];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = ~(t[45] ^ t[11]);
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[36];
  assign t[299] = t[353] ^ x[35];
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[39];
  assign t[301] = t[355] ^ x[38];
  assign t[302] = t[356] ^ x[46];
  assign t[303] = t[357] ^ x[45];
  assign t[304] = t[358] ^ x[49];
  assign t[305] = t[359] ^ x[48];
  assign t[306] = t[360] ^ x[52];
  assign t[307] = t[361] ^ x[51];
  assign t[308] = t[362] ^ x[55];
  assign t[309] = t[363] ^ x[54];
  assign t[30] = ~(t[199]);
  assign t[310] = t[364] ^ x[58];
  assign t[311] = t[365] ^ x[57];
  assign t[312] = t[366] ^ x[61];
  assign t[313] = t[367] ^ x[60];
  assign t[314] = t[368] ^ x[64];
  assign t[315] = t[369] ^ x[63];
  assign t[316] = t[370] ^ x[67];
  assign t[317] = t[371] ^ x[66];
  assign t[318] = t[372] ^ x[70];
  assign t[319] = t[373] ^ x[69];
  assign t[31] = ~(t[200]);
  assign t[320] = t[374] ^ x[73];
  assign t[321] = t[375] ^ x[72];
  assign t[322] = t[376] ^ x[78];
  assign t[323] = t[377] ^ x[77];
  assign t[324] = t[378] ^ x[81];
  assign t[325] = t[379] ^ x[80];
  assign t[326] = t[380] ^ x[88];
  assign t[327] = t[381] ^ x[87];
  assign t[328] = t[382] ^ x[95];
  assign t[329] = t[383] ^ x[94];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[102];
  assign t[331] = t[385] ^ x[101];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = t[8] ? t[52] : t[201];
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = t[8] ? t[53] : t[202];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[34]);
  assign t[353] = (x[34]);
  assign t[354] = (x[37]);
  assign t[355] = (x[37]);
  assign t[356] = (x[44]);
  assign t[357] = (x[44]);
  assign t[358] = (x[47]);
  assign t[359] = (x[47]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[50]);
  assign t[361] = (x[50]);
  assign t[362] = (x[53]);
  assign t[363] = (x[53]);
  assign t[364] = (x[56]);
  assign t[365] = (x[56]);
  assign t[366] = (x[59]);
  assign t[367] = (x[59]);
  assign t[368] = (x[62]);
  assign t[369] = (x[62]);
  assign t[36] = t[56] & t[57];
  assign t[370] = (x[65]);
  assign t[371] = (x[65]);
  assign t[372] = (x[68]);
  assign t[373] = (x[68]);
  assign t[374] = (x[71]);
  assign t[375] = (x[71]);
  assign t[376] = (x[76]);
  assign t[377] = (x[76]);
  assign t[378] = (x[79]);
  assign t[379] = (x[79]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[86]);
  assign t[381] = (x[86]);
  assign t[382] = (x[93]);
  assign t[383] = (x[93]);
  assign t[384] = (x[100]);
  assign t[385] = (x[100]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[62] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[203] ^ t[65];
  assign t[42] = t[66] ^ t[59];
  assign t[43] = t[67] ^ t[68];
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[71] ^ t[72]);
  assign t[46] = t[22] ^ t[73];
  assign t[47] = ~(t[74] ^ t[75]);
  assign t[48] = ~(t[76] & t[77]);
  assign t[49] = t[204] | t[78];
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[203]);
  assign t[51] = ~(t[79] & t[205]);
  assign t[52] = t[201] ^ t[80];
  assign t[53] = t[202] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = t[84] & t[85];
  assign t[56] = ~(t[54] ^ t[86]);
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] ^ t[90];
  assign t[59] = t[91] & t[92];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93];
  assign t[61] = t[63] ^ t[94];
  assign t[62] = t[95];
  assign t[63] = t[96] ^ t[97];
  assign t[64] = t[98] & t[99];
  assign t[65] = t[100] ? t[101] : t[206];
  assign t[66] = t[102] ^ t[103];
  assign t[67] = t[90] ^ t[41];
  assign t[68] = t[66] ^ t[104];
  assign t[69] = t[105] ^ t[106];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[107] & t[108];
  assign t[71] = t[109] ^ t[23];
  assign t[72] = t[110] ^ t[94];
  assign t[73] = t[111] ^ t[103];
  assign t[74] = t[34] ^ t[112];
  assign t[75] = t[113] ^ t[114];
  assign t[76] = ~(t[78] & t[115]);
  assign t[77] = ~(t[207] ^ t[116]);
  assign t[78] = ~(t[117] & t[118]);
  assign t[79] = ~(t[208]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[119] ? x[41] : x[40];
  assign t[81] = t[119] ? x[43] : x[42];
  assign t[82] = ~(t[88]);
  assign t[83] = ~(t[120]);
  assign t[84] = ~(t[33]);
  assign t[85] = t[8] ? t[121] : t[209];
  assign t[86] = t[19] ^ t[120];
  assign t[87] = t[120] ^ t[34];
  assign t[88] = t[85] ^ t[33];
  assign t[89] = t[27] ? t[122] : t[210];
  assign t[8] = ~(t[15]);
  assign t[90] = t[200] ^ t[123];
  assign t[91] = ~(t[58] ^ t[66]);
  assign t[92] = t[67] ^ t[124];
  assign t[93] = t[27] ? t[125] : t[211];
  assign t[94] = t[126] & t[127];
  assign t[95] = t[27] ? t[128] : t[212];
  assign t[96] = t[129] & t[130];
  assign t[97] = t[131] & t[132];
  assign t[98] = ~(t[96] ^ t[133]);
  assign t[99] = t[134] ^ t[135];
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[88]);
  assign t[101] = t[8] ? t[137] : t[214];
  assign t[102] = t[88] ^ t[23];
  assign t[103] = t[138] ? x[61] : x[60];
  assign t[104] = t[138] ? x[63] : x[62];
  assign t[105] = t[139] & t[140];
  assign t[106] = t[141] & t[72];
  assign t[107] = t[8] ? t[142] : t[215];
  assign t[108] = t[207] ^ t[143];
  assign t[109] = ~(t[144] & t[145]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[146] ^ t[216];
  assign t[111] = ~(t[208]);
  assign t[112] = t[147] & t[146];
  assign t[113] = t[148] ^ t[65];
  assign t[114] = ~(t[149] ^ t[39]);
  assign t[115] = t[150] ^ t[151];
  assign t[116] = t[43] ^ t[107];
  assign t[117] = t[70] ^ t[26];
  assign t[118] = t[210] ^ t[152];
  assign t[119] = t[153] ? t[154] : t[217];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[201] ^ t[155];
  assign t[121] = t[27] ? t[156] : t[218];
  assign t[122] = t[157] & t[158];
  assign t[123] = t[159] ^ t[54];
  assign t[124] = t[160] & t[161];
  assign t[125] = t[211] ^ t[162];
  assign t[126] = t[212] ^ t[163];
  assign t[127] = t[27] ? t[164] : t[219];
  assign t[128] = t[165];
  assign t[129] = t[27] ? t[166] : t[220];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[167] & t[168];
  assign t[131] = t[213] ^ t[169];
  assign t[132] = t[170] & t[171];
  assign t[133] = ~(t[172] ^ t[95]);
  assign t[134] = t[150] ^ t[91];
  assign t[135] = ~(t[28]);
  assign t[136] = t[101] ^ t[88];
  assign t[137] = t[214] ^ t[173];
  assign t[138] = ~(t[135]);
  assign t[139] = ~(t[174]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[43]);
  assign t[141] = ~(t[44]);
  assign t[142] = t[215] ^ t[175];
  assign t[143] = t[138] ? x[83] : x[82];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[176] | t[111]);
  assign t[146] = ~(t[221]);
  assign t[147] = ~(t[216]);
  assign t[148] = t[87] ^ t[23];
  assign t[149] = t[177] ^ t[124];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[128] ^ t[61];
  assign t[151] = t[95] ^ t[178];
  assign t[152] = t[97] ? x[88] : x[87];
  assign t[153] = ~(t[15]);
  assign t[154] = t[217] ^ t[179];
  assign t[155] = t[27] ? t[180] : t[222];
  assign t[156] = t[218] ^ t[181];
  assign t[157] = ~(t[105] ^ t[182]);
  assign t[158] = t[116] ^ t[174];
  assign t[159] = t[183] & t[184];
  assign t[15] = ~(t[27]);
  assign t[160] = ~(t[177] ^ t[123]);
  assign t[161] = t[92] ^ t[84];
  assign t[162] = t[97] ? x[93] : x[92];
  assign t[163] = t[97] ? x[95] : x[94];
  assign t[164] = t[219] ^ t[185];
  assign t[165] = t[27] ? t[186] : t[223];
  assign t[166] = t[220] ^ t[187];
  assign t[167] = ~(t[159] ^ t[188]);
  assign t[168] = t[53] ^ t[189];
  assign t[169] = t[28] ? x[100] : x[99];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[190]);
  assign t[171] = ~(t[89]);
  assign t[172] = t[89] ^ t[128];
  assign t[173] = t[97] ? x[102] : x[101];
  assign t[174] = t[72] ^ t[44];
  assign t[175] = t[138] ? x[104] : x[103];
  assign t[176] = ~(t[204]);
  assign t[177] = t[81] ^ t[120];
  assign t[178] = t[191] & t[192];
  assign t[179] = t[193] ? x[106] : x[105];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[222] ^ t[194];
  assign t[181] = t[28] ? x[108] : x[107];
  assign t[182] = t[71] ^ t[43];
  assign t[183] = ~(t[189]);
  assign t[184] = ~(t[81]);
  assign t[185] = t[28] ? x[110] : x[109];
  assign t[186] = t[223] ^ t[195];
  assign t[187] = t[193] ? x[112] : x[111];
  assign t[188] = t[92] ^ t[81];
  assign t[189] = t[84] ^ t[120];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[91] ^ t[128];
  assign t[191] = ~(t[132] ^ t[196]);
  assign t[192] = t[58] ^ t[190];
  assign t[193] = ~(t[135]);
  assign t[194] = t[97] ? x[114] : x[113];
  assign t[195] = t[193] ? x[116] : x[115];
  assign t[196] = t[150] ^ t[89];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[36];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = ~(t[38] ^ t[39]);
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[38];
  assign t[235] = t[262] ^ x[41];
  assign t[236] = t[263] ^ x[44];
  assign t[237] = t[264] ^ x[47];
  assign t[238] = t[265] ^ x[50];
  assign t[239] = t[266] ^ x[53];
  assign t[23] = t[8] ? t[40] : t[198];
  assign t[240] = t[267] ^ x[56];
  assign t[241] = t[268] ^ x[59];
  assign t[242] = t[269] ^ x[66];
  assign t[243] = t[270] ^ x[69];
  assign t[244] = t[271] ^ x[72];
  assign t[245] = t[272] ^ x[75];
  assign t[246] = t[273] ^ x[78];
  assign t[247] = t[274] ^ x[81];
  assign t[248] = t[275] ^ x[86];
  assign t[249] = t[276] ^ x[91];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[277] ^ x[98];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = t[43] ^ t[44];
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = t[45] & t[46];
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[48]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[38];
  assign t[299] = t[353] ^ x[37];
  assign t[29] = ~(t[199]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[41];
  assign t[301] = t[355] ^ x[40];
  assign t[302] = t[356] ^ x[44];
  assign t[303] = t[357] ^ x[43];
  assign t[304] = t[358] ^ x[47];
  assign t[305] = t[359] ^ x[46];
  assign t[306] = t[360] ^ x[50];
  assign t[307] = t[361] ^ x[49];
  assign t[308] = t[362] ^ x[53];
  assign t[309] = t[363] ^ x[52];
  assign t[30] = ~(t[200]);
  assign t[310] = t[364] ^ x[56];
  assign t[311] = t[365] ^ x[55];
  assign t[312] = t[366] ^ x[59];
  assign t[313] = t[367] ^ x[58];
  assign t[314] = t[368] ^ x[66];
  assign t[315] = t[369] ^ x[65];
  assign t[316] = t[370] ^ x[69];
  assign t[317] = t[371] ^ x[68];
  assign t[318] = t[372] ^ x[72];
  assign t[319] = t[373] ^ x[71];
  assign t[31] = ~(t[201]);
  assign t[320] = t[374] ^ x[75];
  assign t[321] = t[375] ^ x[74];
  assign t[322] = t[376] ^ x[78];
  assign t[323] = t[377] ^ x[77];
  assign t[324] = t[378] ^ x[81];
  assign t[325] = t[379] ^ x[80];
  assign t[326] = t[380] ^ x[86];
  assign t[327] = t[381] ^ x[85];
  assign t[328] = t[382] ^ x[91];
  assign t[329] = t[383] ^ x[90];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[98];
  assign t[331] = t[385] ^ x[97];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = ~(t[51] ^ t[52]);
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = t[53] ^ t[54];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[36]);
  assign t[353] = (x[36]);
  assign t[354] = (x[39]);
  assign t[355] = (x[39]);
  assign t[356] = (x[42]);
  assign t[357] = (x[42]);
  assign t[358] = (x[45]);
  assign t[359] = (x[45]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[48]);
  assign t[361] = (x[48]);
  assign t[362] = (x[51]);
  assign t[363] = (x[51]);
  assign t[364] = (x[54]);
  assign t[365] = (x[54]);
  assign t[366] = (x[57]);
  assign t[367] = (x[57]);
  assign t[368] = (x[64]);
  assign t[369] = (x[64]);
  assign t[36] = t[57] ^ t[42];
  assign t[370] = (x[67]);
  assign t[371] = (x[67]);
  assign t[372] = (x[70]);
  assign t[373] = (x[70]);
  assign t[374] = (x[73]);
  assign t[375] = (x[73]);
  assign t[376] = (x[76]);
  assign t[377] = (x[76]);
  assign t[378] = (x[79]);
  assign t[379] = (x[79]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[84]);
  assign t[381] = (x[84]);
  assign t[382] = (x[89]);
  assign t[383] = (x[89]);
  assign t[384] = (x[96]);
  assign t[385] = (x[96]);
  assign t[38] = t[60] ^ t[14];
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[198] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] & t[67];
  assign t[43] = t[8] ? t[68] : t[202];
  assign t[44] = t[8] ? t[69] : t[203];
  assign t[45] = ~(t[25] ^ t[70]);
  assign t[46] = t[71] ^ t[72];
  assign t[47] = ~(t[73] & t[74]);
  assign t[48] = t[204] | t[75];
  assign t[49] = ~(t[205]);
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[76] & t[206]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[71] ^ t[85];
  assign t[56] = t[82] ^ t[86];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] ^ t[61];
  assign t[59] = t[90] & t[91];
  assign t[5] = ~(t[10]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[94];
  assign t[62] = t[95] ^ t[96];
  assign t[63] = t[97] ? x[35] : x[34];
  assign t[64] = t[98] & t[99];
  assign t[65] = t[100] & t[101];
  assign t[66] = ~(t[57] ^ t[41]);
  assign t[67] = t[102] ^ t[101];
  assign t[68] = t[202] ^ t[103];
  assign t[69] = t[203] ^ t[104];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[105] ^ t[106];
  assign t[71] = t[44] ^ t[107];
  assign t[72] = t[8] ? t[108] : t[207];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[208] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[209]);
  assign t[77] = t[13] ^ t[113];
  assign t[78] = ~(t[114] ^ t[115]);
  assign t[79] = t[116] ^ t[106];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[107] ^ t[117];
  assign t[81] = t[27] ? t[118] : t[210];
  assign t[82] = t[205] ^ t[119];
  assign t[83] = ~(t[120]);
  assign t[84] = t[209] ^ t[121];
  assign t[85] = t[70] ^ t[122];
  assign t[86] = t[123] ^ t[124];
  assign t[87] = t[8] ? t[125] : t[211];
  assign t[88] = t[8] ? t[126] : t[212];
  assign t[89] = ~t[127];
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[128]);
  assign t[91] = t[129];
  assign t[92] = t[120] ^ t[82];
  assign t[93] = t[123] ^ t[130];
  assign t[94] = t[27] ? t[131] : t[213];
  assign t[95] = t[132] ^ t[59];
  assign t[96] = t[133] & t[134];
  assign t[97] = ~(t[135]);
  assign t[98] = ~(t[136]);
  assign t[99] = ~(t[87]);
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[88]);
  assign t[101] = t[8] ? t[137] : t[214];
  assign t[102] = t[88] ^ t[23];
  assign t[103] = t[138] ? x[61] : x[60];
  assign t[104] = t[138] ? x[63] : x[62];
  assign t[105] = t[139] & t[140];
  assign t[106] = t[141] & t[72];
  assign t[107] = t[8] ? t[142] : t[215];
  assign t[108] = t[207] ^ t[143];
  assign t[109] = ~(t[144] & t[145]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[146] ^ t[216];
  assign t[111] = ~(t[208]);
  assign t[112] = t[147] & t[146];
  assign t[113] = t[148] ^ t[65];
  assign t[114] = ~(t[149] ^ t[39]);
  assign t[115] = t[150] ^ t[151];
  assign t[116] = t[43] ^ t[107];
  assign t[117] = t[70] ^ t[26];
  assign t[118] = t[210] ^ t[152];
  assign t[119] = t[153] ? t[154] : t[217];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[201] ^ t[155];
  assign t[121] = t[27] ? t[156] : t[218];
  assign t[122] = t[157] & t[158];
  assign t[123] = t[159] ^ t[54];
  assign t[124] = t[160] & t[161];
  assign t[125] = t[211] ^ t[162];
  assign t[126] = t[212] ^ t[163];
  assign t[127] = t[27] ? t[164] : t[219];
  assign t[128] = t[165];
  assign t[129] = t[27] ? t[166] : t[220];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[167] & t[168];
  assign t[131] = t[213] ^ t[169];
  assign t[132] = t[170] & t[171];
  assign t[133] = ~(t[172] ^ t[95]);
  assign t[134] = t[150] ^ t[91];
  assign t[135] = ~(t[28]);
  assign t[136] = t[101] ^ t[88];
  assign t[137] = t[214] ^ t[173];
  assign t[138] = ~(t[135]);
  assign t[139] = ~(t[174]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[43]);
  assign t[141] = ~(t[44]);
  assign t[142] = t[215] ^ t[175];
  assign t[143] = t[138] ? x[83] : x[82];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[176] | t[111]);
  assign t[146] = ~(t[221]);
  assign t[147] = ~(t[216]);
  assign t[148] = t[87] ^ t[23];
  assign t[149] = t[177] ^ t[124];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[128] ^ t[61];
  assign t[151] = t[95] ^ t[178];
  assign t[152] = t[97] ? x[88] : x[87];
  assign t[153] = ~(t[15]);
  assign t[154] = t[217] ^ t[179];
  assign t[155] = t[27] ? t[180] : t[222];
  assign t[156] = t[218] ^ t[181];
  assign t[157] = ~(t[105] ^ t[182]);
  assign t[158] = t[116] ^ t[174];
  assign t[159] = t[183] & t[184];
  assign t[15] = ~(t[27]);
  assign t[160] = ~(t[177] ^ t[123]);
  assign t[161] = t[92] ^ t[84];
  assign t[162] = t[97] ? x[93] : x[92];
  assign t[163] = t[97] ? x[95] : x[94];
  assign t[164] = t[219] ^ t[185];
  assign t[165] = t[27] ? t[186] : t[223];
  assign t[166] = t[220] ^ t[187];
  assign t[167] = ~(t[159] ^ t[188]);
  assign t[168] = t[53] ^ t[189];
  assign t[169] = t[28] ? x[100] : x[99];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[190]);
  assign t[171] = ~(t[89]);
  assign t[172] = t[89] ^ t[128];
  assign t[173] = t[97] ? x[102] : x[101];
  assign t[174] = t[72] ^ t[44];
  assign t[175] = t[138] ? x[104] : x[103];
  assign t[176] = ~(t[204]);
  assign t[177] = t[81] ^ t[120];
  assign t[178] = t[191] & t[192];
  assign t[179] = t[193] ? x[106] : x[105];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[222] ^ t[194];
  assign t[181] = t[28] ? x[108] : x[107];
  assign t[182] = t[71] ^ t[43];
  assign t[183] = ~(t[189]);
  assign t[184] = ~(t[81]);
  assign t[185] = t[28] ? x[110] : x[109];
  assign t[186] = t[223] ^ t[195];
  assign t[187] = t[193] ? x[112] : x[111];
  assign t[188] = t[92] ^ t[81];
  assign t[189] = t[84] ^ t[120];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[91] ^ t[128];
  assign t[191] = ~(t[132] ^ t[196]);
  assign t[192] = t[58] ^ t[190];
  assign t[193] = ~(t[135]);
  assign t[194] = t[97] ? x[114] : x[113];
  assign t[195] = t[193] ? x[116] : x[115];
  assign t[196] = t[150] ^ t[89];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[36];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = ~(t[38] ^ t[39]);
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[38];
  assign t[235] = t[262] ^ x[41];
  assign t[236] = t[263] ^ x[44];
  assign t[237] = t[264] ^ x[47];
  assign t[238] = t[265] ^ x[50];
  assign t[239] = t[266] ^ x[53];
  assign t[23] = t[8] ? t[40] : t[198];
  assign t[240] = t[267] ^ x[56];
  assign t[241] = t[268] ^ x[59];
  assign t[242] = t[269] ^ x[66];
  assign t[243] = t[270] ^ x[69];
  assign t[244] = t[271] ^ x[72];
  assign t[245] = t[272] ^ x[75];
  assign t[246] = t[273] ^ x[78];
  assign t[247] = t[274] ^ x[81];
  assign t[248] = t[275] ^ x[86];
  assign t[249] = t[276] ^ x[91];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[277] ^ x[98];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = t[43] ^ t[44];
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = t[45] & t[46];
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[48]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[38];
  assign t[299] = t[353] ^ x[37];
  assign t[29] = ~(t[199]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[41];
  assign t[301] = t[355] ^ x[40];
  assign t[302] = t[356] ^ x[44];
  assign t[303] = t[357] ^ x[43];
  assign t[304] = t[358] ^ x[47];
  assign t[305] = t[359] ^ x[46];
  assign t[306] = t[360] ^ x[50];
  assign t[307] = t[361] ^ x[49];
  assign t[308] = t[362] ^ x[53];
  assign t[309] = t[363] ^ x[52];
  assign t[30] = ~(t[200]);
  assign t[310] = t[364] ^ x[56];
  assign t[311] = t[365] ^ x[55];
  assign t[312] = t[366] ^ x[59];
  assign t[313] = t[367] ^ x[58];
  assign t[314] = t[368] ^ x[66];
  assign t[315] = t[369] ^ x[65];
  assign t[316] = t[370] ^ x[69];
  assign t[317] = t[371] ^ x[68];
  assign t[318] = t[372] ^ x[72];
  assign t[319] = t[373] ^ x[71];
  assign t[31] = ~(t[201]);
  assign t[320] = t[374] ^ x[75];
  assign t[321] = t[375] ^ x[74];
  assign t[322] = t[376] ^ x[78];
  assign t[323] = t[377] ^ x[77];
  assign t[324] = t[378] ^ x[81];
  assign t[325] = t[379] ^ x[80];
  assign t[326] = t[380] ^ x[86];
  assign t[327] = t[381] ^ x[85];
  assign t[328] = t[382] ^ x[91];
  assign t[329] = t[383] ^ x[90];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[98];
  assign t[331] = t[385] ^ x[97];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = ~(t[51] ^ t[52]);
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = t[53] ^ t[54];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[36]);
  assign t[353] = (x[36]);
  assign t[354] = (x[39]);
  assign t[355] = (x[39]);
  assign t[356] = (x[42]);
  assign t[357] = (x[42]);
  assign t[358] = (x[45]);
  assign t[359] = (x[45]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[48]);
  assign t[361] = (x[48]);
  assign t[362] = (x[51]);
  assign t[363] = (x[51]);
  assign t[364] = (x[54]);
  assign t[365] = (x[54]);
  assign t[366] = (x[57]);
  assign t[367] = (x[57]);
  assign t[368] = (x[64]);
  assign t[369] = (x[64]);
  assign t[36] = t[57] ^ t[42];
  assign t[370] = (x[67]);
  assign t[371] = (x[67]);
  assign t[372] = (x[70]);
  assign t[373] = (x[70]);
  assign t[374] = (x[73]);
  assign t[375] = (x[73]);
  assign t[376] = (x[76]);
  assign t[377] = (x[76]);
  assign t[378] = (x[79]);
  assign t[379] = (x[79]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[84]);
  assign t[381] = (x[84]);
  assign t[382] = (x[89]);
  assign t[383] = (x[89]);
  assign t[384] = (x[96]);
  assign t[385] = (x[96]);
  assign t[38] = t[60] ^ t[14];
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[198] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] & t[67];
  assign t[43] = t[8] ? t[68] : t[202];
  assign t[44] = t[8] ? t[69] : t[203];
  assign t[45] = ~(t[25] ^ t[70]);
  assign t[46] = t[71] ^ t[72];
  assign t[47] = ~(t[73] & t[74]);
  assign t[48] = t[204] | t[75];
  assign t[49] = ~(t[205]);
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[76] & t[206]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[71] ^ t[85];
  assign t[56] = t[82] ^ t[86];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] ^ t[61];
  assign t[59] = t[90] & t[91];
  assign t[5] = ~(t[10]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[94];
  assign t[62] = t[95] ^ t[96];
  assign t[63] = t[97] ? x[35] : x[34];
  assign t[64] = t[98] & t[99];
  assign t[65] = t[100] & t[101];
  assign t[66] = ~(t[57] ^ t[41]);
  assign t[67] = t[102] ^ t[101];
  assign t[68] = t[202] ^ t[103];
  assign t[69] = t[203] ^ t[104];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[105] ^ t[106];
  assign t[71] = t[44] ^ t[107];
  assign t[72] = t[8] ? t[108] : t[207];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[208] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[209]);
  assign t[77] = t[13] ^ t[113];
  assign t[78] = ~(t[114] ^ t[115]);
  assign t[79] = t[116] ^ t[106];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[107] ^ t[117];
  assign t[81] = t[27] ? t[118] : t[210];
  assign t[82] = t[205] ^ t[119];
  assign t[83] = ~(t[120]);
  assign t[84] = t[209] ^ t[121];
  assign t[85] = t[70] ^ t[122];
  assign t[86] = t[123] ^ t[124];
  assign t[87] = t[8] ? t[125] : t[211];
  assign t[88] = t[8] ? t[126] : t[212];
  assign t[89] = ~t[127];
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[128]);
  assign t[91] = t[129];
  assign t[92] = t[120] ^ t[82];
  assign t[93] = t[123] ^ t[130];
  assign t[94] = t[27] ? t[131] : t[213];
  assign t[95] = t[132] ^ t[59];
  assign t[96] = t[133] & t[134];
  assign t[97] = ~(t[135]);
  assign t[98] = ~(t[136]);
  assign t[99] = ~(t[87]);
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind96(x, y);
 input [116:0] x;
 output y;

 wire [378:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[134] ? t[135] : t[209];
  assign t[101] = t[191] ^ t[136];
  assign t[102] = ~(t[68] ^ t[137]);
  assign t[103] = t[138] ^ t[139];
  assign t[104] = t[140] & t[141];
  assign t[105] = ~(t[104] ^ t[142]);
  assign t[106] = t[19] ^ t[143];
  assign t[107] = ~(t[144] & t[145]);
  assign t[108] = t[146] ^ t[210];
  assign t[109] = ~(t[202]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[147] & t[146];
  assign t[111] = t[130] ? x[72] : x[71];
  assign t[112] = t[130] ? x[74] : x[73];
  assign t[113] = t[204] ^ t[148];
  assign t[114] = t[130] ? x[76] : x[75];
  assign t[115] = t[100] ^ t[121];
  assign t[116] = t[149] & t[139];
  assign t[117] = t[33] ^ t[54];
  assign t[118] = t[150] & t[151];
  assign t[119] = t[126] ^ t[152];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[153] ^ t[88];
  assign t[121] = t[198] ^ t[154];
  assign t[122] = t[137] ^ t[69];
  assign t[123] = t[205] ^ t[155];
  assign t[124] = t[206] ^ t[156];
  assign t[125] = t[157] ^ t[158];
  assign t[126] = t[85] ^ t[98];
  assign t[127] = t[27] ? t[159] : t[211];
  assign t[128] = ~(t[153] ^ t[42]);
  assign t[129] = t[23] ^ t[94];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = ~(t[160]);
  assign t[131] = t[8] ? t[161] : t[212];
  assign t[132] = t[207] ^ t[162];
  assign t[133] = t[208] ^ t[163];
  assign t[134] = ~(t[15]);
  assign t[135] = t[209] ^ t[164];
  assign t[136] = t[134] ? t[165] : t[213];
  assign t[137] = t[166] ^ t[116];
  assign t[138] = t[101] ^ t[121];
  assign t[139] = t[192] ^ t[167];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[143]);
  assign t[141] = ~(t[33]);
  assign t[142] = t[46] ^ t[33];
  assign t[143] = t[36] ^ t[54];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[168] | t[109]);
  assign t[146] = ~(t[214]);
  assign t[147] = ~(t[210]);
  assign t[148] = t[130] ? x[90] : x[89];
  assign t[149] = ~(t[101]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[117] ^ t[70]);
  assign t[151] = t[46] ^ t[36];
  assign t[152] = t[125] ^ t[169];
  assign t[153] = t[131] ^ t[40];
  assign t[154] = t[134] ? t[170] : t[215];
  assign t[155] = t[171] ? x[95] : x[94];
  assign t[156] = t[171] ? x[97] : x[96];
  assign t[157] = t[172] & t[173];
  assign t[158] = t[174] & t[127];
  assign t[159] = t[211] ^ t[175];
  assign t[15] = ~(t[27]);
  assign t[160] = ~(t[28]);
  assign t[161] = t[212] ^ t[176];
  assign t[162] = t[130] ? x[99] : x[98];
  assign t[163] = t[28] ? x[101] : x[100];
  assign t[164] = t[177] ? x[103] : x[102];
  assign t[165] = t[213] ^ t[178];
  assign t[166] = t[179] & t[180];
  assign t[167] = t[134] ? t[181] : t[216];
  assign t[168] = ~(t[196]);
  assign t[169] = t[182] & t[183];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[215] ^ t[184];
  assign t[171] = ~(t[160]);
  assign t[172] = ~(t[185]);
  assign t[173] = ~(t[84]);
  assign t[174] = ~(t[85]);
  assign t[175] = t[28] ? x[108] : x[107];
  assign t[176] = t[130] ? x[110] : x[109];
  assign t[177] = ~(t[160]);
  assign t[178] = t[177] ? x[112] : x[111];
  assign t[179] = ~(t[186]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[100]);
  assign t[181] = t[216] ^ t[187];
  assign t[182] = ~(t[157] ^ t[188]);
  assign t[183] = t[189] ^ t[185];
  assign t[184] = t[177] ? x[114] : x[113];
  assign t[185] = t[127] ^ t[85];
  assign t[186] = t[139] ^ t[101];
  assign t[187] = t[177] ? x[116] : x[115];
  assign t[188] = t[126] ^ t[84];
  assign t[189] = t[84] ^ t[98];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] & t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = t[244] ^ x[4];
  assign t[218] = t[245] ^ x[9];
  assign t[219] = t[246] ^ x[12];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[15];
  assign t[221] = t[248] ^ x[18];
  assign t[222] = t[249] ^ x[21];
  assign t[223] = t[250] ^ x[24];
  assign t[224] = t[251] ^ x[27];
  assign t[225] = t[252] ^ x[30];
  assign t[226] = t[253] ^ x[33];
  assign t[227] = t[254] ^ x[36];
  assign t[228] = t[255] ^ x[39];
  assign t[229] = t[256] ^ x[42];
  assign t[22] = ~(t[26] ^ t[39]);
  assign t[230] = t[257] ^ x[45];
  assign t[231] = t[258] ^ x[48];
  assign t[232] = t[259] ^ x[51];
  assign t[233] = t[260] ^ x[54];
  assign t[234] = t[261] ^ x[61];
  assign t[235] = t[262] ^ x[64];
  assign t[236] = t[263] ^ x[67];
  assign t[237] = t[264] ^ x[70];
  assign t[238] = t[265] ^ x[79];
  assign t[239] = t[266] ^ x[82];
  assign t[23] = t[40] ^ t[41];
  assign t[240] = t[267] ^ x[85];
  assign t[241] = t[268] ^ x[88];
  assign t[242] = t[269] ^ x[93];
  assign t[243] = t[270] ^ x[106];
  assign t[244] = (t[271] & ~t[272]);
  assign t[245] = (t[273] & ~t[274]);
  assign t[246] = (t[275] & ~t[276]);
  assign t[247] = (t[277] & ~t[278]);
  assign t[248] = (t[279] & ~t[280]);
  assign t[249] = (t[281] & ~t[282]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[283] & ~t[284]);
  assign t[251] = (t[285] & ~t[286]);
  assign t[252] = (t[287] & ~t[288]);
  assign t[253] = (t[289] & ~t[290]);
  assign t[254] = (t[291] & ~t[292]);
  assign t[255] = (t[293] & ~t[294]);
  assign t[256] = (t[295] & ~t[296]);
  assign t[257] = (t[297] & ~t[298]);
  assign t[258] = (t[299] & ~t[300]);
  assign t[259] = (t[301] & ~t[302]);
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[260] = (t[303] & ~t[304]);
  assign t[261] = (t[305] & ~t[306]);
  assign t[262] = (t[307] & ~t[308]);
  assign t[263] = (t[309] & ~t[310]);
  assign t[264] = (t[311] & ~t[312]);
  assign t[265] = (t[313] & ~t[314]);
  assign t[266] = (t[315] & ~t[316]);
  assign t[267] = (t[317] & ~t[318]);
  assign t[268] = (t[319] & ~t[320]);
  assign t[269] = (t[321] & ~t[322]);
  assign t[26] = t[46] ^ t[47];
  assign t[270] = (t[323] & ~t[324]);
  assign t[271] = t[325] ^ x[4];
  assign t[272] = t[326] ^ x[3];
  assign t[273] = t[327] ^ x[9];
  assign t[274] = t[328] ^ x[8];
  assign t[275] = t[329] ^ x[12];
  assign t[276] = t[330] ^ x[11];
  assign t[277] = t[331] ^ x[15];
  assign t[278] = t[332] ^ x[14];
  assign t[279] = t[333] ^ x[18];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[17];
  assign t[281] = t[335] ^ x[21];
  assign t[282] = t[336] ^ x[20];
  assign t[283] = t[337] ^ x[24];
  assign t[284] = t[338] ^ x[23];
  assign t[285] = t[339] ^ x[27];
  assign t[286] = t[340] ^ x[26];
  assign t[287] = t[341] ^ x[30];
  assign t[288] = t[342] ^ x[29];
  assign t[289] = t[343] ^ x[33];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[32];
  assign t[291] = t[345] ^ x[36];
  assign t[292] = t[346] ^ x[35];
  assign t[293] = t[347] ^ x[39];
  assign t[294] = t[348] ^ x[38];
  assign t[295] = t[349] ^ x[42];
  assign t[296] = t[350] ^ x[41];
  assign t[297] = t[351] ^ x[45];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[48];
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[47];
  assign t[301] = t[355] ^ x[51];
  assign t[302] = t[356] ^ x[50];
  assign t[303] = t[357] ^ x[54];
  assign t[304] = t[358] ^ x[53];
  assign t[305] = t[359] ^ x[61];
  assign t[306] = t[360] ^ x[60];
  assign t[307] = t[361] ^ x[64];
  assign t[308] = t[362] ^ x[63];
  assign t[309] = t[363] ^ x[67];
  assign t[30] = ~(t[192]);
  assign t[310] = t[364] ^ x[66];
  assign t[311] = t[365] ^ x[70];
  assign t[312] = t[366] ^ x[69];
  assign t[313] = t[367] ^ x[79];
  assign t[314] = t[368] ^ x[78];
  assign t[315] = t[369] ^ x[82];
  assign t[316] = t[370] ^ x[81];
  assign t[317] = t[371] ^ x[85];
  assign t[318] = t[372] ^ x[84];
  assign t[319] = t[373] ^ x[88];
  assign t[31] = ~(t[193]);
  assign t[320] = t[374] ^ x[87];
  assign t[321] = t[375] ^ x[93];
  assign t[322] = t[376] ^ x[92];
  assign t[323] = t[377] ^ x[106];
  assign t[324] = t[378] ^ x[105];
  assign t[325] = (x[2]);
  assign t[326] = (x[2]);
  assign t[327] = (x[7]);
  assign t[328] = (x[7]);
  assign t[329] = (x[10]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[10]);
  assign t[331] = (x[13]);
  assign t[332] = (x[13]);
  assign t[333] = (x[16]);
  assign t[334] = (x[16]);
  assign t[335] = (x[19]);
  assign t[336] = (x[19]);
  assign t[337] = (x[22]);
  assign t[338] = (x[22]);
  assign t[339] = (x[25]);
  assign t[33] = t[52];
  assign t[340] = (x[25]);
  assign t[341] = (x[28]);
  assign t[342] = (x[28]);
  assign t[343] = (x[31]);
  assign t[344] = (x[31]);
  assign t[345] = (x[34]);
  assign t[346] = (x[34]);
  assign t[347] = (x[37]);
  assign t[348] = (x[37]);
  assign t[349] = (x[40]);
  assign t[34] = ~t[53];
  assign t[350] = (x[40]);
  assign t[351] = (x[43]);
  assign t[352] = (x[43]);
  assign t[353] = (x[46]);
  assign t[354] = (x[46]);
  assign t[355] = (x[49]);
  assign t[356] = (x[49]);
  assign t[357] = (x[52]);
  assign t[358] = (x[52]);
  assign t[359] = (x[59]);
  assign t[35] = ~(t[54]);
  assign t[360] = (x[59]);
  assign t[361] = (x[62]);
  assign t[362] = (x[62]);
  assign t[363] = (x[65]);
  assign t[364] = (x[65]);
  assign t[365] = (x[68]);
  assign t[366] = (x[68]);
  assign t[367] = (x[77]);
  assign t[368] = (x[77]);
  assign t[369] = (x[80]);
  assign t[36] = t[55];
  assign t[370] = (x[80]);
  assign t[371] = (x[83]);
  assign t[372] = (x[83]);
  assign t[373] = (x[86]);
  assign t[374] = (x[86]);
  assign t[375] = (x[91]);
  assign t[376] = (x[91]);
  assign t[377] = (x[104]);
  assign t[378] = (x[104]);
  assign t[37] = ~(t[56] ^ t[57]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[41] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[61] : t[194];
  assign t[41] = t[8] ? t[62] : t[195];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[65] & t[66];
  assign t[44] = t[13] ^ t[67];
  assign t[45] = t[68] ^ t[69];
  assign t[46] = t[54] ^ t[34];
  assign t[47] = t[70] ^ t[71];
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = t[196] | t[74];
  assign t[4] = t[8] ? t[9] : t[190];
  assign t[50] = ~(t[197]);
  assign t[51] = ~(t[75] & t[198]);
  assign t[52] = t[8] ? t[76] : t[199];
  assign t[53] = t[8] ? t[77] : t[200];
  assign t[54] = ~t[78];
  assign t[55] = t[27] ? t[79] : t[201];
  assign t[56] = t[80] ^ t[81];
  assign t[57] = ~(t[82] ^ t[83]);
  assign t[58] = t[84] ^ t[85];
  assign t[59] = t[86] & t[87];
  assign t[5] = ~(t[10]);
  assign t[60] = t[42] ^ t[88];
  assign t[61] = t[194] ^ t[89];
  assign t[62] = t[195] ^ t[90];
  assign t[63] = t[91] & t[92];
  assign t[64] = t[93] & t[94];
  assign t[65] = ~(t[63] ^ t[95]);
  assign t[66] = t[96] ^ t[97];
  assign t[67] = t[98] ^ t[99];
  assign t[68] = t[100] ^ t[101];
  assign t[69] = t[102] & t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[104] ^ t[20];
  assign t[71] = t[105] & t[106];
  assign t[72] = ~(t[74] & t[107]);
  assign t[73] = ~(t[202] ^ t[108]);
  assign t[74] = ~(t[109] & t[110]);
  assign t[75] = ~(t[203]);
  assign t[76] = t[199] ^ t[111];
  assign t[77] = t[200] ^ t[112];
  assign t[78] = t[8] ? t[113] : t[204];
  assign t[79] = t[201] ^ t[114];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[115] ^ t[116];
  assign t[81] = t[117] ^ t[118];
  assign t[82] = t[119] ^ t[120];
  assign t[83] = t[121] ^ t[122];
  assign t[84] = t[27] ? t[123] : t[205];
  assign t[85] = t[27] ? t[124] : t[206];
  assign t[86] = ~(t[58] ^ t[125]);
  assign t[87] = t[126] ^ t[127];
  assign t[88] = t[128] & t[129];
  assign t[89] = t[130] ? x[56] : x[55];
  assign t[8] = ~(t[15]);
  assign t[90] = t[130] ? x[58] : x[57];
  assign t[91] = ~(t[97]);
  assign t[92] = ~(t[131]);
  assign t[93] = ~(t[40]);
  assign t[94] = t[8] ? t[132] : t[207];
  assign t[95] = t[23] ^ t[131];
  assign t[96] = t[131] ^ t[41];
  assign t[97] = t[94] ^ t[40];
  assign t[98] = t[27] ? t[133] : t[208];
  assign t[99] = t[125] ^ t[59];
  assign t[9] = t[190] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [116:0] x;
 output y;

 wire [378:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[134] ? t[135] : t[209];
  assign t[101] = t[191] ^ t[136];
  assign t[102] = ~(t[68] ^ t[137]);
  assign t[103] = t[138] ^ t[139];
  assign t[104] = t[140] & t[141];
  assign t[105] = ~(t[104] ^ t[142]);
  assign t[106] = t[19] ^ t[143];
  assign t[107] = ~(t[144] & t[145]);
  assign t[108] = t[146] ^ t[210];
  assign t[109] = ~(t[202]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[147] & t[146];
  assign t[111] = t[130] ? x[72] : x[71];
  assign t[112] = t[130] ? x[74] : x[73];
  assign t[113] = t[204] ^ t[148];
  assign t[114] = t[130] ? x[76] : x[75];
  assign t[115] = t[100] ^ t[121];
  assign t[116] = t[149] & t[139];
  assign t[117] = t[33] ^ t[54];
  assign t[118] = t[150] & t[151];
  assign t[119] = t[126] ^ t[152];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[153] ^ t[88];
  assign t[121] = t[198] ^ t[154];
  assign t[122] = t[137] ^ t[69];
  assign t[123] = t[205] ^ t[155];
  assign t[124] = t[206] ^ t[156];
  assign t[125] = t[157] ^ t[158];
  assign t[126] = t[85] ^ t[98];
  assign t[127] = t[27] ? t[159] : t[211];
  assign t[128] = ~(t[153] ^ t[42]);
  assign t[129] = t[23] ^ t[94];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = ~(t[160]);
  assign t[131] = t[8] ? t[161] : t[212];
  assign t[132] = t[207] ^ t[162];
  assign t[133] = t[208] ^ t[163];
  assign t[134] = ~(t[15]);
  assign t[135] = t[209] ^ t[164];
  assign t[136] = t[134] ? t[165] : t[213];
  assign t[137] = t[166] ^ t[116];
  assign t[138] = t[101] ^ t[121];
  assign t[139] = t[192] ^ t[167];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[143]);
  assign t[141] = ~(t[33]);
  assign t[142] = t[46] ^ t[33];
  assign t[143] = t[36] ^ t[54];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[168] | t[109]);
  assign t[146] = ~(t[214]);
  assign t[147] = ~(t[210]);
  assign t[148] = t[130] ? x[90] : x[89];
  assign t[149] = ~(t[101]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[117] ^ t[70]);
  assign t[151] = t[46] ^ t[36];
  assign t[152] = t[125] ^ t[169];
  assign t[153] = t[131] ^ t[40];
  assign t[154] = t[134] ? t[170] : t[215];
  assign t[155] = t[171] ? x[95] : x[94];
  assign t[156] = t[171] ? x[97] : x[96];
  assign t[157] = t[172] & t[173];
  assign t[158] = t[174] & t[127];
  assign t[159] = t[211] ^ t[175];
  assign t[15] = ~(t[27]);
  assign t[160] = ~(t[28]);
  assign t[161] = t[212] ^ t[176];
  assign t[162] = t[130] ? x[99] : x[98];
  assign t[163] = t[28] ? x[101] : x[100];
  assign t[164] = t[177] ? x[103] : x[102];
  assign t[165] = t[213] ^ t[178];
  assign t[166] = t[179] & t[180];
  assign t[167] = t[134] ? t[181] : t[216];
  assign t[168] = ~(t[196]);
  assign t[169] = t[182] & t[183];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[215] ^ t[184];
  assign t[171] = ~(t[160]);
  assign t[172] = ~(t[185]);
  assign t[173] = ~(t[84]);
  assign t[174] = ~(t[85]);
  assign t[175] = t[28] ? x[108] : x[107];
  assign t[176] = t[130] ? x[110] : x[109];
  assign t[177] = ~(t[160]);
  assign t[178] = t[177] ? x[112] : x[111];
  assign t[179] = ~(t[186]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[100]);
  assign t[181] = t[216] ^ t[187];
  assign t[182] = ~(t[157] ^ t[188]);
  assign t[183] = t[189] ^ t[185];
  assign t[184] = t[177] ? x[114] : x[113];
  assign t[185] = t[127] ^ t[85];
  assign t[186] = t[139] ^ t[101];
  assign t[187] = t[177] ? x[116] : x[115];
  assign t[188] = t[126] ^ t[84];
  assign t[189] = t[84] ^ t[98];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] & t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = t[244] ^ x[4];
  assign t[218] = t[245] ^ x[9];
  assign t[219] = t[246] ^ x[12];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[15];
  assign t[221] = t[248] ^ x[18];
  assign t[222] = t[249] ^ x[21];
  assign t[223] = t[250] ^ x[24];
  assign t[224] = t[251] ^ x[27];
  assign t[225] = t[252] ^ x[30];
  assign t[226] = t[253] ^ x[33];
  assign t[227] = t[254] ^ x[36];
  assign t[228] = t[255] ^ x[39];
  assign t[229] = t[256] ^ x[42];
  assign t[22] = ~(t[26] ^ t[39]);
  assign t[230] = t[257] ^ x[45];
  assign t[231] = t[258] ^ x[48];
  assign t[232] = t[259] ^ x[51];
  assign t[233] = t[260] ^ x[54];
  assign t[234] = t[261] ^ x[61];
  assign t[235] = t[262] ^ x[64];
  assign t[236] = t[263] ^ x[67];
  assign t[237] = t[264] ^ x[70];
  assign t[238] = t[265] ^ x[79];
  assign t[239] = t[266] ^ x[82];
  assign t[23] = t[40] ^ t[41];
  assign t[240] = t[267] ^ x[85];
  assign t[241] = t[268] ^ x[88];
  assign t[242] = t[269] ^ x[93];
  assign t[243] = t[270] ^ x[106];
  assign t[244] = (t[271] & ~t[272]);
  assign t[245] = (t[273] & ~t[274]);
  assign t[246] = (t[275] & ~t[276]);
  assign t[247] = (t[277] & ~t[278]);
  assign t[248] = (t[279] & ~t[280]);
  assign t[249] = (t[281] & ~t[282]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[283] & ~t[284]);
  assign t[251] = (t[285] & ~t[286]);
  assign t[252] = (t[287] & ~t[288]);
  assign t[253] = (t[289] & ~t[290]);
  assign t[254] = (t[291] & ~t[292]);
  assign t[255] = (t[293] & ~t[294]);
  assign t[256] = (t[295] & ~t[296]);
  assign t[257] = (t[297] & ~t[298]);
  assign t[258] = (t[299] & ~t[300]);
  assign t[259] = (t[301] & ~t[302]);
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[260] = (t[303] & ~t[304]);
  assign t[261] = (t[305] & ~t[306]);
  assign t[262] = (t[307] & ~t[308]);
  assign t[263] = (t[309] & ~t[310]);
  assign t[264] = (t[311] & ~t[312]);
  assign t[265] = (t[313] & ~t[314]);
  assign t[266] = (t[315] & ~t[316]);
  assign t[267] = (t[317] & ~t[318]);
  assign t[268] = (t[319] & ~t[320]);
  assign t[269] = (t[321] & ~t[322]);
  assign t[26] = t[46] ^ t[47];
  assign t[270] = (t[323] & ~t[324]);
  assign t[271] = t[325] ^ x[4];
  assign t[272] = t[326] ^ x[3];
  assign t[273] = t[327] ^ x[9];
  assign t[274] = t[328] ^ x[8];
  assign t[275] = t[329] ^ x[12];
  assign t[276] = t[330] ^ x[11];
  assign t[277] = t[331] ^ x[15];
  assign t[278] = t[332] ^ x[14];
  assign t[279] = t[333] ^ x[18];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[17];
  assign t[281] = t[335] ^ x[21];
  assign t[282] = t[336] ^ x[20];
  assign t[283] = t[337] ^ x[24];
  assign t[284] = t[338] ^ x[23];
  assign t[285] = t[339] ^ x[27];
  assign t[286] = t[340] ^ x[26];
  assign t[287] = t[341] ^ x[30];
  assign t[288] = t[342] ^ x[29];
  assign t[289] = t[343] ^ x[33];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[32];
  assign t[291] = t[345] ^ x[36];
  assign t[292] = t[346] ^ x[35];
  assign t[293] = t[347] ^ x[39];
  assign t[294] = t[348] ^ x[38];
  assign t[295] = t[349] ^ x[42];
  assign t[296] = t[350] ^ x[41];
  assign t[297] = t[351] ^ x[45];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[48];
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[47];
  assign t[301] = t[355] ^ x[51];
  assign t[302] = t[356] ^ x[50];
  assign t[303] = t[357] ^ x[54];
  assign t[304] = t[358] ^ x[53];
  assign t[305] = t[359] ^ x[61];
  assign t[306] = t[360] ^ x[60];
  assign t[307] = t[361] ^ x[64];
  assign t[308] = t[362] ^ x[63];
  assign t[309] = t[363] ^ x[67];
  assign t[30] = ~(t[192]);
  assign t[310] = t[364] ^ x[66];
  assign t[311] = t[365] ^ x[70];
  assign t[312] = t[366] ^ x[69];
  assign t[313] = t[367] ^ x[79];
  assign t[314] = t[368] ^ x[78];
  assign t[315] = t[369] ^ x[82];
  assign t[316] = t[370] ^ x[81];
  assign t[317] = t[371] ^ x[85];
  assign t[318] = t[372] ^ x[84];
  assign t[319] = t[373] ^ x[88];
  assign t[31] = ~(t[193]);
  assign t[320] = t[374] ^ x[87];
  assign t[321] = t[375] ^ x[93];
  assign t[322] = t[376] ^ x[92];
  assign t[323] = t[377] ^ x[106];
  assign t[324] = t[378] ^ x[105];
  assign t[325] = (x[2]);
  assign t[326] = (x[2]);
  assign t[327] = (x[7]);
  assign t[328] = (x[7]);
  assign t[329] = (x[10]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (x[10]);
  assign t[331] = (x[13]);
  assign t[332] = (x[13]);
  assign t[333] = (x[16]);
  assign t[334] = (x[16]);
  assign t[335] = (x[19]);
  assign t[336] = (x[19]);
  assign t[337] = (x[22]);
  assign t[338] = (x[22]);
  assign t[339] = (x[25]);
  assign t[33] = t[52];
  assign t[340] = (x[25]);
  assign t[341] = (x[28]);
  assign t[342] = (x[28]);
  assign t[343] = (x[31]);
  assign t[344] = (x[31]);
  assign t[345] = (x[34]);
  assign t[346] = (x[34]);
  assign t[347] = (x[37]);
  assign t[348] = (x[37]);
  assign t[349] = (x[40]);
  assign t[34] = ~t[53];
  assign t[350] = (x[40]);
  assign t[351] = (x[43]);
  assign t[352] = (x[43]);
  assign t[353] = (x[46]);
  assign t[354] = (x[46]);
  assign t[355] = (x[49]);
  assign t[356] = (x[49]);
  assign t[357] = (x[52]);
  assign t[358] = (x[52]);
  assign t[359] = (x[59]);
  assign t[35] = ~(t[54]);
  assign t[360] = (x[59]);
  assign t[361] = (x[62]);
  assign t[362] = (x[62]);
  assign t[363] = (x[65]);
  assign t[364] = (x[65]);
  assign t[365] = (x[68]);
  assign t[366] = (x[68]);
  assign t[367] = (x[77]);
  assign t[368] = (x[77]);
  assign t[369] = (x[80]);
  assign t[36] = t[55];
  assign t[370] = (x[80]);
  assign t[371] = (x[83]);
  assign t[372] = (x[83]);
  assign t[373] = (x[86]);
  assign t[374] = (x[86]);
  assign t[375] = (x[91]);
  assign t[376] = (x[91]);
  assign t[377] = (x[104]);
  assign t[378] = (x[104]);
  assign t[37] = ~(t[56] ^ t[57]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[41] ^ t[60];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[61] : t[194];
  assign t[41] = t[8] ? t[62] : t[195];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[65] & t[66];
  assign t[44] = t[13] ^ t[67];
  assign t[45] = t[68] ^ t[69];
  assign t[46] = t[54] ^ t[34];
  assign t[47] = t[70] ^ t[71];
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = t[196] | t[74];
  assign t[4] = t[8] ? t[9] : t[190];
  assign t[50] = ~(t[197]);
  assign t[51] = ~(t[75] & t[198]);
  assign t[52] = t[8] ? t[76] : t[199];
  assign t[53] = t[8] ? t[77] : t[200];
  assign t[54] = ~t[78];
  assign t[55] = t[27] ? t[79] : t[201];
  assign t[56] = t[80] ^ t[81];
  assign t[57] = ~(t[82] ^ t[83]);
  assign t[58] = t[84] ^ t[85];
  assign t[59] = t[86] & t[87];
  assign t[5] = ~(t[10]);
  assign t[60] = t[42] ^ t[88];
  assign t[61] = t[194] ^ t[89];
  assign t[62] = t[195] ^ t[90];
  assign t[63] = t[91] & t[92];
  assign t[64] = t[93] & t[94];
  assign t[65] = ~(t[63] ^ t[95]);
  assign t[66] = t[96] ^ t[97];
  assign t[67] = t[98] ^ t[99];
  assign t[68] = t[100] ^ t[101];
  assign t[69] = t[102] & t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[104] ^ t[20];
  assign t[71] = t[105] & t[106];
  assign t[72] = ~(t[74] & t[107]);
  assign t[73] = ~(t[202] ^ t[108]);
  assign t[74] = ~(t[109] & t[110]);
  assign t[75] = ~(t[203]);
  assign t[76] = t[199] ^ t[111];
  assign t[77] = t[200] ^ t[112];
  assign t[78] = t[8] ? t[113] : t[204];
  assign t[79] = t[201] ^ t[114];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[115] ^ t[116];
  assign t[81] = t[117] ^ t[118];
  assign t[82] = t[119] ^ t[120];
  assign t[83] = t[121] ^ t[122];
  assign t[84] = t[27] ? t[123] : t[205];
  assign t[85] = t[27] ? t[124] : t[206];
  assign t[86] = ~(t[58] ^ t[125]);
  assign t[87] = t[126] ^ t[127];
  assign t[88] = t[128] & t[129];
  assign t[89] = t[130] ? x[56] : x[55];
  assign t[8] = ~(t[15]);
  assign t[90] = t[130] ? x[58] : x[57];
  assign t[91] = ~(t[97]);
  assign t[92] = ~(t[131]);
  assign t[93] = ~(t[40]);
  assign t[94] = t[8] ? t[132] : t[207];
  assign t[95] = t[23] ^ t[131];
  assign t[96] = t[131] ^ t[41];
  assign t[97] = t[94] ^ t[40];
  assign t[98] = t[27] ? t[133] : t[208];
  assign t[99] = t[125] ^ t[59];
  assign t[9] = t[190] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [116:0] x;
 output y;

 wire [396:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[8]);
  assign t[101] = t[31] ? x[50] : x[49];
  assign t[102] = ~(t[137] ^ t[65]);
  assign t[103] = t[40] ^ t[106];
  assign t[104] = t[67] ? t[138] : t[223];
  assign t[105] = ~(t[64]);
  assign t[106] = t[67] ? t[139] : t[224];
  assign t[107] = t[8] ? t[140] : t[225];
  assign t[108] = t[8] ? t[141] : t[226];
  assign t[109] = t[142] ^ t[126];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[143] & t[144];
  assign t[111] = t[67] ? t[145] : t[227];
  assign t[112] = t[146] ^ t[147];
  assign t[113] = t[45] ^ t[148];
  assign t[114] = t[149] ^ t[150];
  assign t[115] = t[8] ? t[151] : t[228];
  assign t[116] = ~(t[78] ^ t[109]);
  assign t[117] = t[72] ^ t[152];
  assign t[118] = t[153] & t[154];
  assign t[119] = ~(t[209]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[108] ^ t[155];
  assign t[121] = t[156] ^ t[157];
  assign t[122] = t[158] & t[159];
  assign t[123] = t[157] ^ t[149];
  assign t[124] = t[160] ^ t[161];
  assign t[125] = t[115] ^ t[108];
  assign t[126] = t[162] & t[152];
  assign t[127] = t[221] ^ t[163];
  assign t[128] = t[222] ^ t[164];
  assign t[129] = t[165] & t[166];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[167] & t[95];
  assign t[131] = t[8] ? t[168] : t[229];
  assign t[132] = t[31] ? x[73] : x[72];
  assign t[133] = ~(t[136]);
  assign t[134] = ~(t[104]);
  assign t[135] = t[40] ^ t[104];
  assign t[136] = t[106] ^ t[64];
  assign t[137] = t[104] ^ t[64];
  assign t[138] = t[223] ^ t[169];
  assign t[139] = t[224] ^ t[170];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[225] ^ t[171];
  assign t[141] = t[226] ^ t[172];
  assign t[142] = t[173] & t[174];
  assign t[143] = ~(t[142] ^ t[175]);
  assign t[144] = t[125] ^ t[176];
  assign t[145] = t[227] ^ t[177];
  assign t[146] = t[156] ^ t[149];
  assign t[147] = t[178] & t[179];
  assign t[148] = t[137] ^ t[69];
  assign t[149] = t[217] ^ t[180];
  assign t[14] = ~(t[26] ^ t[27]);
  assign t[150] = t[160] ^ t[122];
  assign t[151] = t[228] ^ t[181];
  assign t[152] = t[8] ? t[182] : t[230];
  assign t[153] = ~(t[129] ^ t[183]);
  assign t[154] = t[184] ^ t[185];
  assign t[155] = t[109] ^ t[79];
  assign t[156] = t[186] ? t[187] : t[231];
  assign t[157] = t[211] ^ t[188];
  assign t[158] = ~(t[121] ^ t[160]);
  assign t[159] = t[123] ^ t[179];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[189] ^ t[147];
  assign t[161] = t[190] & t[191];
  assign t[162] = ~(t[107]);
  assign t[163] = t[31] ? x[81] : x[80];
  assign t[164] = t[31] ? x[83] : x[82];
  assign t[165] = ~(t[185]);
  assign t[166] = ~(t[60]);
  assign t[167] = ~(t[61]);
  assign t[168] = t[229] ^ t[192];
  assign t[169] = t[31] ? x[85] : x[84];
  assign t[16] = t[209] | t[30];
  assign t[170] = t[31] ? x[87] : x[86];
  assign t[171] = t[193] ? x[89] : x[88];
  assign t[172] = t[86] ? x[91] : x[90];
  assign t[173] = ~(t[176]);
  assign t[174] = ~(t[115]);
  assign t[175] = t[72] ^ t[115];
  assign t[176] = t[152] ^ t[107];
  assign t[177] = t[31] ? x[93] : x[92];
  assign t[178] = ~(t[157]);
  assign t[179] = t[212] ^ t[194];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[186] ? t[195] : t[232];
  assign t[181] = t[193] ? x[98] : x[97];
  assign t[182] = t[230] ^ t[196];
  assign t[183] = t[80] ^ t[60];
  assign t[184] = t[60] ^ t[74];
  assign t[185] = t[95] ^ t[61];
  assign t[186] = ~(t[100]);
  assign t[187] = t[231] ^ t[197];
  assign t[188] = t[186] ? t[198] : t[233];
  assign t[189] = t[199] & t[200];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = ~(t[189] ^ t[201]);
  assign t[191] = t[146] ^ t[202];
  assign t[192] = t[31] ? x[103] : x[102];
  assign t[193] = ~(t[54]);
  assign t[194] = t[186] ? t[203] : t[234];
  assign t[195] = t[232] ^ t[204];
  assign t[196] = t[86] ? x[108] : x[107];
  assign t[197] = t[205] ? x[110] : x[109];
  assign t[198] = t[233] ^ t[206];
  assign t[199] = ~(t[202]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[156]);
  assign t[201] = t[123] ^ t[156];
  assign t[202] = t[179] ^ t[157];
  assign t[203] = t[234] ^ t[207];
  assign t[204] = t[205] ? x[112] : x[111];
  assign t[205] = ~(t[54]);
  assign t[206] = t[205] ? x[114] : x[113];
  assign t[207] = t[205] ? x[116] : x[115];
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[36] ^ t[37];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = t[262] ^ x[4];
  assign t[236] = t[263] ^ x[7];
  assign t[237] = t[264] ^ x[12];
  assign t[238] = t[265] ^ x[15];
  assign t[239] = t[266] ^ x[18];
  assign t[23] = t[42] ^ t[43];
  assign t[240] = t[267] ^ x[21];
  assign t[241] = t[268] ^ x[24];
  assign t[242] = t[269] ^ x[27];
  assign t[243] = t[270] ^ x[30];
  assign t[244] = t[271] ^ x[33];
  assign t[245] = t[272] ^ x[36];
  assign t[246] = t[273] ^ x[39];
  assign t[247] = t[274] ^ x[42];
  assign t[248] = t[275] ^ x[45];
  assign t[249] = t[276] ^ x[48];
  assign t[24] = t[44] ^ t[45];
  assign t[250] = t[277] ^ x[53];
  assign t[251] = t[278] ^ x[56];
  assign t[252] = t[279] ^ x[59];
  assign t[253] = t[280] ^ x[62];
  assign t[254] = t[281] ^ x[65];
  assign t[255] = t[282] ^ x[68];
  assign t[256] = t[283] ^ x[71];
  assign t[257] = t[284] ^ x[76];
  assign t[258] = t[285] ^ x[79];
  assign t[259] = t[286] ^ x[96];
  assign t[25] = ~(t[36] ^ t[46]);
  assign t[260] = t[287] ^ x[101];
  assign t[261] = t[288] ^ x[106];
  assign t[262] = (t[289] & ~t[290]);
  assign t[263] = (t[291] & ~t[292]);
  assign t[264] = (t[293] & ~t[294]);
  assign t[265] = (t[295] & ~t[296]);
  assign t[266] = (t[297] & ~t[298]);
  assign t[267] = (t[299] & ~t[300]);
  assign t[268] = (t[301] & ~t[302]);
  assign t[269] = (t[303] & ~t[304]);
  assign t[26] = t[47] ^ t[48];
  assign t[270] = (t[305] & ~t[306]);
  assign t[271] = (t[307] & ~t[308]);
  assign t[272] = (t[309] & ~t[310]);
  assign t[273] = (t[311] & ~t[312]);
  assign t[274] = (t[313] & ~t[314]);
  assign t[275] = (t[315] & ~t[316]);
  assign t[276] = (t[317] & ~t[318]);
  assign t[277] = (t[319] & ~t[320]);
  assign t[278] = (t[321] & ~t[322]);
  assign t[279] = (t[323] & ~t[324]);
  assign t[27] = ~(t[49] ^ t[23]);
  assign t[280] = (t[325] & ~t[326]);
  assign t[281] = (t[327] & ~t[328]);
  assign t[282] = (t[329] & ~t[330]);
  assign t[283] = (t[331] & ~t[332]);
  assign t[284] = (t[333] & ~t[334]);
  assign t[285] = (t[335] & ~t[336]);
  assign t[286] = (t[337] & ~t[338]);
  assign t[287] = (t[339] & ~t[340]);
  assign t[288] = (t[341] & ~t[342]);
  assign t[289] = t[343] ^ x[4];
  assign t[28] = ~(t[30] & t[50]);
  assign t[290] = t[344] ^ x[3];
  assign t[291] = t[345] ^ x[7];
  assign t[292] = t[346] ^ x[6];
  assign t[293] = t[347] ^ x[12];
  assign t[294] = t[348] ^ x[11];
  assign t[295] = t[349] ^ x[15];
  assign t[296] = t[350] ^ x[14];
  assign t[297] = t[351] ^ x[18];
  assign t[298] = t[352] ^ x[17];
  assign t[299] = t[353] ^ x[21];
  assign t[29] = ~(t[210] ^ t[51]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[20];
  assign t[301] = t[355] ^ x[24];
  assign t[302] = t[356] ^ x[23];
  assign t[303] = t[357] ^ x[27];
  assign t[304] = t[358] ^ x[26];
  assign t[305] = t[359] ^ x[30];
  assign t[306] = t[360] ^ x[29];
  assign t[307] = t[361] ^ x[33];
  assign t[308] = t[362] ^ x[32];
  assign t[309] = t[363] ^ x[36];
  assign t[30] = ~(t[52] & t[53]);
  assign t[310] = t[364] ^ x[35];
  assign t[311] = t[365] ^ x[39];
  assign t[312] = t[366] ^ x[38];
  assign t[313] = t[367] ^ x[42];
  assign t[314] = t[368] ^ x[41];
  assign t[315] = t[369] ^ x[45];
  assign t[316] = t[370] ^ x[44];
  assign t[317] = t[371] ^ x[48];
  assign t[318] = t[372] ^ x[47];
  assign t[319] = t[373] ^ x[53];
  assign t[31] = ~(t[54]);
  assign t[320] = t[374] ^ x[52];
  assign t[321] = t[375] ^ x[56];
  assign t[322] = t[376] ^ x[55];
  assign t[323] = t[377] ^ x[59];
  assign t[324] = t[378] ^ x[58];
  assign t[325] = t[379] ^ x[62];
  assign t[326] = t[380] ^ x[61];
  assign t[327] = t[381] ^ x[65];
  assign t[328] = t[382] ^ x[64];
  assign t[329] = t[383] ^ x[68];
  assign t[32] = ~(t[211]);
  assign t[330] = t[384] ^ x[67];
  assign t[331] = t[385] ^ x[71];
  assign t[332] = t[386] ^ x[70];
  assign t[333] = t[387] ^ x[76];
  assign t[334] = t[388] ^ x[75];
  assign t[335] = t[389] ^ x[79];
  assign t[336] = t[390] ^ x[78];
  assign t[337] = t[391] ^ x[96];
  assign t[338] = t[392] ^ x[95];
  assign t[339] = t[393] ^ x[101];
  assign t[33] = ~(t[212]);
  assign t[340] = t[394] ^ x[100];
  assign t[341] = t[395] ^ x[106];
  assign t[342] = t[396] ^ x[105];
  assign t[343] = (x[2]);
  assign t[344] = (x[2]);
  assign t[345] = (x[5]);
  assign t[346] = (x[5]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[213]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = ~(t[57] ^ t[49]);
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[51]);
  assign t[374] = (x[51]);
  assign t[375] = (x[54]);
  assign t[376] = (x[54]);
  assign t[377] = (x[57]);
  assign t[378] = (x[57]);
  assign t[379] = (x[60]);
  assign t[37] = ~(t[58] ^ t[59]);
  assign t[380] = (x[60]);
  assign t[381] = (x[63]);
  assign t[382] = (x[63]);
  assign t[383] = (x[66]);
  assign t[384] = (x[66]);
  assign t[385] = (x[69]);
  assign t[386] = (x[69]);
  assign t[387] = (x[74]);
  assign t[388] = (x[74]);
  assign t[389] = (x[77]);
  assign t[38] = t[60] ^ t[61];
  assign t[390] = (x[77]);
  assign t[391] = (x[94]);
  assign t[392] = (x[94]);
  assign t[393] = (x[99]);
  assign t[394] = (x[99]);
  assign t[395] = (x[104]);
  assign t[396] = (x[104]);
  assign t[39] = t[62] & t[63];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[42];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] ? t[68] : t[214];
  assign t[43] = t[65] ^ t[69];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = ~(t[76] ^ t[77]);
  assign t[48] = t[78] ^ t[79];
  assign t[49] = t[80] ^ t[81];
  assign t[4] = t[8] ? t[9] : t[208];
  assign t[50] = ~(t[82] & t[83]);
  assign t[51] = t[84] ^ t[215];
  assign t[52] = ~(t[210]);
  assign t[53] = t[85] & t[84];
  assign t[54] = ~(t[86]);
  assign t[55] = ~(t[216]);
  assign t[56] = ~(t[87] & t[217]);
  assign t[57] = ~(t[88] ^ t[89]);
  assign t[58] = t[90] ^ t[91];
  assign t[59] = ~(t[46] ^ t[23]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[92];
  assign t[61] = ~t[93];
  assign t[62] = ~(t[38] ^ t[94]);
  assign t[63] = t[80] ^ t[95];
  assign t[64] = t[67] ? t[96] : t[218];
  assign t[65] = t[97] ^ t[71];
  assign t[66] = t[98] & t[99];
  assign t[67] = ~(t[100]);
  assign t[68] = t[214] ^ t[101];
  assign t[69] = t[102] & t[103];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[104] ^ t[42];
  assign t[71] = t[105] & t[106];
  assign t[72] = t[107] ^ t[108];
  assign t[73] = t[109] ^ t[110];
  assign t[74] = ~t[111];
  assign t[75] = t[94] ^ t[39];
  assign t[76] = t[112] ^ t[21];
  assign t[77] = ~(t[113] ^ t[114]);
  assign t[78] = t[115] ^ t[107];
  assign t[79] = t[116] & t[117];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[61] ^ t[74];
  assign t[81] = t[94] ^ t[118];
  assign t[82] = ~(t[85] | t[84]);
  assign t[83] = ~(t[119] | t[52]);
  assign t[84] = ~(t[219]);
  assign t[85] = ~(t[215]);
  assign t[86] = ~(t[16]);
  assign t[87] = ~(t[220]);
  assign t[88] = t[22] ^ t[120];
  assign t[89] = t[121] ^ t[122];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[123] ^ t[124];
  assign t[91] = t[125] ^ t[126];
  assign t[92] = t[67] ? t[127] : t[221];
  assign t[93] = t[67] ? t[128] : t[222];
  assign t[94] = t[129] ^ t[130];
  assign t[95] = t[131];
  assign t[96] = t[218] ^ t[132];
  assign t[97] = t[133] & t[134];
  assign t[98] = ~(t[97] ^ t[135]);
  assign t[99] = t[70] ^ t[136];
  assign t[9] = t[208] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [116:0] x;
 output y;

 wire [396:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[8]);
  assign t[101] = t[31] ? x[50] : x[49];
  assign t[102] = ~(t[137] ^ t[65]);
  assign t[103] = t[40] ^ t[106];
  assign t[104] = t[67] ? t[138] : t[223];
  assign t[105] = ~(t[64]);
  assign t[106] = t[67] ? t[139] : t[224];
  assign t[107] = t[8] ? t[140] : t[225];
  assign t[108] = t[8] ? t[141] : t[226];
  assign t[109] = t[142] ^ t[126];
  assign t[10] = ~(t[18] | t[19]);
  assign t[110] = t[143] & t[144];
  assign t[111] = t[67] ? t[145] : t[227];
  assign t[112] = t[146] ^ t[147];
  assign t[113] = t[45] ^ t[148];
  assign t[114] = t[149] ^ t[150];
  assign t[115] = t[8] ? t[151] : t[228];
  assign t[116] = ~(t[78] ^ t[109]);
  assign t[117] = t[72] ^ t[152];
  assign t[118] = t[153] & t[154];
  assign t[119] = ~(t[209]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[108] ^ t[155];
  assign t[121] = t[156] ^ t[157];
  assign t[122] = t[158] & t[159];
  assign t[123] = t[157] ^ t[149];
  assign t[124] = t[160] ^ t[161];
  assign t[125] = t[115] ^ t[108];
  assign t[126] = t[162] & t[152];
  assign t[127] = t[221] ^ t[163];
  assign t[128] = t[222] ^ t[164];
  assign t[129] = t[165] & t[166];
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[130] = t[167] & t[95];
  assign t[131] = t[8] ? t[168] : t[229];
  assign t[132] = t[31] ? x[73] : x[72];
  assign t[133] = ~(t[136]);
  assign t[134] = ~(t[104]);
  assign t[135] = t[40] ^ t[104];
  assign t[136] = t[106] ^ t[64];
  assign t[137] = t[104] ^ t[64];
  assign t[138] = t[223] ^ t[169];
  assign t[139] = t[224] ^ t[170];
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[140] = t[225] ^ t[171];
  assign t[141] = t[226] ^ t[172];
  assign t[142] = t[173] & t[174];
  assign t[143] = ~(t[142] ^ t[175]);
  assign t[144] = t[125] ^ t[176];
  assign t[145] = t[227] ^ t[177];
  assign t[146] = t[156] ^ t[149];
  assign t[147] = t[178] & t[179];
  assign t[148] = t[137] ^ t[69];
  assign t[149] = t[217] ^ t[180];
  assign t[14] = ~(t[26] ^ t[27]);
  assign t[150] = t[160] ^ t[122];
  assign t[151] = t[228] ^ t[181];
  assign t[152] = t[8] ? t[182] : t[230];
  assign t[153] = ~(t[129] ^ t[183]);
  assign t[154] = t[184] ^ t[185];
  assign t[155] = t[109] ^ t[79];
  assign t[156] = t[186] ? t[187] : t[231];
  assign t[157] = t[211] ^ t[188];
  assign t[158] = ~(t[121] ^ t[160]);
  assign t[159] = t[123] ^ t[179];
  assign t[15] = ~(t[28] & t[29]);
  assign t[160] = t[189] ^ t[147];
  assign t[161] = t[190] & t[191];
  assign t[162] = ~(t[107]);
  assign t[163] = t[31] ? x[81] : x[80];
  assign t[164] = t[31] ? x[83] : x[82];
  assign t[165] = ~(t[185]);
  assign t[166] = ~(t[60]);
  assign t[167] = ~(t[61]);
  assign t[168] = t[229] ^ t[192];
  assign t[169] = t[31] ? x[85] : x[84];
  assign t[16] = t[209] | t[30];
  assign t[170] = t[31] ? x[87] : x[86];
  assign t[171] = t[193] ? x[89] : x[88];
  assign t[172] = t[86] ? x[91] : x[90];
  assign t[173] = ~(t[176]);
  assign t[174] = ~(t[115]);
  assign t[175] = t[72] ^ t[115];
  assign t[176] = t[152] ^ t[107];
  assign t[177] = t[31] ? x[93] : x[92];
  assign t[178] = ~(t[157]);
  assign t[179] = t[212] ^ t[194];
  assign t[17] = t[31] ? x[9] : x[8];
  assign t[180] = t[186] ? t[195] : t[232];
  assign t[181] = t[193] ? x[98] : x[97];
  assign t[182] = t[230] ^ t[196];
  assign t[183] = t[80] ^ t[60];
  assign t[184] = t[60] ^ t[74];
  assign t[185] = t[95] ^ t[61];
  assign t[186] = ~(t[100]);
  assign t[187] = t[231] ^ t[197];
  assign t[188] = t[186] ? t[198] : t[233];
  assign t[189] = t[199] & t[200];
  assign t[18] = ~(t[32] & t[33]);
  assign t[190] = ~(t[189] ^ t[201]);
  assign t[191] = t[146] ^ t[202];
  assign t[192] = t[31] ? x[103] : x[102];
  assign t[193] = ~(t[54]);
  assign t[194] = t[186] ? t[203] : t[234];
  assign t[195] = t[232] ^ t[204];
  assign t[196] = t[86] ? x[108] : x[107];
  assign t[197] = t[205] ? x[110] : x[109];
  assign t[198] = t[233] ^ t[206];
  assign t[199] = ~(t[202]);
  assign t[19] = ~(t[34] & t[35]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[156]);
  assign t[201] = t[123] ^ t[156];
  assign t[202] = t[179] ^ t[157];
  assign t[203] = t[234] ^ t[207];
  assign t[204] = t[205] ? x[112] : x[111];
  assign t[205] = ~(t[54]);
  assign t[206] = t[205] ? x[114] : x[113];
  assign t[207] = t[205] ? x[116] : x[115];
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[36] ^ t[37];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[38] ^ t[39];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[40] ^ t[41];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = t[262] ^ x[4];
  assign t[236] = t[263] ^ x[7];
  assign t[237] = t[264] ^ x[12];
  assign t[238] = t[265] ^ x[15];
  assign t[239] = t[266] ^ x[18];
  assign t[23] = t[42] ^ t[43];
  assign t[240] = t[267] ^ x[21];
  assign t[241] = t[268] ^ x[24];
  assign t[242] = t[269] ^ x[27];
  assign t[243] = t[270] ^ x[30];
  assign t[244] = t[271] ^ x[33];
  assign t[245] = t[272] ^ x[36];
  assign t[246] = t[273] ^ x[39];
  assign t[247] = t[274] ^ x[42];
  assign t[248] = t[275] ^ x[45];
  assign t[249] = t[276] ^ x[48];
  assign t[24] = t[44] ^ t[45];
  assign t[250] = t[277] ^ x[53];
  assign t[251] = t[278] ^ x[56];
  assign t[252] = t[279] ^ x[59];
  assign t[253] = t[280] ^ x[62];
  assign t[254] = t[281] ^ x[65];
  assign t[255] = t[282] ^ x[68];
  assign t[256] = t[283] ^ x[71];
  assign t[257] = t[284] ^ x[76];
  assign t[258] = t[285] ^ x[79];
  assign t[259] = t[286] ^ x[96];
  assign t[25] = ~(t[36] ^ t[46]);
  assign t[260] = t[287] ^ x[101];
  assign t[261] = t[288] ^ x[106];
  assign t[262] = (t[289] & ~t[290]);
  assign t[263] = (t[291] & ~t[292]);
  assign t[264] = (t[293] & ~t[294]);
  assign t[265] = (t[295] & ~t[296]);
  assign t[266] = (t[297] & ~t[298]);
  assign t[267] = (t[299] & ~t[300]);
  assign t[268] = (t[301] & ~t[302]);
  assign t[269] = (t[303] & ~t[304]);
  assign t[26] = t[47] ^ t[48];
  assign t[270] = (t[305] & ~t[306]);
  assign t[271] = (t[307] & ~t[308]);
  assign t[272] = (t[309] & ~t[310]);
  assign t[273] = (t[311] & ~t[312]);
  assign t[274] = (t[313] & ~t[314]);
  assign t[275] = (t[315] & ~t[316]);
  assign t[276] = (t[317] & ~t[318]);
  assign t[277] = (t[319] & ~t[320]);
  assign t[278] = (t[321] & ~t[322]);
  assign t[279] = (t[323] & ~t[324]);
  assign t[27] = ~(t[49] ^ t[23]);
  assign t[280] = (t[325] & ~t[326]);
  assign t[281] = (t[327] & ~t[328]);
  assign t[282] = (t[329] & ~t[330]);
  assign t[283] = (t[331] & ~t[332]);
  assign t[284] = (t[333] & ~t[334]);
  assign t[285] = (t[335] & ~t[336]);
  assign t[286] = (t[337] & ~t[338]);
  assign t[287] = (t[339] & ~t[340]);
  assign t[288] = (t[341] & ~t[342]);
  assign t[289] = t[343] ^ x[4];
  assign t[28] = ~(t[30] & t[50]);
  assign t[290] = t[344] ^ x[3];
  assign t[291] = t[345] ^ x[7];
  assign t[292] = t[346] ^ x[6];
  assign t[293] = t[347] ^ x[12];
  assign t[294] = t[348] ^ x[11];
  assign t[295] = t[349] ^ x[15];
  assign t[296] = t[350] ^ x[14];
  assign t[297] = t[351] ^ x[18];
  assign t[298] = t[352] ^ x[17];
  assign t[299] = t[353] ^ x[21];
  assign t[29] = ~(t[210] ^ t[51]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[20];
  assign t[301] = t[355] ^ x[24];
  assign t[302] = t[356] ^ x[23];
  assign t[303] = t[357] ^ x[27];
  assign t[304] = t[358] ^ x[26];
  assign t[305] = t[359] ^ x[30];
  assign t[306] = t[360] ^ x[29];
  assign t[307] = t[361] ^ x[33];
  assign t[308] = t[362] ^ x[32];
  assign t[309] = t[363] ^ x[36];
  assign t[30] = ~(t[52] & t[53]);
  assign t[310] = t[364] ^ x[35];
  assign t[311] = t[365] ^ x[39];
  assign t[312] = t[366] ^ x[38];
  assign t[313] = t[367] ^ x[42];
  assign t[314] = t[368] ^ x[41];
  assign t[315] = t[369] ^ x[45];
  assign t[316] = t[370] ^ x[44];
  assign t[317] = t[371] ^ x[48];
  assign t[318] = t[372] ^ x[47];
  assign t[319] = t[373] ^ x[53];
  assign t[31] = ~(t[54]);
  assign t[320] = t[374] ^ x[52];
  assign t[321] = t[375] ^ x[56];
  assign t[322] = t[376] ^ x[55];
  assign t[323] = t[377] ^ x[59];
  assign t[324] = t[378] ^ x[58];
  assign t[325] = t[379] ^ x[62];
  assign t[326] = t[380] ^ x[61];
  assign t[327] = t[381] ^ x[65];
  assign t[328] = t[382] ^ x[64];
  assign t[329] = t[383] ^ x[68];
  assign t[32] = ~(t[211]);
  assign t[330] = t[384] ^ x[67];
  assign t[331] = t[385] ^ x[71];
  assign t[332] = t[386] ^ x[70];
  assign t[333] = t[387] ^ x[76];
  assign t[334] = t[388] ^ x[75];
  assign t[335] = t[389] ^ x[79];
  assign t[336] = t[390] ^ x[78];
  assign t[337] = t[391] ^ x[96];
  assign t[338] = t[392] ^ x[95];
  assign t[339] = t[393] ^ x[101];
  assign t[33] = ~(t[212]);
  assign t[340] = t[394] ^ x[100];
  assign t[341] = t[395] ^ x[106];
  assign t[342] = t[396] ^ x[105];
  assign t[343] = (x[2]);
  assign t[344] = (x[2]);
  assign t[345] = (x[5]);
  assign t[346] = (x[5]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[213]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = ~(t[57] ^ t[49]);
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[51]);
  assign t[374] = (x[51]);
  assign t[375] = (x[54]);
  assign t[376] = (x[54]);
  assign t[377] = (x[57]);
  assign t[378] = (x[57]);
  assign t[379] = (x[60]);
  assign t[37] = ~(t[58] ^ t[59]);
  assign t[380] = (x[60]);
  assign t[381] = (x[63]);
  assign t[382] = (x[63]);
  assign t[383] = (x[66]);
  assign t[384] = (x[66]);
  assign t[385] = (x[69]);
  assign t[386] = (x[69]);
  assign t[387] = (x[74]);
  assign t[388] = (x[74]);
  assign t[389] = (x[77]);
  assign t[38] = t[60] ^ t[61];
  assign t[390] = (x[77]);
  assign t[391] = (x[94]);
  assign t[392] = (x[94]);
  assign t[393] = (x[99]);
  assign t[394] = (x[99]);
  assign t[395] = (x[104]);
  assign t[396] = (x[104]);
  assign t[39] = t[62] & t[63];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[42];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] ? t[68] : t[214];
  assign t[43] = t[65] ^ t[69];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = ~(t[76] ^ t[77]);
  assign t[48] = t[78] ^ t[79];
  assign t[49] = t[80] ^ t[81];
  assign t[4] = t[8] ? t[9] : t[208];
  assign t[50] = ~(t[82] & t[83]);
  assign t[51] = t[84] ^ t[215];
  assign t[52] = ~(t[210]);
  assign t[53] = t[85] & t[84];
  assign t[54] = ~(t[86]);
  assign t[55] = ~(t[216]);
  assign t[56] = ~(t[87] & t[217]);
  assign t[57] = ~(t[88] ^ t[89]);
  assign t[58] = t[90] ^ t[91];
  assign t[59] = ~(t[46] ^ t[23]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[92];
  assign t[61] = ~t[93];
  assign t[62] = ~(t[38] ^ t[94]);
  assign t[63] = t[80] ^ t[95];
  assign t[64] = t[67] ? t[96] : t[218];
  assign t[65] = t[97] ^ t[71];
  assign t[66] = t[98] & t[99];
  assign t[67] = ~(t[100]);
  assign t[68] = t[214] ^ t[101];
  assign t[69] = t[102] & t[103];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[104] ^ t[42];
  assign t[71] = t[105] & t[106];
  assign t[72] = t[107] ^ t[108];
  assign t[73] = t[109] ^ t[110];
  assign t[74] = ~t[111];
  assign t[75] = t[94] ^ t[39];
  assign t[76] = t[112] ^ t[21];
  assign t[77] = ~(t[113] ^ t[114]);
  assign t[78] = t[115] ^ t[107];
  assign t[79] = t[116] & t[117];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[61] ^ t[74];
  assign t[81] = t[94] ^ t[118];
  assign t[82] = ~(t[85] | t[84]);
  assign t[83] = ~(t[119] | t[52]);
  assign t[84] = ~(t[219]);
  assign t[85] = ~(t[215]);
  assign t[86] = ~(t[16]);
  assign t[87] = ~(t[220]);
  assign t[88] = t[22] ^ t[120];
  assign t[89] = t[121] ^ t[122];
  assign t[8] = ~(t[15] & t[16]);
  assign t[90] = t[123] ^ t[124];
  assign t[91] = t[125] ^ t[126];
  assign t[92] = t[67] ? t[127] : t[221];
  assign t[93] = t[67] ? t[128] : t[222];
  assign t[94] = t[129] ^ t[130];
  assign t[95] = t[131];
  assign t[96] = t[218] ^ t[132];
  assign t[97] = t[133] & t[134];
  assign t[98] = ~(t[97] ^ t[135]);
  assign t[99] = t[70] ^ t[136];
  assign t[9] = t[208] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[98] ^ t[136]);
  assign t[101] = t[137] ^ t[138];
  assign t[102] = t[80] ? x[53] : x[52];
  assign t[103] = t[139] & t[140];
  assign t[104] = t[141] & t[126];
  assign t[105] = t[142] & t[143];
  assign t[106] = t[8] ? t[144] : t[213];
  assign t[107] = t[8] ? t[145] : t[214];
  assign t[108] = ~(t[70] ^ t[146]);
  assign t[109] = t[147] ^ t[148];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[147] ^ t[149];
  assign t[111] = t[150] ^ t[63];
  assign t[112] = t[91] ^ t[41];
  assign t[113] = t[35] ^ t[151];
  assign t[114] = t[8] ? t[152] : t[215];
  assign t[115] = t[146] ^ t[71];
  assign t[116] = ~(t[153] & t[154]);
  assign t[117] = t[155] ^ t[216];
  assign t[118] = ~(t[207]);
  assign t[119] = t[156] & t[155];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[28] ? x[67] : x[66];
  assign t[121] = t[28] ? x[69] : x[68];
  assign t[122] = t[157];
  assign t[123] = t[27] ? t[158] : t[217];
  assign t[124] = t[209] ^ t[159];
  assign t[125] = t[210] ^ t[160];
  assign t[126] = t[27] ? t[161] : t[218];
  assign t[127] = ~(t[15]);
  assign t[128] = t[211] ^ t[162];
  assign t[129] = ~(t[111] ^ t[64]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[39] ^ t[135];
  assign t[131] = t[212] ^ t[163];
  assign t[132] = ~(t[138]);
  assign t[133] = ~(t[150]);
  assign t[134] = ~(t[63]);
  assign t[135] = t[199] ^ t[164];
  assign t[136] = t[39] ^ t[150];
  assign t[137] = t[150] ^ t[61];
  assign t[138] = t[135] ^ t[63];
  assign t[139] = ~(t[165]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = ~(t[91]);
  assign t[141] = ~(t[92]);
  assign t[142] = ~(t[103] ^ t[166]);
  assign t[143] = t[112] ^ t[165];
  assign t[144] = t[213] ^ t[167];
  assign t[145] = t[214] ^ t[168];
  assign t[146] = t[169] ^ t[170];
  assign t[147] = t[107] ^ t[114];
  assign t[148] = t[8] ? t[171] : t[219];
  assign t[149] = t[146] ^ t[172];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[127] ? t[173] : t[220];
  assign t[151] = t[174] & t[175];
  assign t[152] = t[215] ^ t[176];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[177] | t[118]);
  assign t[155] = ~(t[221]);
  assign t[156] = ~(t[216]);
  assign t[157] = t[8] ? t[178] : t[222];
  assign t[158] = t[217] ^ t[179];
  assign t[159] = t[180] ? x[89] : x[88];
  assign t[15] = ~(t[27]);
  assign t[160] = t[180] ? x[91] : x[90];
  assign t[161] = t[218] ^ t[181];
  assign t[162] = t[182] ? x[93] : x[92];
  assign t[163] = t[182] ? x[95] : x[94];
  assign t[164] = t[127] ? t[183] : t[223];
  assign t[165] = t[126] ^ t[92];
  assign t[166] = t[68] ^ t[91];
  assign t[167] = t[28] ? x[100] : x[99];
  assign t[168] = t[28] ? x[102] : x[101];
  assign t[169] = t[184] & t[185];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[186] & t[148];
  assign t[171] = t[219] ^ t[187];
  assign t[172] = t[188] & t[189];
  assign t[173] = t[220] ^ t[190];
  assign t[174] = ~(t[191] ^ t[35]);
  assign t[175] = t[19] ^ t[87];
  assign t[176] = t[28] ? x[104] : x[103];
  assign t[177] = ~(t[202]);
  assign t[178] = t[222] ^ t[192];
  assign t[179] = t[28] ? x[106] : x[105];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[50]);
  assign t[181] = t[80] ? x[108] : x[107];
  assign t[182] = ~(t[50]);
  assign t[183] = t[223] ^ t[193];
  assign t[184] = ~(t[194]);
  assign t[185] = ~(t[106]);
  assign t[186] = ~(t[107]);
  assign t[187] = t[28] ? x[110] : x[109];
  assign t[188] = ~(t[169] ^ t[195]);
  assign t[189] = t[196] ^ t[194];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[182] ? x[112] : x[111];
  assign t[191] = t[122] ^ t[33];
  assign t[192] = t[28] ? x[114] : x[113];
  assign t[193] = t[182] ? x[116] : x[115];
  assign t[194] = t[148] ^ t[107];
  assign t[195] = t[147] ^ t[106];
  assign t[196] = t[106] ^ t[114];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = t[39] ^ t[40];
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[36];
  assign t[235] = t[262] ^ x[39];
  assign t[236] = t[263] ^ x[42];
  assign t[237] = t[264] ^ x[45];
  assign t[238] = t[265] ^ x[48];
  assign t[239] = t[266] ^ x[51];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[56];
  assign t[241] = t[268] ^ x[59];
  assign t[242] = t[269] ^ x[62];
  assign t[243] = t[270] ^ x[65];
  assign t[244] = t[271] ^ x[72];
  assign t[245] = t[272] ^ x[75];
  assign t[246] = t[273] ^ x[78];
  assign t[247] = t[274] ^ x[81];
  assign t[248] = t[275] ^ x[84];
  assign t[249] = t[276] ^ x[87];
  assign t[24] = t[43] ^ t[44];
  assign t[250] = t[277] ^ x[98];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = ~(t[45] ^ t[11]);
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[36];
  assign t[299] = t[353] ^ x[35];
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[39];
  assign t[301] = t[355] ^ x[38];
  assign t[302] = t[356] ^ x[42];
  assign t[303] = t[357] ^ x[41];
  assign t[304] = t[358] ^ x[45];
  assign t[305] = t[359] ^ x[44];
  assign t[306] = t[360] ^ x[48];
  assign t[307] = t[361] ^ x[47];
  assign t[308] = t[362] ^ x[51];
  assign t[309] = t[363] ^ x[50];
  assign t[30] = ~(t[199]);
  assign t[310] = t[364] ^ x[56];
  assign t[311] = t[365] ^ x[55];
  assign t[312] = t[366] ^ x[59];
  assign t[313] = t[367] ^ x[58];
  assign t[314] = t[368] ^ x[62];
  assign t[315] = t[369] ^ x[61];
  assign t[316] = t[370] ^ x[65];
  assign t[317] = t[371] ^ x[64];
  assign t[318] = t[372] ^ x[72];
  assign t[319] = t[373] ^ x[71];
  assign t[31] = ~(t[200]);
  assign t[320] = t[374] ^ x[75];
  assign t[321] = t[375] ^ x[74];
  assign t[322] = t[376] ^ x[78];
  assign t[323] = t[377] ^ x[77];
  assign t[324] = t[378] ^ x[81];
  assign t[325] = t[379] ^ x[80];
  assign t[326] = t[380] ^ x[84];
  assign t[327] = t[381] ^ x[83];
  assign t[328] = t[382] ^ x[87];
  assign t[329] = t[383] ^ x[86];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[384] ^ x[98];
  assign t[331] = t[385] ^ x[97];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = ~t[53];
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = ~t[54];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[34]);
  assign t[353] = (x[34]);
  assign t[354] = (x[37]);
  assign t[355] = (x[37]);
  assign t[356] = (x[40]);
  assign t[357] = (x[40]);
  assign t[358] = (x[43]);
  assign t[359] = (x[43]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[46]);
  assign t[361] = (x[46]);
  assign t[362] = (x[49]);
  assign t[363] = (x[49]);
  assign t[364] = (x[54]);
  assign t[365] = (x[54]);
  assign t[366] = (x[57]);
  assign t[367] = (x[57]);
  assign t[368] = (x[60]);
  assign t[369] = (x[60]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[63]);
  assign t[371] = (x[63]);
  assign t[372] = (x[70]);
  assign t[373] = (x[70]);
  assign t[374] = (x[73]);
  assign t[375] = (x[73]);
  assign t[376] = (x[76]);
  assign t[377] = (x[76]);
  assign t[378] = (x[79]);
  assign t[379] = (x[79]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[82]);
  assign t[381] = (x[82]);
  assign t[382] = (x[85]);
  assign t[383] = (x[85]);
  assign t[384] = (x[96]);
  assign t[385] = (x[96]);
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[27] ? t[66] : t[201];
  assign t[42] = t[67] ^ t[60];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = ~(t[72] ^ t[73]);
  assign t[46] = t[22] ^ t[74];
  assign t[47] = ~(t[75] ^ t[76]);
  assign t[48] = ~(t[77] & t[78]);
  assign t[49] = t[202] | t[79];
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[80]);
  assign t[51] = ~(t[203]);
  assign t[52] = ~(t[81] & t[204]);
  assign t[53] = t[8] ? t[82] : t[205];
  assign t[54] = t[8] ? t[83] : t[206];
  assign t[55] = t[84] & t[85];
  assign t[56] = t[86] & t[87];
  assign t[57] = ~(t[55] ^ t[88]);
  assign t[58] = t[89] ^ t[90];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] & t[94];
  assign t[61] = t[204] ^ t[95];
  assign t[62] = t[64] ^ t[96];
  assign t[63] = t[198] ^ t[97];
  assign t[64] = t[98] ^ t[99];
  assign t[65] = t[100] & t[101];
  assign t[66] = t[201] ^ t[102];
  assign t[67] = t[103] ^ t[104];
  assign t[68] = t[92] ^ t[41];
  assign t[69] = t[67] ^ t[105];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[106] ^ t[107];
  assign t[71] = t[108] & t[109];
  assign t[72] = t[110] ^ t[23];
  assign t[73] = t[111] ^ t[96];
  assign t[74] = t[112] ^ t[104];
  assign t[75] = t[34] ^ t[113];
  assign t[76] = t[114] ^ t[115];
  assign t[77] = ~(t[79] & t[116]);
  assign t[78] = ~(t[207] ^ t[117]);
  assign t[79] = ~(t[118] & t[119]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[49]);
  assign t[81] = ~(t[208]);
  assign t[82] = t[205] ^ t[120];
  assign t[83] = t[206] ^ t[121];
  assign t[84] = ~(t[90]);
  assign t[85] = ~(t[122]);
  assign t[86] = ~(t[33]);
  assign t[87] = t[123];
  assign t[88] = t[19] ^ t[122];
  assign t[89] = t[122] ^ t[34];
  assign t[8] = ~(t[15]);
  assign t[90] = t[87] ^ t[33];
  assign t[91] = t[27] ? t[124] : t[209];
  assign t[92] = t[27] ? t[125] : t[210];
  assign t[93] = ~(t[59] ^ t[67]);
  assign t[94] = t[68] ^ t[126];
  assign t[95] = t[127] ? t[128] : t[211];
  assign t[96] = t[129] & t[130];
  assign t[97] = t[127] ? t[131] : t[212];
  assign t[98] = t[132] & t[133];
  assign t[99] = t[134] & t[135];
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind101(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[98] ^ t[136]);
  assign t[101] = t[137] ^ t[138];
  assign t[102] = t[80] ? x[53] : x[52];
  assign t[103] = t[139] & t[140];
  assign t[104] = t[141] & t[126];
  assign t[105] = t[142] & t[143];
  assign t[106] = t[8] ? t[144] : t[213];
  assign t[107] = t[8] ? t[145] : t[214];
  assign t[108] = ~(t[70] ^ t[146]);
  assign t[109] = t[147] ^ t[148];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[147] ^ t[149];
  assign t[111] = t[150] ^ t[63];
  assign t[112] = t[91] ^ t[41];
  assign t[113] = t[35] ^ t[151];
  assign t[114] = t[8] ? t[152] : t[215];
  assign t[115] = t[146] ^ t[71];
  assign t[116] = ~(t[153] & t[154]);
  assign t[117] = t[155] ^ t[216];
  assign t[118] = ~(t[207]);
  assign t[119] = t[156] & t[155];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[28] ? x[67] : x[66];
  assign t[121] = t[28] ? x[69] : x[68];
  assign t[122] = t[157];
  assign t[123] = t[27] ? t[158] : t[217];
  assign t[124] = t[209] ^ t[159];
  assign t[125] = t[210] ^ t[160];
  assign t[126] = t[27] ? t[161] : t[218];
  assign t[127] = ~(t[15]);
  assign t[128] = t[211] ^ t[162];
  assign t[129] = ~(t[111] ^ t[64]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[39] ^ t[135];
  assign t[131] = t[212] ^ t[163];
  assign t[132] = ~(t[138]);
  assign t[133] = ~(t[150]);
  assign t[134] = ~(t[63]);
  assign t[135] = t[199] ^ t[164];
  assign t[136] = t[39] ^ t[150];
  assign t[137] = t[150] ^ t[61];
  assign t[138] = t[135] ^ t[63];
  assign t[139] = ~(t[165]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = ~(t[91]);
  assign t[141] = ~(t[92]);
  assign t[142] = ~(t[103] ^ t[166]);
  assign t[143] = t[112] ^ t[165];
  assign t[144] = t[213] ^ t[167];
  assign t[145] = t[214] ^ t[168];
  assign t[146] = t[169] ^ t[170];
  assign t[147] = t[107] ^ t[114];
  assign t[148] = t[8] ? t[171] : t[219];
  assign t[149] = t[146] ^ t[172];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[127] ? t[173] : t[220];
  assign t[151] = t[174] & t[175];
  assign t[152] = t[215] ^ t[176];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[177] | t[118]);
  assign t[155] = ~(t[221]);
  assign t[156] = ~(t[216]);
  assign t[157] = t[8] ? t[178] : t[222];
  assign t[158] = t[217] ^ t[179];
  assign t[159] = t[180] ? x[89] : x[88];
  assign t[15] = ~(t[27]);
  assign t[160] = t[180] ? x[91] : x[90];
  assign t[161] = t[218] ^ t[181];
  assign t[162] = t[182] ? x[93] : x[92];
  assign t[163] = t[182] ? x[95] : x[94];
  assign t[164] = t[127] ? t[183] : t[223];
  assign t[165] = t[126] ^ t[92];
  assign t[166] = t[68] ^ t[91];
  assign t[167] = t[28] ? x[100] : x[99];
  assign t[168] = t[28] ? x[102] : x[101];
  assign t[169] = t[184] & t[185];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[186] & t[148];
  assign t[171] = t[219] ^ t[187];
  assign t[172] = t[188] & t[189];
  assign t[173] = t[220] ^ t[190];
  assign t[174] = ~(t[191] ^ t[35]);
  assign t[175] = t[19] ^ t[87];
  assign t[176] = t[28] ? x[104] : x[103];
  assign t[177] = ~(t[202]);
  assign t[178] = t[222] ^ t[192];
  assign t[179] = t[28] ? x[106] : x[105];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[50]);
  assign t[181] = t[80] ? x[108] : x[107];
  assign t[182] = ~(t[50]);
  assign t[183] = t[223] ^ t[193];
  assign t[184] = ~(t[194]);
  assign t[185] = ~(t[106]);
  assign t[186] = ~(t[107]);
  assign t[187] = t[28] ? x[110] : x[109];
  assign t[188] = ~(t[169] ^ t[195]);
  assign t[189] = t[196] ^ t[194];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[182] ? x[112] : x[111];
  assign t[191] = t[122] ^ t[33];
  assign t[192] = t[28] ? x[114] : x[113];
  assign t[193] = t[182] ? x[116] : x[115];
  assign t[194] = t[148] ^ t[107];
  assign t[195] = t[147] ^ t[106];
  assign t[196] = t[106] ^ t[114];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = t[39] ^ t[40];
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[36];
  assign t[235] = t[262] ^ x[39];
  assign t[236] = t[263] ^ x[42];
  assign t[237] = t[264] ^ x[45];
  assign t[238] = t[265] ^ x[48];
  assign t[239] = t[266] ^ x[51];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[56];
  assign t[241] = t[268] ^ x[59];
  assign t[242] = t[269] ^ x[62];
  assign t[243] = t[270] ^ x[65];
  assign t[244] = t[271] ^ x[72];
  assign t[245] = t[272] ^ x[75];
  assign t[246] = t[273] ^ x[78];
  assign t[247] = t[274] ^ x[81];
  assign t[248] = t[275] ^ x[84];
  assign t[249] = t[276] ^ x[87];
  assign t[24] = t[43] ^ t[44];
  assign t[250] = t[277] ^ x[98];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = ~(t[45] ^ t[11]);
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[36];
  assign t[299] = t[353] ^ x[35];
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[39];
  assign t[301] = t[355] ^ x[38];
  assign t[302] = t[356] ^ x[42];
  assign t[303] = t[357] ^ x[41];
  assign t[304] = t[358] ^ x[45];
  assign t[305] = t[359] ^ x[44];
  assign t[306] = t[360] ^ x[48];
  assign t[307] = t[361] ^ x[47];
  assign t[308] = t[362] ^ x[51];
  assign t[309] = t[363] ^ x[50];
  assign t[30] = ~(t[199]);
  assign t[310] = t[364] ^ x[56];
  assign t[311] = t[365] ^ x[55];
  assign t[312] = t[366] ^ x[59];
  assign t[313] = t[367] ^ x[58];
  assign t[314] = t[368] ^ x[62];
  assign t[315] = t[369] ^ x[61];
  assign t[316] = t[370] ^ x[65];
  assign t[317] = t[371] ^ x[64];
  assign t[318] = t[372] ^ x[72];
  assign t[319] = t[373] ^ x[71];
  assign t[31] = ~(t[200]);
  assign t[320] = t[374] ^ x[75];
  assign t[321] = t[375] ^ x[74];
  assign t[322] = t[376] ^ x[78];
  assign t[323] = t[377] ^ x[77];
  assign t[324] = t[378] ^ x[81];
  assign t[325] = t[379] ^ x[80];
  assign t[326] = t[380] ^ x[84];
  assign t[327] = t[381] ^ x[83];
  assign t[328] = t[382] ^ x[87];
  assign t[329] = t[383] ^ x[86];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[384] ^ x[98];
  assign t[331] = t[385] ^ x[97];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = ~t[53];
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = ~t[54];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[34]);
  assign t[353] = (x[34]);
  assign t[354] = (x[37]);
  assign t[355] = (x[37]);
  assign t[356] = (x[40]);
  assign t[357] = (x[40]);
  assign t[358] = (x[43]);
  assign t[359] = (x[43]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[46]);
  assign t[361] = (x[46]);
  assign t[362] = (x[49]);
  assign t[363] = (x[49]);
  assign t[364] = (x[54]);
  assign t[365] = (x[54]);
  assign t[366] = (x[57]);
  assign t[367] = (x[57]);
  assign t[368] = (x[60]);
  assign t[369] = (x[60]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[63]);
  assign t[371] = (x[63]);
  assign t[372] = (x[70]);
  assign t[373] = (x[70]);
  assign t[374] = (x[73]);
  assign t[375] = (x[73]);
  assign t[376] = (x[76]);
  assign t[377] = (x[76]);
  assign t[378] = (x[79]);
  assign t[379] = (x[79]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[82]);
  assign t[381] = (x[82]);
  assign t[382] = (x[85]);
  assign t[383] = (x[85]);
  assign t[384] = (x[96]);
  assign t[385] = (x[96]);
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[27] ? t[66] : t[201];
  assign t[42] = t[67] ^ t[60];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = ~(t[72] ^ t[73]);
  assign t[46] = t[22] ^ t[74];
  assign t[47] = ~(t[75] ^ t[76]);
  assign t[48] = ~(t[77] & t[78]);
  assign t[49] = t[202] | t[79];
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[80]);
  assign t[51] = ~(t[203]);
  assign t[52] = ~(t[81] & t[204]);
  assign t[53] = t[8] ? t[82] : t[205];
  assign t[54] = t[8] ? t[83] : t[206];
  assign t[55] = t[84] & t[85];
  assign t[56] = t[86] & t[87];
  assign t[57] = ~(t[55] ^ t[88]);
  assign t[58] = t[89] ^ t[90];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] & t[94];
  assign t[61] = t[204] ^ t[95];
  assign t[62] = t[64] ^ t[96];
  assign t[63] = t[198] ^ t[97];
  assign t[64] = t[98] ^ t[99];
  assign t[65] = t[100] & t[101];
  assign t[66] = t[201] ^ t[102];
  assign t[67] = t[103] ^ t[104];
  assign t[68] = t[92] ^ t[41];
  assign t[69] = t[67] ^ t[105];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[106] ^ t[107];
  assign t[71] = t[108] & t[109];
  assign t[72] = t[110] ^ t[23];
  assign t[73] = t[111] ^ t[96];
  assign t[74] = t[112] ^ t[104];
  assign t[75] = t[34] ^ t[113];
  assign t[76] = t[114] ^ t[115];
  assign t[77] = ~(t[79] & t[116]);
  assign t[78] = ~(t[207] ^ t[117]);
  assign t[79] = ~(t[118] & t[119]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[49]);
  assign t[81] = ~(t[208]);
  assign t[82] = t[205] ^ t[120];
  assign t[83] = t[206] ^ t[121];
  assign t[84] = ~(t[90]);
  assign t[85] = ~(t[122]);
  assign t[86] = ~(t[33]);
  assign t[87] = t[123];
  assign t[88] = t[19] ^ t[122];
  assign t[89] = t[122] ^ t[34];
  assign t[8] = ~(t[15]);
  assign t[90] = t[87] ^ t[33];
  assign t[91] = t[27] ? t[124] : t[209];
  assign t[92] = t[27] ? t[125] : t[210];
  assign t[93] = ~(t[59] ^ t[67]);
  assign t[94] = t[68] ^ t[126];
  assign t[95] = t[127] ? t[128] : t[211];
  assign t[96] = t[129] & t[130];
  assign t[97] = t[127] ? t[131] : t[212];
  assign t[98] = t[132] & t[133];
  assign t[99] = t[134] & t[135];
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[88]);
  assign t[101] = t[138];
  assign t[102] = t[88] ^ t[23];
  assign t[103] = t[136] ? x[61] : x[60];
  assign t[104] = t[136] ? x[63] : x[62];
  assign t[105] = t[139] & t[140];
  assign t[106] = t[141] & t[72];
  assign t[107] = t[8] ? t[142] : t[215];
  assign t[108] = t[207] ^ t[143];
  assign t[109] = ~(t[144] & t[145]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[146] ^ t[216];
  assign t[111] = ~(t[208]);
  assign t[112] = t[147] & t[146];
  assign t[113] = t[148] ^ t[65];
  assign t[114] = ~(t[149] ^ t[39]);
  assign t[115] = t[150] ^ t[151];
  assign t[116] = t[43] ^ t[107];
  assign t[117] = t[70] ^ t[26];
  assign t[118] = t[210] ^ t[152];
  assign t[119] = t[211] ^ t[153];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[27] ? t[154] : t[217];
  assign t[121] = t[212] ^ t[155];
  assign t[122] = t[156] & t[157];
  assign t[123] = t[158] ^ t[54];
  assign t[124] = t[159] & t[160];
  assign t[125] = t[8] ? t[161] : t[218];
  assign t[126] = t[8] ? t[162] : t[219];
  assign t[127] = ~(t[15]);
  assign t[128] = t[213] ^ t[163];
  assign t[129] = t[198] ^ t[164];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[127] ? t[165] : t[220];
  assign t[131] = t[166] & t[167];
  assign t[132] = t[214] ^ t[168];
  assign t[133] = t[169] & t[170];
  assign t[134] = ~(t[171] ^ t[95]);
  assign t[135] = t[150] ^ t[91];
  assign t[136] = ~(t[172]);
  assign t[137] = t[101] ^ t[88];
  assign t[138] = t[27] ? t[173] : t[221];
  assign t[139] = ~(t[174]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[43]);
  assign t[141] = ~(t[44]);
  assign t[142] = t[215] ^ t[175];
  assign t[143] = t[136] ? x[86] : x[85];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[176] | t[111]);
  assign t[146] = ~(t[222]);
  assign t[147] = ~(t[216]);
  assign t[148] = t[87] ^ t[23];
  assign t[149] = t[177] ^ t[124];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[129] ^ t[61];
  assign t[151] = t[95] ^ t[178];
  assign t[152] = t[179] ? x[91] : x[90];
  assign t[153] = t[28] ? x[93] : x[92];
  assign t[154] = t[217] ^ t[180];
  assign t[155] = t[28] ? x[95] : x[94];
  assign t[156] = ~(t[105] ^ t[181]);
  assign t[157] = t[116] ^ t[174];
  assign t[158] = t[182] & t[183];
  assign t[159] = ~(t[177] ^ t[123]);
  assign t[15] = ~(t[27]);
  assign t[160] = t[92] ^ t[84];
  assign t[161] = t[218] ^ t[184];
  assign t[162] = t[219] ^ t[185];
  assign t[163] = t[186] ? x[97] : x[96];
  assign t[164] = t[127] ? t[187] : t[223];
  assign t[165] = t[220] ^ t[188];
  assign t[166] = ~(t[158] ^ t[189]);
  assign t[167] = t[53] ^ t[190];
  assign t[168] = t[186] ? x[102] : x[101];
  assign t[169] = ~(t[191]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[89]);
  assign t[171] = t[89] ^ t[129];
  assign t[172] = ~(t[28]);
  assign t[173] = t[221] ^ t[192];
  assign t[174] = t[72] ^ t[44];
  assign t[175] = t[136] ? x[104] : x[103];
  assign t[176] = ~(t[204]);
  assign t[177] = t[81] ^ t[120];
  assign t[178] = t[193] & t[194];
  assign t[179] = ~(t[172]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[179] ? x[106] : x[105];
  assign t[181] = t[71] ^ t[43];
  assign t[182] = ~(t[190]);
  assign t[183] = ~(t[81]);
  assign t[184] = t[136] ? x[108] : x[107];
  assign t[185] = t[136] ? x[110] : x[109];
  assign t[186] = ~(t[172]);
  assign t[187] = t[223] ^ t[195];
  assign t[188] = t[186] ? x[112] : x[111];
  assign t[189] = t[92] ^ t[81];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[84] ^ t[120];
  assign t[191] = t[91] ^ t[129];
  assign t[192] = t[136] ? x[114] : x[113];
  assign t[193] = ~(t[133] ^ t[196]);
  assign t[194] = t[58] ^ t[191];
  assign t[195] = t[186] ? x[116] : x[115];
  assign t[196] = t[150] ^ t[89];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[36];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = ~(t[38] ^ t[39]);
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[36];
  assign t[235] = t[262] ^ x[39];
  assign t[236] = t[263] ^ x[42];
  assign t[237] = t[264] ^ x[45];
  assign t[238] = t[265] ^ x[48];
  assign t[239] = t[266] ^ x[51];
  assign t[23] = ~t[40];
  assign t[240] = t[267] ^ x[54];
  assign t[241] = t[268] ^ x[57];
  assign t[242] = t[269] ^ x[66];
  assign t[243] = t[270] ^ x[69];
  assign t[244] = t[271] ^ x[72];
  assign t[245] = t[272] ^ x[75];
  assign t[246] = t[273] ^ x[78];
  assign t[247] = t[274] ^ x[81];
  assign t[248] = t[275] ^ x[84];
  assign t[249] = t[276] ^ x[89];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[277] ^ x[100];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = t[43] ^ t[44];
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = t[45] & t[46];
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[48]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[36];
  assign t[299] = t[353] ^ x[35];
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[39];
  assign t[301] = t[355] ^ x[38];
  assign t[302] = t[356] ^ x[42];
  assign t[303] = t[357] ^ x[41];
  assign t[304] = t[358] ^ x[45];
  assign t[305] = t[359] ^ x[44];
  assign t[306] = t[360] ^ x[48];
  assign t[307] = t[361] ^ x[47];
  assign t[308] = t[362] ^ x[51];
  assign t[309] = t[363] ^ x[50];
  assign t[30] = ~(t[199]);
  assign t[310] = t[364] ^ x[54];
  assign t[311] = t[365] ^ x[53];
  assign t[312] = t[366] ^ x[57];
  assign t[313] = t[367] ^ x[56];
  assign t[314] = t[368] ^ x[66];
  assign t[315] = t[369] ^ x[65];
  assign t[316] = t[370] ^ x[69];
  assign t[317] = t[371] ^ x[68];
  assign t[318] = t[372] ^ x[72];
  assign t[319] = t[373] ^ x[71];
  assign t[31] = ~(t[200]);
  assign t[320] = t[374] ^ x[75];
  assign t[321] = t[375] ^ x[74];
  assign t[322] = t[376] ^ x[78];
  assign t[323] = t[377] ^ x[77];
  assign t[324] = t[378] ^ x[81];
  assign t[325] = t[379] ^ x[80];
  assign t[326] = t[380] ^ x[84];
  assign t[327] = t[381] ^ x[83];
  assign t[328] = t[382] ^ x[89];
  assign t[329] = t[383] ^ x[88];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[100];
  assign t[331] = t[385] ^ x[99];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = ~(t[51] ^ t[52]);
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = t[53] ^ t[54];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[34]);
  assign t[353] = (x[34]);
  assign t[354] = (x[37]);
  assign t[355] = (x[37]);
  assign t[356] = (x[40]);
  assign t[357] = (x[40]);
  assign t[358] = (x[43]);
  assign t[359] = (x[43]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[46]);
  assign t[361] = (x[46]);
  assign t[362] = (x[49]);
  assign t[363] = (x[49]);
  assign t[364] = (x[52]);
  assign t[365] = (x[52]);
  assign t[366] = (x[55]);
  assign t[367] = (x[55]);
  assign t[368] = (x[64]);
  assign t[369] = (x[64]);
  assign t[36] = t[57] ^ t[42];
  assign t[370] = (x[67]);
  assign t[371] = (x[67]);
  assign t[372] = (x[70]);
  assign t[373] = (x[70]);
  assign t[374] = (x[73]);
  assign t[375] = (x[73]);
  assign t[376] = (x[76]);
  assign t[377] = (x[76]);
  assign t[378] = (x[79]);
  assign t[379] = (x[79]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[82]);
  assign t[381] = (x[82]);
  assign t[382] = (x[87]);
  assign t[383] = (x[87]);
  assign t[384] = (x[98]);
  assign t[385] = (x[98]);
  assign t[38] = t[60] ^ t[14];
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[63] : t[201];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] & t[67];
  assign t[43] = t[8] ? t[68] : t[202];
  assign t[44] = t[8] ? t[69] : t[203];
  assign t[45] = ~(t[25] ^ t[70]);
  assign t[46] = t[71] ^ t[72];
  assign t[47] = ~(t[73] & t[74]);
  assign t[48] = t[204] | t[75];
  assign t[49] = ~(t[205]);
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[76] & t[206]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[71] ^ t[85];
  assign t[56] = t[82] ^ t[86];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] ^ t[61];
  assign t[59] = t[90] & t[91];
  assign t[5] = ~(t[10]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[206] ^ t[94];
  assign t[62] = t[95] ^ t[96];
  assign t[63] = t[201] ^ t[97];
  assign t[64] = t[98] & t[99];
  assign t[65] = t[100] & t[101];
  assign t[66] = ~(t[57] ^ t[41]);
  assign t[67] = t[102] ^ t[101];
  assign t[68] = t[202] ^ t[103];
  assign t[69] = t[203] ^ t[104];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[105] ^ t[106];
  assign t[71] = t[44] ^ t[107];
  assign t[72] = t[8] ? t[108] : t[207];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[208] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[209]);
  assign t[77] = t[13] ^ t[113];
  assign t[78] = ~(t[114] ^ t[115]);
  assign t[79] = t[116] ^ t[106];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[107] ^ t[117];
  assign t[81] = t[27] ? t[118] : t[210];
  assign t[82] = t[27] ? t[119] : t[211];
  assign t[83] = ~(t[120]);
  assign t[84] = t[27] ? t[121] : t[212];
  assign t[85] = t[70] ^ t[122];
  assign t[86] = t[123] ^ t[124];
  assign t[87] = t[125];
  assign t[88] = ~t[126];
  assign t[89] = t[127] ? t[128] : t[213];
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[129]);
  assign t[91] = t[199] ^ t[130];
  assign t[92] = t[120] ^ t[82];
  assign t[93] = t[123] ^ t[131];
  assign t[94] = t[127] ? t[132] : t[214];
  assign t[95] = t[133] ^ t[59];
  assign t[96] = t[134] & t[135];
  assign t[97] = t[136] ? x[59] : x[58];
  assign t[98] = ~(t[137]);
  assign t[99] = ~(t[87]);
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[88]);
  assign t[101] = t[138];
  assign t[102] = t[88] ^ t[23];
  assign t[103] = t[136] ? x[61] : x[60];
  assign t[104] = t[136] ? x[63] : x[62];
  assign t[105] = t[139] & t[140];
  assign t[106] = t[141] & t[72];
  assign t[107] = t[8] ? t[142] : t[215];
  assign t[108] = t[207] ^ t[143];
  assign t[109] = ~(t[144] & t[145]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[146] ^ t[216];
  assign t[111] = ~(t[208]);
  assign t[112] = t[147] & t[146];
  assign t[113] = t[148] ^ t[65];
  assign t[114] = ~(t[149] ^ t[39]);
  assign t[115] = t[150] ^ t[151];
  assign t[116] = t[43] ^ t[107];
  assign t[117] = t[70] ^ t[26];
  assign t[118] = t[210] ^ t[152];
  assign t[119] = t[211] ^ t[153];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[27] ? t[154] : t[217];
  assign t[121] = t[212] ^ t[155];
  assign t[122] = t[156] & t[157];
  assign t[123] = t[158] ^ t[54];
  assign t[124] = t[159] & t[160];
  assign t[125] = t[8] ? t[161] : t[218];
  assign t[126] = t[8] ? t[162] : t[219];
  assign t[127] = ~(t[15]);
  assign t[128] = t[213] ^ t[163];
  assign t[129] = t[198] ^ t[164];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[127] ? t[165] : t[220];
  assign t[131] = t[166] & t[167];
  assign t[132] = t[214] ^ t[168];
  assign t[133] = t[169] & t[170];
  assign t[134] = ~(t[171] ^ t[95]);
  assign t[135] = t[150] ^ t[91];
  assign t[136] = ~(t[172]);
  assign t[137] = t[101] ^ t[88];
  assign t[138] = t[27] ? t[173] : t[221];
  assign t[139] = ~(t[174]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = ~(t[43]);
  assign t[141] = ~(t[44]);
  assign t[142] = t[215] ^ t[175];
  assign t[143] = t[136] ? x[86] : x[85];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[176] | t[111]);
  assign t[146] = ~(t[222]);
  assign t[147] = ~(t[216]);
  assign t[148] = t[87] ^ t[23];
  assign t[149] = t[177] ^ t[124];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[129] ^ t[61];
  assign t[151] = t[95] ^ t[178];
  assign t[152] = t[179] ? x[91] : x[90];
  assign t[153] = t[28] ? x[93] : x[92];
  assign t[154] = t[217] ^ t[180];
  assign t[155] = t[28] ? x[95] : x[94];
  assign t[156] = ~(t[105] ^ t[181]);
  assign t[157] = t[116] ^ t[174];
  assign t[158] = t[182] & t[183];
  assign t[159] = ~(t[177] ^ t[123]);
  assign t[15] = ~(t[27]);
  assign t[160] = t[92] ^ t[84];
  assign t[161] = t[218] ^ t[184];
  assign t[162] = t[219] ^ t[185];
  assign t[163] = t[186] ? x[97] : x[96];
  assign t[164] = t[127] ? t[187] : t[223];
  assign t[165] = t[220] ^ t[188];
  assign t[166] = ~(t[158] ^ t[189]);
  assign t[167] = t[53] ^ t[190];
  assign t[168] = t[186] ? x[102] : x[101];
  assign t[169] = ~(t[191]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[89]);
  assign t[171] = t[89] ^ t[129];
  assign t[172] = ~(t[28]);
  assign t[173] = t[221] ^ t[192];
  assign t[174] = t[72] ^ t[44];
  assign t[175] = t[136] ? x[104] : x[103];
  assign t[176] = ~(t[204]);
  assign t[177] = t[81] ^ t[120];
  assign t[178] = t[193] & t[194];
  assign t[179] = ~(t[172]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[179] ? x[106] : x[105];
  assign t[181] = t[71] ^ t[43];
  assign t[182] = ~(t[190]);
  assign t[183] = ~(t[81]);
  assign t[184] = t[136] ? x[108] : x[107];
  assign t[185] = t[136] ? x[110] : x[109];
  assign t[186] = ~(t[172]);
  assign t[187] = t[223] ^ t[195];
  assign t[188] = t[186] ? x[112] : x[111];
  assign t[189] = t[92] ^ t[81];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[84] ^ t[120];
  assign t[191] = t[91] ^ t[129];
  assign t[192] = t[136] ? x[114] : x[113];
  assign t[193] = ~(t[133] ^ t[196]);
  assign t[194] = t[58] ^ t[191];
  assign t[195] = t[186] ? x[116] : x[115];
  assign t[196] = t[150] ^ t[89];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[36];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = ~(t[38] ^ t[39]);
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[36];
  assign t[235] = t[262] ^ x[39];
  assign t[236] = t[263] ^ x[42];
  assign t[237] = t[264] ^ x[45];
  assign t[238] = t[265] ^ x[48];
  assign t[239] = t[266] ^ x[51];
  assign t[23] = ~t[40];
  assign t[240] = t[267] ^ x[54];
  assign t[241] = t[268] ^ x[57];
  assign t[242] = t[269] ^ x[66];
  assign t[243] = t[270] ^ x[69];
  assign t[244] = t[271] ^ x[72];
  assign t[245] = t[272] ^ x[75];
  assign t[246] = t[273] ^ x[78];
  assign t[247] = t[274] ^ x[81];
  assign t[248] = t[275] ^ x[84];
  assign t[249] = t[276] ^ x[89];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[277] ^ x[100];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = t[43] ^ t[44];
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = t[45] & t[46];
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[48]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[36];
  assign t[299] = t[353] ^ x[35];
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[39];
  assign t[301] = t[355] ^ x[38];
  assign t[302] = t[356] ^ x[42];
  assign t[303] = t[357] ^ x[41];
  assign t[304] = t[358] ^ x[45];
  assign t[305] = t[359] ^ x[44];
  assign t[306] = t[360] ^ x[48];
  assign t[307] = t[361] ^ x[47];
  assign t[308] = t[362] ^ x[51];
  assign t[309] = t[363] ^ x[50];
  assign t[30] = ~(t[199]);
  assign t[310] = t[364] ^ x[54];
  assign t[311] = t[365] ^ x[53];
  assign t[312] = t[366] ^ x[57];
  assign t[313] = t[367] ^ x[56];
  assign t[314] = t[368] ^ x[66];
  assign t[315] = t[369] ^ x[65];
  assign t[316] = t[370] ^ x[69];
  assign t[317] = t[371] ^ x[68];
  assign t[318] = t[372] ^ x[72];
  assign t[319] = t[373] ^ x[71];
  assign t[31] = ~(t[200]);
  assign t[320] = t[374] ^ x[75];
  assign t[321] = t[375] ^ x[74];
  assign t[322] = t[376] ^ x[78];
  assign t[323] = t[377] ^ x[77];
  assign t[324] = t[378] ^ x[81];
  assign t[325] = t[379] ^ x[80];
  assign t[326] = t[380] ^ x[84];
  assign t[327] = t[381] ^ x[83];
  assign t[328] = t[382] ^ x[89];
  assign t[329] = t[383] ^ x[88];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[100];
  assign t[331] = t[385] ^ x[99];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = ~(t[51] ^ t[52]);
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = t[53] ^ t[54];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[34]);
  assign t[353] = (x[34]);
  assign t[354] = (x[37]);
  assign t[355] = (x[37]);
  assign t[356] = (x[40]);
  assign t[357] = (x[40]);
  assign t[358] = (x[43]);
  assign t[359] = (x[43]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[46]);
  assign t[361] = (x[46]);
  assign t[362] = (x[49]);
  assign t[363] = (x[49]);
  assign t[364] = (x[52]);
  assign t[365] = (x[52]);
  assign t[366] = (x[55]);
  assign t[367] = (x[55]);
  assign t[368] = (x[64]);
  assign t[369] = (x[64]);
  assign t[36] = t[57] ^ t[42];
  assign t[370] = (x[67]);
  assign t[371] = (x[67]);
  assign t[372] = (x[70]);
  assign t[373] = (x[70]);
  assign t[374] = (x[73]);
  assign t[375] = (x[73]);
  assign t[376] = (x[76]);
  assign t[377] = (x[76]);
  assign t[378] = (x[79]);
  assign t[379] = (x[79]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[82]);
  assign t[381] = (x[82]);
  assign t[382] = (x[87]);
  assign t[383] = (x[87]);
  assign t[384] = (x[98]);
  assign t[385] = (x[98]);
  assign t[38] = t[60] ^ t[14];
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[8] ? t[63] : t[201];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] & t[67];
  assign t[43] = t[8] ? t[68] : t[202];
  assign t[44] = t[8] ? t[69] : t[203];
  assign t[45] = ~(t[25] ^ t[70]);
  assign t[46] = t[71] ^ t[72];
  assign t[47] = ~(t[73] & t[74]);
  assign t[48] = t[204] | t[75];
  assign t[49] = ~(t[205]);
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[76] & t[206]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[71] ^ t[85];
  assign t[56] = t[82] ^ t[86];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] ^ t[61];
  assign t[59] = t[90] & t[91];
  assign t[5] = ~(t[10]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[206] ^ t[94];
  assign t[62] = t[95] ^ t[96];
  assign t[63] = t[201] ^ t[97];
  assign t[64] = t[98] & t[99];
  assign t[65] = t[100] & t[101];
  assign t[66] = ~(t[57] ^ t[41]);
  assign t[67] = t[102] ^ t[101];
  assign t[68] = t[202] ^ t[103];
  assign t[69] = t[203] ^ t[104];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[105] ^ t[106];
  assign t[71] = t[44] ^ t[107];
  assign t[72] = t[8] ? t[108] : t[207];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[208] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[209]);
  assign t[77] = t[13] ^ t[113];
  assign t[78] = ~(t[114] ^ t[115]);
  assign t[79] = t[116] ^ t[106];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[107] ^ t[117];
  assign t[81] = t[27] ? t[118] : t[210];
  assign t[82] = t[27] ? t[119] : t[211];
  assign t[83] = ~(t[120]);
  assign t[84] = t[27] ? t[121] : t[212];
  assign t[85] = t[70] ^ t[122];
  assign t[86] = t[123] ^ t[124];
  assign t[87] = t[125];
  assign t[88] = ~t[126];
  assign t[89] = t[127] ? t[128] : t[213];
  assign t[8] = ~(t[15]);
  assign t[90] = ~(t[129]);
  assign t[91] = t[199] ^ t[130];
  assign t[92] = t[120] ^ t[82];
  assign t[93] = t[123] ^ t[131];
  assign t[94] = t[127] ? t[132] : t[214];
  assign t[95] = t[133] ^ t[59];
  assign t[96] = t[134] & t[135];
  assign t[97] = t[136] ? x[59] : x[58];
  assign t[98] = ~(t[137]);
  assign t[99] = ~(t[87]);
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [116:0] x;
 output y;

 wire [378:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[8] ? t[136] : t[207];
  assign t[101] = t[127] ^ t[60];
  assign t[102] = t[137] ? t[138] : t[208];
  assign t[103] = t[137] ? t[139] : t[209];
  assign t[104] = ~(t[69] ^ t[140]);
  assign t[105] = t[141] ^ t[142];
  assign t[106] = t[143] & t[144];
  assign t[107] = ~(t[106] ^ t[145]);
  assign t[108] = t[19] ^ t[146];
  assign t[109] = ~(t[147] & t[148]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[149] ^ t[210];
  assign t[111] = ~(t[203]);
  assign t[112] = t[150] & t[149];
  assign t[113] = ~(t[50]);
  assign t[114] = t[113] ? x[70] : x[69];
  assign t[115] = t[204] ^ t[151];
  assign t[116] = t[113] ? x[72] : x[71];
  assign t[117] = t[102] ^ t[123];
  assign t[118] = t[152] & t[142];
  assign t[119] = t[33] ^ t[55];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[153] & t[154];
  assign t[121] = t[128] ^ t[155];
  assign t[122] = t[156] ^ t[90];
  assign t[123] = t[137] ? t[157] : t[211];
  assign t[124] = t[140] ^ t[70];
  assign t[125] = t[205] ^ t[158];
  assign t[126] = t[206] ^ t[159];
  assign t[127] = t[160] ^ t[161];
  assign t[128] = t[87] ^ t[100];
  assign t[129] = t[8] ? t[162] : t[212];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = ~(t[156] ^ t[42]);
  assign t[131] = t[23] ^ t[96];
  assign t[132] = t[113] ? x[80] : x[79];
  assign t[133] = t[76] ? x[82] : x[81];
  assign t[134] = t[163];
  assign t[135] = t[8] ? t[164] : t[213];
  assign t[136] = t[207] ^ t[165];
  assign t[137] = ~(t[15]);
  assign t[138] = t[208] ^ t[166];
  assign t[139] = t[209] ^ t[167];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[168] ^ t[118];
  assign t[141] = t[103] ^ t[123];
  assign t[142] = t[137] ? t[169] : t[214];
  assign t[143] = ~(t[146]);
  assign t[144] = ~(t[33]);
  assign t[145] = t[46] ^ t[33];
  assign t[146] = t[36] ^ t[55];
  assign t[147] = ~(t[150] | t[149]);
  assign t[148] = ~(t[170] | t[111]);
  assign t[149] = ~(t[215]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[210]);
  assign t[151] = t[113] ? x[93] : x[92];
  assign t[152] = ~(t[103]);
  assign t[153] = ~(t[119] ^ t[71]);
  assign t[154] = t[46] ^ t[36];
  assign t[155] = t[127] ^ t[171];
  assign t[156] = t[134] ^ t[40];
  assign t[157] = t[211] ^ t[172];
  assign t[158] = t[28] ? x[95] : x[94];
  assign t[159] = t[28] ? x[97] : x[96];
  assign t[15] = ~(t[27]);
  assign t[160] = t[173] & t[174];
  assign t[161] = t[175] & t[129];
  assign t[162] = t[212] ^ t[176];
  assign t[163] = t[8] ? t[177] : t[216];
  assign t[164] = t[213] ^ t[178];
  assign t[165] = t[76] ? x[102] : x[101];
  assign t[166] = t[179] ? x[104] : x[103];
  assign t[167] = t[179] ? x[106] : x[105];
  assign t[168] = t[180] & t[181];
  assign t[169] = t[214] ^ t[182];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[197]);
  assign t[171] = t[183] & t[184];
  assign t[172] = t[179] ? x[108] : x[107];
  assign t[173] = ~(t[185]);
  assign t[174] = ~(t[86]);
  assign t[175] = ~(t[87]);
  assign t[176] = t[28] ? x[110] : x[109];
  assign t[177] = t[216] ^ t[186];
  assign t[178] = t[76] ? x[112] : x[111];
  assign t[179] = ~(t[50]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[187]);
  assign t[181] = ~(t[102]);
  assign t[182] = t[179] ? x[114] : x[113];
  assign t[183] = ~(t[160] ^ t[188]);
  assign t[184] = t[189] ^ t[185];
  assign t[185] = t[129] ^ t[87];
  assign t[186] = t[76] ? x[116] : x[115];
  assign t[187] = t[142] ^ t[103];
  assign t[188] = t[128] ^ t[86];
  assign t[189] = t[86] ^ t[100];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] & t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = t[244] ^ x[4];
  assign t[218] = t[245] ^ x[9];
  assign t[219] = t[246] ^ x[12];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[15];
  assign t[221] = t[248] ^ x[18];
  assign t[222] = t[249] ^ x[21];
  assign t[223] = t[250] ^ x[24];
  assign t[224] = t[251] ^ x[27];
  assign t[225] = t[252] ^ x[30];
  assign t[226] = t[253] ^ x[33];
  assign t[227] = t[254] ^ x[36];
  assign t[228] = t[255] ^ x[39];
  assign t[229] = t[256] ^ x[42];
  assign t[22] = ~(t[26] ^ t[39]);
  assign t[230] = t[257] ^ x[45];
  assign t[231] = t[258] ^ x[50];
  assign t[232] = t[259] ^ x[53];
  assign t[233] = t[260] ^ x[56];
  assign t[234] = t[261] ^ x[59];
  assign t[235] = t[262] ^ x[62];
  assign t[236] = t[263] ^ x[65];
  assign t[237] = t[264] ^ x[68];
  assign t[238] = t[265] ^ x[75];
  assign t[239] = t[266] ^ x[78];
  assign t[23] = t[40] ^ t[41];
  assign t[240] = t[267] ^ x[85];
  assign t[241] = t[268] ^ x[88];
  assign t[242] = t[269] ^ x[91];
  assign t[243] = t[270] ^ x[100];
  assign t[244] = (t[271] & ~t[272]);
  assign t[245] = (t[273] & ~t[274]);
  assign t[246] = (t[275] & ~t[276]);
  assign t[247] = (t[277] & ~t[278]);
  assign t[248] = (t[279] & ~t[280]);
  assign t[249] = (t[281] & ~t[282]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[283] & ~t[284]);
  assign t[251] = (t[285] & ~t[286]);
  assign t[252] = (t[287] & ~t[288]);
  assign t[253] = (t[289] & ~t[290]);
  assign t[254] = (t[291] & ~t[292]);
  assign t[255] = (t[293] & ~t[294]);
  assign t[256] = (t[295] & ~t[296]);
  assign t[257] = (t[297] & ~t[298]);
  assign t[258] = (t[299] & ~t[300]);
  assign t[259] = (t[301] & ~t[302]);
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[260] = (t[303] & ~t[304]);
  assign t[261] = (t[305] & ~t[306]);
  assign t[262] = (t[307] & ~t[308]);
  assign t[263] = (t[309] & ~t[310]);
  assign t[264] = (t[311] & ~t[312]);
  assign t[265] = (t[313] & ~t[314]);
  assign t[266] = (t[315] & ~t[316]);
  assign t[267] = (t[317] & ~t[318]);
  assign t[268] = (t[319] & ~t[320]);
  assign t[269] = (t[321] & ~t[322]);
  assign t[26] = t[46] ^ t[47];
  assign t[270] = (t[323] & ~t[324]);
  assign t[271] = t[325] ^ x[4];
  assign t[272] = t[326] ^ x[3];
  assign t[273] = t[327] ^ x[9];
  assign t[274] = t[328] ^ x[8];
  assign t[275] = t[329] ^ x[12];
  assign t[276] = t[330] ^ x[11];
  assign t[277] = t[331] ^ x[15];
  assign t[278] = t[332] ^ x[14];
  assign t[279] = t[333] ^ x[18];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[17];
  assign t[281] = t[335] ^ x[21];
  assign t[282] = t[336] ^ x[20];
  assign t[283] = t[337] ^ x[24];
  assign t[284] = t[338] ^ x[23];
  assign t[285] = t[339] ^ x[27];
  assign t[286] = t[340] ^ x[26];
  assign t[287] = t[341] ^ x[30];
  assign t[288] = t[342] ^ x[29];
  assign t[289] = t[343] ^ x[33];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[32];
  assign t[291] = t[345] ^ x[36];
  assign t[292] = t[346] ^ x[35];
  assign t[293] = t[347] ^ x[39];
  assign t[294] = t[348] ^ x[38];
  assign t[295] = t[349] ^ x[42];
  assign t[296] = t[350] ^ x[41];
  assign t[297] = t[351] ^ x[45];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[50];
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[49];
  assign t[301] = t[355] ^ x[53];
  assign t[302] = t[356] ^ x[52];
  assign t[303] = t[357] ^ x[56];
  assign t[304] = t[358] ^ x[55];
  assign t[305] = t[359] ^ x[59];
  assign t[306] = t[360] ^ x[58];
  assign t[307] = t[361] ^ x[62];
  assign t[308] = t[362] ^ x[61];
  assign t[309] = t[363] ^ x[65];
  assign t[30] = ~(t[192]);
  assign t[310] = t[364] ^ x[64];
  assign t[311] = t[365] ^ x[68];
  assign t[312] = t[366] ^ x[67];
  assign t[313] = t[367] ^ x[75];
  assign t[314] = t[368] ^ x[74];
  assign t[315] = t[369] ^ x[78];
  assign t[316] = t[370] ^ x[77];
  assign t[317] = t[371] ^ x[85];
  assign t[318] = t[372] ^ x[84];
  assign t[319] = t[373] ^ x[88];
  assign t[31] = ~(t[193]);
  assign t[320] = t[374] ^ x[87];
  assign t[321] = t[375] ^ x[91];
  assign t[322] = t[376] ^ x[90];
  assign t[323] = t[377] ^ x[100];
  assign t[324] = t[378] ^ x[99];
  assign t[325] = (x[2]);
  assign t[326] = (x[2]);
  assign t[327] = (x[7]);
  assign t[328] = (x[7]);
  assign t[329] = (x[10]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[10]);
  assign t[331] = (x[13]);
  assign t[332] = (x[13]);
  assign t[333] = (x[16]);
  assign t[334] = (x[16]);
  assign t[335] = (x[19]);
  assign t[336] = (x[19]);
  assign t[337] = (x[22]);
  assign t[338] = (x[22]);
  assign t[339] = (x[25]);
  assign t[33] = t[8] ? t[53] : t[194];
  assign t[340] = (x[25]);
  assign t[341] = (x[28]);
  assign t[342] = (x[28]);
  assign t[343] = (x[31]);
  assign t[344] = (x[31]);
  assign t[345] = (x[34]);
  assign t[346] = (x[34]);
  assign t[347] = (x[37]);
  assign t[348] = (x[37]);
  assign t[349] = (x[40]);
  assign t[34] = t[195] ^ t[54];
  assign t[350] = (x[40]);
  assign t[351] = (x[43]);
  assign t[352] = (x[43]);
  assign t[353] = (x[48]);
  assign t[354] = (x[48]);
  assign t[355] = (x[51]);
  assign t[356] = (x[51]);
  assign t[357] = (x[54]);
  assign t[358] = (x[54]);
  assign t[359] = (x[57]);
  assign t[35] = ~(t[55]);
  assign t[360] = (x[57]);
  assign t[361] = (x[60]);
  assign t[362] = (x[60]);
  assign t[363] = (x[63]);
  assign t[364] = (x[63]);
  assign t[365] = (x[66]);
  assign t[366] = (x[66]);
  assign t[367] = (x[73]);
  assign t[368] = (x[73]);
  assign t[369] = (x[76]);
  assign t[36] = t[196] ^ t[56];
  assign t[370] = (x[76]);
  assign t[371] = (x[83]);
  assign t[372] = (x[83]);
  assign t[373] = (x[86]);
  assign t[374] = (x[86]);
  assign t[375] = (x[89]);
  assign t[376] = (x[89]);
  assign t[377] = (x[98]);
  assign t[378] = (x[98]);
  assign t[37] = ~(t[57] ^ t[58]);
  assign t[38] = t[59] ^ t[60];
  assign t[39] = t[41] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~t[62];
  assign t[41] = t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[13] ^ t[68];
  assign t[45] = t[69] ^ t[70];
  assign t[46] = t[55] ^ t[34];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[197] | t[75];
  assign t[4] = t[8] ? t[9] : t[190];
  assign t[50] = ~(t[76]);
  assign t[51] = ~(t[195]);
  assign t[52] = ~(t[77] & t[198]);
  assign t[53] = t[194] ^ t[78];
  assign t[54] = t[8] ? t[79] : t[199];
  assign t[55] = t[193] ^ t[80];
  assign t[56] = t[8] ? t[81] : t[200];
  assign t[57] = t[82] ^ t[83];
  assign t[58] = ~(t[84] ^ t[85]);
  assign t[59] = t[86] ^ t[87];
  assign t[5] = ~(t[10]);
  assign t[60] = t[88] & t[89];
  assign t[61] = t[42] ^ t[90];
  assign t[62] = t[8] ? t[91] : t[201];
  assign t[63] = t[8] ? t[92] : t[202];
  assign t[64] = t[93] & t[94];
  assign t[65] = t[95] & t[96];
  assign t[66] = ~(t[64] ^ t[97]);
  assign t[67] = t[98] ^ t[99];
  assign t[68] = t[100] ^ t[101];
  assign t[69] = t[102] ^ t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[104] & t[105];
  assign t[71] = t[106] ^ t[20];
  assign t[72] = t[107] & t[108];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[203] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[49]);
  assign t[77] = ~(t[196]);
  assign t[78] = t[113] ? x[47] : x[46];
  assign t[79] = t[199] ^ t[114];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[115] : t[204];
  assign t[81] = t[200] ^ t[116];
  assign t[82] = t[117] ^ t[118];
  assign t[83] = t[119] ^ t[120];
  assign t[84] = t[121] ^ t[122];
  assign t[85] = t[123] ^ t[124];
  assign t[86] = t[8] ? t[125] : t[205];
  assign t[87] = t[8] ? t[126] : t[206];
  assign t[88] = ~(t[59] ^ t[127]);
  assign t[89] = t[128] ^ t[129];
  assign t[8] = ~(t[15]);
  assign t[90] = t[130] & t[131];
  assign t[91] = t[201] ^ t[132];
  assign t[92] = t[202] ^ t[133];
  assign t[93] = ~(t[99]);
  assign t[94] = ~(t[134]);
  assign t[95] = ~(t[40]);
  assign t[96] = t[135];
  assign t[97] = t[23] ^ t[134];
  assign t[98] = t[134] ^ t[41];
  assign t[99] = t[96] ^ t[40];
  assign t[9] = t[190] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [116:0] x;
 output y;

 wire [378:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[8] ? t[136] : t[207];
  assign t[101] = t[127] ^ t[60];
  assign t[102] = t[137] ? t[138] : t[208];
  assign t[103] = t[137] ? t[139] : t[209];
  assign t[104] = ~(t[69] ^ t[140]);
  assign t[105] = t[141] ^ t[142];
  assign t[106] = t[143] & t[144];
  assign t[107] = ~(t[106] ^ t[145]);
  assign t[108] = t[19] ^ t[146];
  assign t[109] = ~(t[147] & t[148]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[149] ^ t[210];
  assign t[111] = ~(t[203]);
  assign t[112] = t[150] & t[149];
  assign t[113] = ~(t[50]);
  assign t[114] = t[113] ? x[70] : x[69];
  assign t[115] = t[204] ^ t[151];
  assign t[116] = t[113] ? x[72] : x[71];
  assign t[117] = t[102] ^ t[123];
  assign t[118] = t[152] & t[142];
  assign t[119] = t[33] ^ t[55];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[153] & t[154];
  assign t[121] = t[128] ^ t[155];
  assign t[122] = t[156] ^ t[90];
  assign t[123] = t[137] ? t[157] : t[211];
  assign t[124] = t[140] ^ t[70];
  assign t[125] = t[205] ^ t[158];
  assign t[126] = t[206] ^ t[159];
  assign t[127] = t[160] ^ t[161];
  assign t[128] = t[87] ^ t[100];
  assign t[129] = t[8] ? t[162] : t[212];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = ~(t[156] ^ t[42]);
  assign t[131] = t[23] ^ t[96];
  assign t[132] = t[113] ? x[80] : x[79];
  assign t[133] = t[76] ? x[82] : x[81];
  assign t[134] = t[163];
  assign t[135] = t[8] ? t[164] : t[213];
  assign t[136] = t[207] ^ t[165];
  assign t[137] = ~(t[15]);
  assign t[138] = t[208] ^ t[166];
  assign t[139] = t[209] ^ t[167];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[168] ^ t[118];
  assign t[141] = t[103] ^ t[123];
  assign t[142] = t[137] ? t[169] : t[214];
  assign t[143] = ~(t[146]);
  assign t[144] = ~(t[33]);
  assign t[145] = t[46] ^ t[33];
  assign t[146] = t[36] ^ t[55];
  assign t[147] = ~(t[150] | t[149]);
  assign t[148] = ~(t[170] | t[111]);
  assign t[149] = ~(t[215]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[210]);
  assign t[151] = t[113] ? x[93] : x[92];
  assign t[152] = ~(t[103]);
  assign t[153] = ~(t[119] ^ t[71]);
  assign t[154] = t[46] ^ t[36];
  assign t[155] = t[127] ^ t[171];
  assign t[156] = t[134] ^ t[40];
  assign t[157] = t[211] ^ t[172];
  assign t[158] = t[28] ? x[95] : x[94];
  assign t[159] = t[28] ? x[97] : x[96];
  assign t[15] = ~(t[27]);
  assign t[160] = t[173] & t[174];
  assign t[161] = t[175] & t[129];
  assign t[162] = t[212] ^ t[176];
  assign t[163] = t[8] ? t[177] : t[216];
  assign t[164] = t[213] ^ t[178];
  assign t[165] = t[76] ? x[102] : x[101];
  assign t[166] = t[179] ? x[104] : x[103];
  assign t[167] = t[179] ? x[106] : x[105];
  assign t[168] = t[180] & t[181];
  assign t[169] = t[214] ^ t[182];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[197]);
  assign t[171] = t[183] & t[184];
  assign t[172] = t[179] ? x[108] : x[107];
  assign t[173] = ~(t[185]);
  assign t[174] = ~(t[86]);
  assign t[175] = ~(t[87]);
  assign t[176] = t[28] ? x[110] : x[109];
  assign t[177] = t[216] ^ t[186];
  assign t[178] = t[76] ? x[112] : x[111];
  assign t[179] = ~(t[50]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[187]);
  assign t[181] = ~(t[102]);
  assign t[182] = t[179] ? x[114] : x[113];
  assign t[183] = ~(t[160] ^ t[188]);
  assign t[184] = t[189] ^ t[185];
  assign t[185] = t[129] ^ t[87];
  assign t[186] = t[76] ? x[116] : x[115];
  assign t[187] = t[142] ^ t[103];
  assign t[188] = t[128] ^ t[86];
  assign t[189] = t[86] ^ t[100];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] & t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = t[244] ^ x[4];
  assign t[218] = t[245] ^ x[9];
  assign t[219] = t[246] ^ x[12];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[15];
  assign t[221] = t[248] ^ x[18];
  assign t[222] = t[249] ^ x[21];
  assign t[223] = t[250] ^ x[24];
  assign t[224] = t[251] ^ x[27];
  assign t[225] = t[252] ^ x[30];
  assign t[226] = t[253] ^ x[33];
  assign t[227] = t[254] ^ x[36];
  assign t[228] = t[255] ^ x[39];
  assign t[229] = t[256] ^ x[42];
  assign t[22] = ~(t[26] ^ t[39]);
  assign t[230] = t[257] ^ x[45];
  assign t[231] = t[258] ^ x[50];
  assign t[232] = t[259] ^ x[53];
  assign t[233] = t[260] ^ x[56];
  assign t[234] = t[261] ^ x[59];
  assign t[235] = t[262] ^ x[62];
  assign t[236] = t[263] ^ x[65];
  assign t[237] = t[264] ^ x[68];
  assign t[238] = t[265] ^ x[75];
  assign t[239] = t[266] ^ x[78];
  assign t[23] = t[40] ^ t[41];
  assign t[240] = t[267] ^ x[85];
  assign t[241] = t[268] ^ x[88];
  assign t[242] = t[269] ^ x[91];
  assign t[243] = t[270] ^ x[100];
  assign t[244] = (t[271] & ~t[272]);
  assign t[245] = (t[273] & ~t[274]);
  assign t[246] = (t[275] & ~t[276]);
  assign t[247] = (t[277] & ~t[278]);
  assign t[248] = (t[279] & ~t[280]);
  assign t[249] = (t[281] & ~t[282]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[283] & ~t[284]);
  assign t[251] = (t[285] & ~t[286]);
  assign t[252] = (t[287] & ~t[288]);
  assign t[253] = (t[289] & ~t[290]);
  assign t[254] = (t[291] & ~t[292]);
  assign t[255] = (t[293] & ~t[294]);
  assign t[256] = (t[295] & ~t[296]);
  assign t[257] = (t[297] & ~t[298]);
  assign t[258] = (t[299] & ~t[300]);
  assign t[259] = (t[301] & ~t[302]);
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[260] = (t[303] & ~t[304]);
  assign t[261] = (t[305] & ~t[306]);
  assign t[262] = (t[307] & ~t[308]);
  assign t[263] = (t[309] & ~t[310]);
  assign t[264] = (t[311] & ~t[312]);
  assign t[265] = (t[313] & ~t[314]);
  assign t[266] = (t[315] & ~t[316]);
  assign t[267] = (t[317] & ~t[318]);
  assign t[268] = (t[319] & ~t[320]);
  assign t[269] = (t[321] & ~t[322]);
  assign t[26] = t[46] ^ t[47];
  assign t[270] = (t[323] & ~t[324]);
  assign t[271] = t[325] ^ x[4];
  assign t[272] = t[326] ^ x[3];
  assign t[273] = t[327] ^ x[9];
  assign t[274] = t[328] ^ x[8];
  assign t[275] = t[329] ^ x[12];
  assign t[276] = t[330] ^ x[11];
  assign t[277] = t[331] ^ x[15];
  assign t[278] = t[332] ^ x[14];
  assign t[279] = t[333] ^ x[18];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[17];
  assign t[281] = t[335] ^ x[21];
  assign t[282] = t[336] ^ x[20];
  assign t[283] = t[337] ^ x[24];
  assign t[284] = t[338] ^ x[23];
  assign t[285] = t[339] ^ x[27];
  assign t[286] = t[340] ^ x[26];
  assign t[287] = t[341] ^ x[30];
  assign t[288] = t[342] ^ x[29];
  assign t[289] = t[343] ^ x[33];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[32];
  assign t[291] = t[345] ^ x[36];
  assign t[292] = t[346] ^ x[35];
  assign t[293] = t[347] ^ x[39];
  assign t[294] = t[348] ^ x[38];
  assign t[295] = t[349] ^ x[42];
  assign t[296] = t[350] ^ x[41];
  assign t[297] = t[351] ^ x[45];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[50];
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[49];
  assign t[301] = t[355] ^ x[53];
  assign t[302] = t[356] ^ x[52];
  assign t[303] = t[357] ^ x[56];
  assign t[304] = t[358] ^ x[55];
  assign t[305] = t[359] ^ x[59];
  assign t[306] = t[360] ^ x[58];
  assign t[307] = t[361] ^ x[62];
  assign t[308] = t[362] ^ x[61];
  assign t[309] = t[363] ^ x[65];
  assign t[30] = ~(t[192]);
  assign t[310] = t[364] ^ x[64];
  assign t[311] = t[365] ^ x[68];
  assign t[312] = t[366] ^ x[67];
  assign t[313] = t[367] ^ x[75];
  assign t[314] = t[368] ^ x[74];
  assign t[315] = t[369] ^ x[78];
  assign t[316] = t[370] ^ x[77];
  assign t[317] = t[371] ^ x[85];
  assign t[318] = t[372] ^ x[84];
  assign t[319] = t[373] ^ x[88];
  assign t[31] = ~(t[193]);
  assign t[320] = t[374] ^ x[87];
  assign t[321] = t[375] ^ x[91];
  assign t[322] = t[376] ^ x[90];
  assign t[323] = t[377] ^ x[100];
  assign t[324] = t[378] ^ x[99];
  assign t[325] = (x[2]);
  assign t[326] = (x[2]);
  assign t[327] = (x[7]);
  assign t[328] = (x[7]);
  assign t[329] = (x[10]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[10]);
  assign t[331] = (x[13]);
  assign t[332] = (x[13]);
  assign t[333] = (x[16]);
  assign t[334] = (x[16]);
  assign t[335] = (x[19]);
  assign t[336] = (x[19]);
  assign t[337] = (x[22]);
  assign t[338] = (x[22]);
  assign t[339] = (x[25]);
  assign t[33] = t[8] ? t[53] : t[194];
  assign t[340] = (x[25]);
  assign t[341] = (x[28]);
  assign t[342] = (x[28]);
  assign t[343] = (x[31]);
  assign t[344] = (x[31]);
  assign t[345] = (x[34]);
  assign t[346] = (x[34]);
  assign t[347] = (x[37]);
  assign t[348] = (x[37]);
  assign t[349] = (x[40]);
  assign t[34] = t[195] ^ t[54];
  assign t[350] = (x[40]);
  assign t[351] = (x[43]);
  assign t[352] = (x[43]);
  assign t[353] = (x[48]);
  assign t[354] = (x[48]);
  assign t[355] = (x[51]);
  assign t[356] = (x[51]);
  assign t[357] = (x[54]);
  assign t[358] = (x[54]);
  assign t[359] = (x[57]);
  assign t[35] = ~(t[55]);
  assign t[360] = (x[57]);
  assign t[361] = (x[60]);
  assign t[362] = (x[60]);
  assign t[363] = (x[63]);
  assign t[364] = (x[63]);
  assign t[365] = (x[66]);
  assign t[366] = (x[66]);
  assign t[367] = (x[73]);
  assign t[368] = (x[73]);
  assign t[369] = (x[76]);
  assign t[36] = t[196] ^ t[56];
  assign t[370] = (x[76]);
  assign t[371] = (x[83]);
  assign t[372] = (x[83]);
  assign t[373] = (x[86]);
  assign t[374] = (x[86]);
  assign t[375] = (x[89]);
  assign t[376] = (x[89]);
  assign t[377] = (x[98]);
  assign t[378] = (x[98]);
  assign t[37] = ~(t[57] ^ t[58]);
  assign t[38] = t[59] ^ t[60];
  assign t[39] = t[41] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~t[62];
  assign t[41] = t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[13] ^ t[68];
  assign t[45] = t[69] ^ t[70];
  assign t[46] = t[55] ^ t[34];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[197] | t[75];
  assign t[4] = t[8] ? t[9] : t[190];
  assign t[50] = ~(t[76]);
  assign t[51] = ~(t[195]);
  assign t[52] = ~(t[77] & t[198]);
  assign t[53] = t[194] ^ t[78];
  assign t[54] = t[8] ? t[79] : t[199];
  assign t[55] = t[193] ^ t[80];
  assign t[56] = t[8] ? t[81] : t[200];
  assign t[57] = t[82] ^ t[83];
  assign t[58] = ~(t[84] ^ t[85]);
  assign t[59] = t[86] ^ t[87];
  assign t[5] = ~(t[10]);
  assign t[60] = t[88] & t[89];
  assign t[61] = t[42] ^ t[90];
  assign t[62] = t[8] ? t[91] : t[201];
  assign t[63] = t[8] ? t[92] : t[202];
  assign t[64] = t[93] & t[94];
  assign t[65] = t[95] & t[96];
  assign t[66] = ~(t[64] ^ t[97]);
  assign t[67] = t[98] ^ t[99];
  assign t[68] = t[100] ^ t[101];
  assign t[69] = t[102] ^ t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[104] & t[105];
  assign t[71] = t[106] ^ t[20];
  assign t[72] = t[107] & t[108];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[203] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[49]);
  assign t[77] = ~(t[196]);
  assign t[78] = t[113] ? x[47] : x[46];
  assign t[79] = t[199] ^ t[114];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[115] : t[204];
  assign t[81] = t[200] ^ t[116];
  assign t[82] = t[117] ^ t[118];
  assign t[83] = t[119] ^ t[120];
  assign t[84] = t[121] ^ t[122];
  assign t[85] = t[123] ^ t[124];
  assign t[86] = t[8] ? t[125] : t[205];
  assign t[87] = t[8] ? t[126] : t[206];
  assign t[88] = ~(t[59] ^ t[127]);
  assign t[89] = t[128] ^ t[129];
  assign t[8] = ~(t[15]);
  assign t[90] = t[130] & t[131];
  assign t[91] = t[201] ^ t[132];
  assign t[92] = t[202] ^ t[133];
  assign t[93] = ~(t[99]);
  assign t[94] = ~(t[134]);
  assign t[95] = ~(t[40]);
  assign t[96] = t[135];
  assign t[97] = t[23] ^ t[134];
  assign t[98] = t[134] ^ t[41];
  assign t[99] = t[96] ^ t[40];
  assign t[9] = t[190] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind106(x, y);
 input [116:0] x;
 output y;

 wire [396:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[8] ? t[137] : t[222];
  assign t[101] = t[138] ^ t[121];
  assign t[102] = t[139] & t[140];
  assign t[103] = t[8] ? t[141] : t[223];
  assign t[104] = t[142] ^ t[143];
  assign t[105] = t[42] ^ t[144];
  assign t[106] = t[145] ^ t[146];
  assign t[107] = t[8] ? t[147] : t[224];
  assign t[108] = ~(t[72] ^ t[101]);
  assign t[109] = t[66] ^ t[148];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[149] & t[150];
  assign t[111] = ~(t[151] & t[152]);
  assign t[112] = t[153] ^ t[225];
  assign t[113] = ~(t[217]);
  assign t[114] = t[154] & t[153];
  assign t[115] = t[100] ^ t[155];
  assign t[116] = t[156] ^ t[157];
  assign t[117] = t[158] & t[159];
  assign t[118] = t[157] ^ t[145];
  assign t[119] = t[160] ^ t[161];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[107] ^ t[100];
  assign t[121] = t[162] & t[148];
  assign t[122] = t[163] ? x[59] : x[58];
  assign t[123] = t[219] ^ t[164];
  assign t[124] = t[165] & t[166];
  assign t[125] = t[167] & t[88];
  assign t[126] = t[8] ? t[168] : t[226];
  assign t[127] = t[220] ^ t[169];
  assign t[128] = ~(t[131]);
  assign t[129] = ~(t[96]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[37] ^ t[96];
  assign t[131] = t[98] ^ t[59];
  assign t[132] = t[79] ? x[64] : x[63];
  assign t[133] = t[96] ^ t[59];
  assign t[134] = t[8] ? t[170] : t[227];
  assign t[135] = t[8] ? t[171] : t[228];
  assign t[136] = t[221] ^ t[172];
  assign t[137] = t[222] ^ t[173];
  assign t[138] = t[174] & t[175];
  assign t[139] = ~(t[138] ^ t[176]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[120] ^ t[177];
  assign t[141] = t[223] ^ t[178];
  assign t[142] = t[156] ^ t[145];
  assign t[143] = t[179] & t[180];
  assign t[144] = t[133] ^ t[63];
  assign t[145] = t[181] ? t[182] : t[229];
  assign t[146] = t[160] ^ t[117];
  assign t[147] = t[224] ^ t[183];
  assign t[148] = t[8] ? t[184] : t[230];
  assign t[149] = ~(t[124] ^ t[185]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[186] ^ t[187];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[188] | t[113]);
  assign t[153] = ~(t[231]);
  assign t[154] = ~(t[225]);
  assign t[155] = t[101] ^ t[73];
  assign t[156] = t[181] ? t[189] : t[232];
  assign t[157] = t[181] ? t[190] : t[233];
  assign t[158] = ~(t[116] ^ t[160]);
  assign t[159] = t[118] ^ t[180];
  assign t[15] = ~(t[27]);
  assign t[160] = t[191] ^ t[143];
  assign t[161] = t[192] & t[193];
  assign t[162] = ~(t[99]);
  assign t[163] = ~(t[49]);
  assign t[164] = t[163] ? x[87] : x[86];
  assign t[165] = ~(t[187]);
  assign t[166] = ~(t[55]);
  assign t[167] = ~(t[56]);
  assign t[168] = t[226] ^ t[194];
  assign t[169] = t[163] ? x[89] : x[88];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[227] ^ t[195];
  assign t[171] = t[228] ^ t[196];
  assign t[172] = t[28] ? x[91] : x[90];
  assign t[173] = t[79] ? x[93] : x[92];
  assign t[174] = ~(t[177]);
  assign t[175] = ~(t[107]);
  assign t[176] = t[66] ^ t[107];
  assign t[177] = t[148] ^ t[99];
  assign t[178] = t[163] ? x[95] : x[94];
  assign t[179] = ~(t[157]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[181] ? t[197] : t[234];
  assign t[181] = ~(t[15]);
  assign t[182] = t[229] ^ t[198];
  assign t[183] = t[28] ? x[100] : x[99];
  assign t[184] = t[230] ^ t[199];
  assign t[185] = t[74] ^ t[55];
  assign t[186] = t[55] ^ t[68];
  assign t[187] = t[88] ^ t[56];
  assign t[188] = ~(t[212]);
  assign t[189] = t[232] ^ t[200];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[233] ^ t[201];
  assign t[191] = t[202] & t[203];
  assign t[192] = ~(t[191] ^ t[204]);
  assign t[193] = t[142] ^ t[205];
  assign t[194] = t[163] ? x[102] : x[101];
  assign t[195] = t[79] ? x[104] : x[103];
  assign t[196] = t[79] ? x[106] : x[105];
  assign t[197] = t[234] ^ t[206];
  assign t[198] = t[207] ? x[108] : x[107];
  assign t[199] = t[28] ? x[110] : x[109];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[207] ? x[112] : x[111];
  assign t[201] = t[207] ? x[114] : x[113];
  assign t[202] = ~(t[205]);
  assign t[203] = ~(t[156]);
  assign t[204] = t[118] ^ t[156];
  assign t[205] = t[180] ^ t[157];
  assign t[206] = t[207] ? x[116] : x[115];
  assign t[207] = ~(t[49]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = t[262] ^ x[4];
  assign t[236] = t[263] ^ x[9];
  assign t[237] = t[264] ^ x[12];
  assign t[238] = t[265] ^ x[15];
  assign t[239] = t[266] ^ x[18];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[21];
  assign t[241] = t[268] ^ x[24];
  assign t[242] = t[269] ^ x[27];
  assign t[243] = t[270] ^ x[30];
  assign t[244] = t[271] ^ x[33];
  assign t[245] = t[272] ^ x[36];
  assign t[246] = t[273] ^ x[39];
  assign t[247] = t[274] ^ x[42];
  assign t[248] = t[275] ^ x[45];
  assign t[249] = t[276] ^ x[48];
  assign t[24] = ~(t[33] ^ t[43]);
  assign t[250] = t[277] ^ x[51];
  assign t[251] = t[278] ^ x[54];
  assign t[252] = t[279] ^ x[57];
  assign t[253] = t[280] ^ x[62];
  assign t[254] = t[281] ^ x[67];
  assign t[255] = t[282] ^ x[70];
  assign t[256] = t[283] ^ x[73];
  assign t[257] = t[284] ^ x[76];
  assign t[258] = t[285] ^ x[79];
  assign t[259] = t[286] ^ x[82];
  assign t[25] = t[44] ^ t[45];
  assign t[260] = t[287] ^ x[85];
  assign t[261] = t[288] ^ x[98];
  assign t[262] = (t[289] & ~t[290]);
  assign t[263] = (t[291] & ~t[292]);
  assign t[264] = (t[293] & ~t[294]);
  assign t[265] = (t[295] & ~t[296]);
  assign t[266] = (t[297] & ~t[298]);
  assign t[267] = (t[299] & ~t[300]);
  assign t[268] = (t[301] & ~t[302]);
  assign t[269] = (t[303] & ~t[304]);
  assign t[26] = ~(t[46] ^ t[22]);
  assign t[270] = (t[305] & ~t[306]);
  assign t[271] = (t[307] & ~t[308]);
  assign t[272] = (t[309] & ~t[310]);
  assign t[273] = (t[311] & ~t[312]);
  assign t[274] = (t[313] & ~t[314]);
  assign t[275] = (t[315] & ~t[316]);
  assign t[276] = (t[317] & ~t[318]);
  assign t[277] = (t[319] & ~t[320]);
  assign t[278] = (t[321] & ~t[322]);
  assign t[279] = (t[323] & ~t[324]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[325] & ~t[326]);
  assign t[281] = (t[327] & ~t[328]);
  assign t[282] = (t[329] & ~t[330]);
  assign t[283] = (t[331] & ~t[332]);
  assign t[284] = (t[333] & ~t[334]);
  assign t[285] = (t[335] & ~t[336]);
  assign t[286] = (t[337] & ~t[338]);
  assign t[287] = (t[339] & ~t[340]);
  assign t[288] = (t[341] & ~t[342]);
  assign t[289] = t[343] ^ x[4];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[3];
  assign t[291] = t[345] ^ x[9];
  assign t[292] = t[346] ^ x[8];
  assign t[293] = t[347] ^ x[12];
  assign t[294] = t[348] ^ x[11];
  assign t[295] = t[349] ^ x[15];
  assign t[296] = t[350] ^ x[14];
  assign t[297] = t[351] ^ x[18];
  assign t[298] = t[352] ^ x[17];
  assign t[299] = t[353] ^ x[21];
  assign t[29] = ~(t[209]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[20];
  assign t[301] = t[355] ^ x[24];
  assign t[302] = t[356] ^ x[23];
  assign t[303] = t[357] ^ x[27];
  assign t[304] = t[358] ^ x[26];
  assign t[305] = t[359] ^ x[30];
  assign t[306] = t[360] ^ x[29];
  assign t[307] = t[361] ^ x[33];
  assign t[308] = t[362] ^ x[32];
  assign t[309] = t[363] ^ x[36];
  assign t[30] = ~(t[210]);
  assign t[310] = t[364] ^ x[35];
  assign t[311] = t[365] ^ x[39];
  assign t[312] = t[366] ^ x[38];
  assign t[313] = t[367] ^ x[42];
  assign t[314] = t[368] ^ x[41];
  assign t[315] = t[369] ^ x[45];
  assign t[316] = t[370] ^ x[44];
  assign t[317] = t[371] ^ x[48];
  assign t[318] = t[372] ^ x[47];
  assign t[319] = t[373] ^ x[51];
  assign t[31] = ~(t[211]);
  assign t[320] = t[374] ^ x[50];
  assign t[321] = t[375] ^ x[54];
  assign t[322] = t[376] ^ x[53];
  assign t[323] = t[377] ^ x[57];
  assign t[324] = t[378] ^ x[56];
  assign t[325] = t[379] ^ x[62];
  assign t[326] = t[380] ^ x[61];
  assign t[327] = t[381] ^ x[67];
  assign t[328] = t[382] ^ x[66];
  assign t[329] = t[383] ^ x[70];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[69];
  assign t[331] = t[385] ^ x[73];
  assign t[332] = t[386] ^ x[72];
  assign t[333] = t[387] ^ x[76];
  assign t[334] = t[388] ^ x[75];
  assign t[335] = t[389] ^ x[79];
  assign t[336] = t[390] ^ x[78];
  assign t[337] = t[391] ^ x[82];
  assign t[338] = t[392] ^ x[81];
  assign t[339] = t[393] ^ x[85];
  assign t[33] = ~(t[52] ^ t[46]);
  assign t[340] = t[394] ^ x[84];
  assign t[341] = t[395] ^ x[98];
  assign t[342] = t[396] ^ x[97];
  assign t[343] = (x[2]);
  assign t[344] = (x[2]);
  assign t[345] = (x[7]);
  assign t[346] = (x[7]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[49]);
  assign t[374] = (x[49]);
  assign t[375] = (x[52]);
  assign t[376] = (x[52]);
  assign t[377] = (x[55]);
  assign t[378] = (x[55]);
  assign t[379] = (x[60]);
  assign t[37] = t[59] ^ t[39];
  assign t[380] = (x[60]);
  assign t[381] = (x[65]);
  assign t[382] = (x[65]);
  assign t[383] = (x[68]);
  assign t[384] = (x[68]);
  assign t[385] = (x[71]);
  assign t[386] = (x[71]);
  assign t[387] = (x[74]);
  assign t[388] = (x[74]);
  assign t[389] = (x[77]);
  assign t[38] = t[60] ^ t[61];
  assign t[390] = (x[77]);
  assign t[391] = (x[80]);
  assign t[392] = (x[80]);
  assign t[393] = (x[83]);
  assign t[394] = (x[83]);
  assign t[395] = (x[96]);
  assign t[396] = (x[96]);
  assign t[39] = t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[60] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = ~(t[70] ^ t[71]);
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = t[212] | t[78];
  assign t[49] = ~(t[79]);
  assign t[4] = t[8] ? t[9] : t[208];
  assign t[50] = ~(t[213]);
  assign t[51] = ~(t[80] & t[214]);
  assign t[52] = ~(t[81] ^ t[82]);
  assign t[53] = t[83] ^ t[84];
  assign t[54] = ~(t[43] ^ t[22]);
  assign t[55] = t[8] ? t[85] : t[215];
  assign t[56] = t[211] ^ t[86];
  assign t[57] = ~(t[35] ^ t[87]);
  assign t[58] = t[74] ^ t[88];
  assign t[59] = ~t[89];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[65];
  assign t[61] = t[91] & t[92];
  assign t[62] = t[8] ? t[93] : t[216];
  assign t[63] = t[94] & t[95];
  assign t[64] = t[96] ^ t[39];
  assign t[65] = t[97] & t[98];
  assign t[66] = t[99] ^ t[100];
  assign t[67] = t[101] ^ t[102];
  assign t[68] = t[213] ^ t[103];
  assign t[69] = t[87] ^ t[36];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[104] ^ t[20];
  assign t[71] = ~(t[105] ^ t[106]);
  assign t[72] = t[107] ^ t[99];
  assign t[73] = t[108] & t[109];
  assign t[74] = t[56] ^ t[68];
  assign t[75] = t[87] ^ t[110];
  assign t[76] = ~(t[78] & t[111]);
  assign t[77] = ~(t[217] ^ t[112]);
  assign t[78] = ~(t[113] & t[114]);
  assign t[79] = ~(t[48]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[218]);
  assign t[81] = t[21] ^ t[115];
  assign t[82] = t[116] ^ t[117];
  assign t[83] = t[118] ^ t[119];
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[215] ^ t[122];
  assign t[86] = t[8] ? t[123] : t[219];
  assign t[87] = t[124] ^ t[125];
  assign t[88] = t[218] ^ t[126];
  assign t[89] = t[8] ? t[127] : t[220];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] & t[129];
  assign t[91] = ~(t[90] ^ t[130]);
  assign t[92] = t[64] ^ t[131];
  assign t[93] = t[216] ^ t[132];
  assign t[94] = ~(t[133] ^ t[60]);
  assign t[95] = t[37] ^ t[98];
  assign t[96] = t[134];
  assign t[97] = ~(t[59]);
  assign t[98] = t[135];
  assign t[99] = t[8] ? t[136] : t[221];
  assign t[9] = t[208] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [116:0] x;
 output y;

 wire [396:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[8] ? t[137] : t[222];
  assign t[101] = t[138] ^ t[121];
  assign t[102] = t[139] & t[140];
  assign t[103] = t[8] ? t[141] : t[223];
  assign t[104] = t[142] ^ t[143];
  assign t[105] = t[42] ^ t[144];
  assign t[106] = t[145] ^ t[146];
  assign t[107] = t[8] ? t[147] : t[224];
  assign t[108] = ~(t[72] ^ t[101]);
  assign t[109] = t[66] ^ t[148];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[149] & t[150];
  assign t[111] = ~(t[151] & t[152]);
  assign t[112] = t[153] ^ t[225];
  assign t[113] = ~(t[217]);
  assign t[114] = t[154] & t[153];
  assign t[115] = t[100] ^ t[155];
  assign t[116] = t[156] ^ t[157];
  assign t[117] = t[158] & t[159];
  assign t[118] = t[157] ^ t[145];
  assign t[119] = t[160] ^ t[161];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[107] ^ t[100];
  assign t[121] = t[162] & t[148];
  assign t[122] = t[163] ? x[59] : x[58];
  assign t[123] = t[219] ^ t[164];
  assign t[124] = t[165] & t[166];
  assign t[125] = t[167] & t[88];
  assign t[126] = t[8] ? t[168] : t[226];
  assign t[127] = t[220] ^ t[169];
  assign t[128] = ~(t[131]);
  assign t[129] = ~(t[96]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[37] ^ t[96];
  assign t[131] = t[98] ^ t[59];
  assign t[132] = t[79] ? x[64] : x[63];
  assign t[133] = t[96] ^ t[59];
  assign t[134] = t[8] ? t[170] : t[227];
  assign t[135] = t[8] ? t[171] : t[228];
  assign t[136] = t[221] ^ t[172];
  assign t[137] = t[222] ^ t[173];
  assign t[138] = t[174] & t[175];
  assign t[139] = ~(t[138] ^ t[176]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[120] ^ t[177];
  assign t[141] = t[223] ^ t[178];
  assign t[142] = t[156] ^ t[145];
  assign t[143] = t[179] & t[180];
  assign t[144] = t[133] ^ t[63];
  assign t[145] = t[181] ? t[182] : t[229];
  assign t[146] = t[160] ^ t[117];
  assign t[147] = t[224] ^ t[183];
  assign t[148] = t[8] ? t[184] : t[230];
  assign t[149] = ~(t[124] ^ t[185]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[186] ^ t[187];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[188] | t[113]);
  assign t[153] = ~(t[231]);
  assign t[154] = ~(t[225]);
  assign t[155] = t[101] ^ t[73];
  assign t[156] = t[181] ? t[189] : t[232];
  assign t[157] = t[181] ? t[190] : t[233];
  assign t[158] = ~(t[116] ^ t[160]);
  assign t[159] = t[118] ^ t[180];
  assign t[15] = ~(t[27]);
  assign t[160] = t[191] ^ t[143];
  assign t[161] = t[192] & t[193];
  assign t[162] = ~(t[99]);
  assign t[163] = ~(t[49]);
  assign t[164] = t[163] ? x[87] : x[86];
  assign t[165] = ~(t[187]);
  assign t[166] = ~(t[55]);
  assign t[167] = ~(t[56]);
  assign t[168] = t[226] ^ t[194];
  assign t[169] = t[163] ? x[89] : x[88];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[227] ^ t[195];
  assign t[171] = t[228] ^ t[196];
  assign t[172] = t[28] ? x[91] : x[90];
  assign t[173] = t[79] ? x[93] : x[92];
  assign t[174] = ~(t[177]);
  assign t[175] = ~(t[107]);
  assign t[176] = t[66] ^ t[107];
  assign t[177] = t[148] ^ t[99];
  assign t[178] = t[163] ? x[95] : x[94];
  assign t[179] = ~(t[157]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[181] ? t[197] : t[234];
  assign t[181] = ~(t[15]);
  assign t[182] = t[229] ^ t[198];
  assign t[183] = t[28] ? x[100] : x[99];
  assign t[184] = t[230] ^ t[199];
  assign t[185] = t[74] ^ t[55];
  assign t[186] = t[55] ^ t[68];
  assign t[187] = t[88] ^ t[56];
  assign t[188] = ~(t[212]);
  assign t[189] = t[232] ^ t[200];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[233] ^ t[201];
  assign t[191] = t[202] & t[203];
  assign t[192] = ~(t[191] ^ t[204]);
  assign t[193] = t[142] ^ t[205];
  assign t[194] = t[163] ? x[102] : x[101];
  assign t[195] = t[79] ? x[104] : x[103];
  assign t[196] = t[79] ? x[106] : x[105];
  assign t[197] = t[234] ^ t[206];
  assign t[198] = t[207] ? x[108] : x[107];
  assign t[199] = t[28] ? x[110] : x[109];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[207] ? x[112] : x[111];
  assign t[201] = t[207] ? x[114] : x[113];
  assign t[202] = ~(t[205]);
  assign t[203] = ~(t[156]);
  assign t[204] = t[118] ^ t[156];
  assign t[205] = t[180] ^ t[157];
  assign t[206] = t[207] ? x[116] : x[115];
  assign t[207] = ~(t[49]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = t[262] ^ x[4];
  assign t[236] = t[263] ^ x[9];
  assign t[237] = t[264] ^ x[12];
  assign t[238] = t[265] ^ x[15];
  assign t[239] = t[266] ^ x[18];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[21];
  assign t[241] = t[268] ^ x[24];
  assign t[242] = t[269] ^ x[27];
  assign t[243] = t[270] ^ x[30];
  assign t[244] = t[271] ^ x[33];
  assign t[245] = t[272] ^ x[36];
  assign t[246] = t[273] ^ x[39];
  assign t[247] = t[274] ^ x[42];
  assign t[248] = t[275] ^ x[45];
  assign t[249] = t[276] ^ x[48];
  assign t[24] = ~(t[33] ^ t[43]);
  assign t[250] = t[277] ^ x[51];
  assign t[251] = t[278] ^ x[54];
  assign t[252] = t[279] ^ x[57];
  assign t[253] = t[280] ^ x[62];
  assign t[254] = t[281] ^ x[67];
  assign t[255] = t[282] ^ x[70];
  assign t[256] = t[283] ^ x[73];
  assign t[257] = t[284] ^ x[76];
  assign t[258] = t[285] ^ x[79];
  assign t[259] = t[286] ^ x[82];
  assign t[25] = t[44] ^ t[45];
  assign t[260] = t[287] ^ x[85];
  assign t[261] = t[288] ^ x[98];
  assign t[262] = (t[289] & ~t[290]);
  assign t[263] = (t[291] & ~t[292]);
  assign t[264] = (t[293] & ~t[294]);
  assign t[265] = (t[295] & ~t[296]);
  assign t[266] = (t[297] & ~t[298]);
  assign t[267] = (t[299] & ~t[300]);
  assign t[268] = (t[301] & ~t[302]);
  assign t[269] = (t[303] & ~t[304]);
  assign t[26] = ~(t[46] ^ t[22]);
  assign t[270] = (t[305] & ~t[306]);
  assign t[271] = (t[307] & ~t[308]);
  assign t[272] = (t[309] & ~t[310]);
  assign t[273] = (t[311] & ~t[312]);
  assign t[274] = (t[313] & ~t[314]);
  assign t[275] = (t[315] & ~t[316]);
  assign t[276] = (t[317] & ~t[318]);
  assign t[277] = (t[319] & ~t[320]);
  assign t[278] = (t[321] & ~t[322]);
  assign t[279] = (t[323] & ~t[324]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[325] & ~t[326]);
  assign t[281] = (t[327] & ~t[328]);
  assign t[282] = (t[329] & ~t[330]);
  assign t[283] = (t[331] & ~t[332]);
  assign t[284] = (t[333] & ~t[334]);
  assign t[285] = (t[335] & ~t[336]);
  assign t[286] = (t[337] & ~t[338]);
  assign t[287] = (t[339] & ~t[340]);
  assign t[288] = (t[341] & ~t[342]);
  assign t[289] = t[343] ^ x[4];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[3];
  assign t[291] = t[345] ^ x[9];
  assign t[292] = t[346] ^ x[8];
  assign t[293] = t[347] ^ x[12];
  assign t[294] = t[348] ^ x[11];
  assign t[295] = t[349] ^ x[15];
  assign t[296] = t[350] ^ x[14];
  assign t[297] = t[351] ^ x[18];
  assign t[298] = t[352] ^ x[17];
  assign t[299] = t[353] ^ x[21];
  assign t[29] = ~(t[209]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[20];
  assign t[301] = t[355] ^ x[24];
  assign t[302] = t[356] ^ x[23];
  assign t[303] = t[357] ^ x[27];
  assign t[304] = t[358] ^ x[26];
  assign t[305] = t[359] ^ x[30];
  assign t[306] = t[360] ^ x[29];
  assign t[307] = t[361] ^ x[33];
  assign t[308] = t[362] ^ x[32];
  assign t[309] = t[363] ^ x[36];
  assign t[30] = ~(t[210]);
  assign t[310] = t[364] ^ x[35];
  assign t[311] = t[365] ^ x[39];
  assign t[312] = t[366] ^ x[38];
  assign t[313] = t[367] ^ x[42];
  assign t[314] = t[368] ^ x[41];
  assign t[315] = t[369] ^ x[45];
  assign t[316] = t[370] ^ x[44];
  assign t[317] = t[371] ^ x[48];
  assign t[318] = t[372] ^ x[47];
  assign t[319] = t[373] ^ x[51];
  assign t[31] = ~(t[211]);
  assign t[320] = t[374] ^ x[50];
  assign t[321] = t[375] ^ x[54];
  assign t[322] = t[376] ^ x[53];
  assign t[323] = t[377] ^ x[57];
  assign t[324] = t[378] ^ x[56];
  assign t[325] = t[379] ^ x[62];
  assign t[326] = t[380] ^ x[61];
  assign t[327] = t[381] ^ x[67];
  assign t[328] = t[382] ^ x[66];
  assign t[329] = t[383] ^ x[70];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[69];
  assign t[331] = t[385] ^ x[73];
  assign t[332] = t[386] ^ x[72];
  assign t[333] = t[387] ^ x[76];
  assign t[334] = t[388] ^ x[75];
  assign t[335] = t[389] ^ x[79];
  assign t[336] = t[390] ^ x[78];
  assign t[337] = t[391] ^ x[82];
  assign t[338] = t[392] ^ x[81];
  assign t[339] = t[393] ^ x[85];
  assign t[33] = ~(t[52] ^ t[46]);
  assign t[340] = t[394] ^ x[84];
  assign t[341] = t[395] ^ x[98];
  assign t[342] = t[396] ^ x[97];
  assign t[343] = (x[2]);
  assign t[344] = (x[2]);
  assign t[345] = (x[7]);
  assign t[346] = (x[7]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[49]);
  assign t[374] = (x[49]);
  assign t[375] = (x[52]);
  assign t[376] = (x[52]);
  assign t[377] = (x[55]);
  assign t[378] = (x[55]);
  assign t[379] = (x[60]);
  assign t[37] = t[59] ^ t[39];
  assign t[380] = (x[60]);
  assign t[381] = (x[65]);
  assign t[382] = (x[65]);
  assign t[383] = (x[68]);
  assign t[384] = (x[68]);
  assign t[385] = (x[71]);
  assign t[386] = (x[71]);
  assign t[387] = (x[74]);
  assign t[388] = (x[74]);
  assign t[389] = (x[77]);
  assign t[38] = t[60] ^ t[61];
  assign t[390] = (x[77]);
  assign t[391] = (x[80]);
  assign t[392] = (x[80]);
  assign t[393] = (x[83]);
  assign t[394] = (x[83]);
  assign t[395] = (x[96]);
  assign t[396] = (x[96]);
  assign t[39] = t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[60] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = ~(t[70] ^ t[71]);
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = t[212] | t[78];
  assign t[49] = ~(t[79]);
  assign t[4] = t[8] ? t[9] : t[208];
  assign t[50] = ~(t[213]);
  assign t[51] = ~(t[80] & t[214]);
  assign t[52] = ~(t[81] ^ t[82]);
  assign t[53] = t[83] ^ t[84];
  assign t[54] = ~(t[43] ^ t[22]);
  assign t[55] = t[8] ? t[85] : t[215];
  assign t[56] = t[211] ^ t[86];
  assign t[57] = ~(t[35] ^ t[87]);
  assign t[58] = t[74] ^ t[88];
  assign t[59] = ~t[89];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[65];
  assign t[61] = t[91] & t[92];
  assign t[62] = t[8] ? t[93] : t[216];
  assign t[63] = t[94] & t[95];
  assign t[64] = t[96] ^ t[39];
  assign t[65] = t[97] & t[98];
  assign t[66] = t[99] ^ t[100];
  assign t[67] = t[101] ^ t[102];
  assign t[68] = t[213] ^ t[103];
  assign t[69] = t[87] ^ t[36];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[104] ^ t[20];
  assign t[71] = ~(t[105] ^ t[106]);
  assign t[72] = t[107] ^ t[99];
  assign t[73] = t[108] & t[109];
  assign t[74] = t[56] ^ t[68];
  assign t[75] = t[87] ^ t[110];
  assign t[76] = ~(t[78] & t[111]);
  assign t[77] = ~(t[217] ^ t[112]);
  assign t[78] = ~(t[113] & t[114]);
  assign t[79] = ~(t[48]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[218]);
  assign t[81] = t[21] ^ t[115];
  assign t[82] = t[116] ^ t[117];
  assign t[83] = t[118] ^ t[119];
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[215] ^ t[122];
  assign t[86] = t[8] ? t[123] : t[219];
  assign t[87] = t[124] ^ t[125];
  assign t[88] = t[218] ^ t[126];
  assign t[89] = t[8] ? t[127] : t[220];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] & t[129];
  assign t[91] = ~(t[90] ^ t[130]);
  assign t[92] = t[64] ^ t[131];
  assign t[93] = t[216] ^ t[132];
  assign t[94] = ~(t[133] ^ t[60]);
  assign t[95] = t[37] ^ t[98];
  assign t[96] = t[134];
  assign t[97] = ~(t[59]);
  assign t[98] = t[135];
  assign t[99] = t[8] ? t[136] : t[221];
  assign t[9] = t[208] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[134] & t[135];
  assign t[101] = ~(t[99] ^ t[136]);
  assign t[102] = t[137] ^ t[138];
  assign t[103] = t[80] ? x[53] : x[52];
  assign t[104] = t[139] & t[140];
  assign t[105] = t[141] & t[127];
  assign t[106] = t[142] & t[143];
  assign t[107] = t[144];
  assign t[108] = ~t[145];
  assign t[109] = ~(t[70] ^ t[146]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[147] ^ t[148];
  assign t[111] = t[147] ^ t[149];
  assign t[112] = t[150] ^ t[63];
  assign t[113] = t[91] ^ t[41];
  assign t[114] = t[35] ^ t[151];
  assign t[115] = t[152];
  assign t[116] = t[146] ^ t[71];
  assign t[117] = ~(t[153] & t[154]);
  assign t[118] = t[155] ^ t[213];
  assign t[119] = ~(t[209]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[156] & t[155];
  assign t[121] = t[157] ? x[58] : x[57];
  assign t[122] = t[157] ? x[60] : x[59];
  assign t[123] = t[8] ? t[158] : t[214];
  assign t[124] = t[8] ? t[159] : t[215];
  assign t[125] = t[211] ^ t[160];
  assign t[126] = t[212] ^ t[161];
  assign t[127] = t[8] ? t[162] : t[216];
  assign t[128] = t[163] ? x[71] : x[70];
  assign t[129] = ~(t[112] ^ t[64]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[39] ^ t[135];
  assign t[131] = t[163] ? x[73] : x[72];
  assign t[132] = ~(t[138]);
  assign t[133] = ~(t[150]);
  assign t[134] = ~(t[63]);
  assign t[135] = t[95] ? t[164] : t[217];
  assign t[136] = t[39] ^ t[150];
  assign t[137] = t[150] ^ t[61];
  assign t[138] = t[135] ^ t[63];
  assign t[139] = ~(t[165]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = ~(t[91]);
  assign t[141] = ~(t[92]);
  assign t[142] = ~(t[104] ^ t[166]);
  assign t[143] = t[113] ^ t[165];
  assign t[144] = t[8] ? t[167] : t[218];
  assign t[145] = t[8] ? t[168] : t[219];
  assign t[146] = t[169] ^ t[170];
  assign t[147] = t[108] ^ t[115];
  assign t[148] = t[171];
  assign t[149] = t[146] ^ t[172];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[95] ? t[173] : t[220];
  assign t[151] = t[174] & t[175];
  assign t[152] = t[8] ? t[176] : t[221];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[177] | t[119]);
  assign t[155] = ~(t[222]);
  assign t[156] = ~(t[213]);
  assign t[157] = ~(t[50]);
  assign t[158] = t[214] ^ t[178];
  assign t[159] = t[215] ^ t[179];
  assign t[15] = ~(t[27]);
  assign t[160] = t[28] ? x[93] : x[92];
  assign t[161] = t[28] ? x[95] : x[94];
  assign t[162] = t[216] ^ t[180];
  assign t[163] = ~(t[50]);
  assign t[164] = t[217] ^ t[181];
  assign t[165] = t[127] ^ t[92];
  assign t[166] = t[68] ^ t[91];
  assign t[167] = t[218] ^ t[182];
  assign t[168] = t[219] ^ t[183];
  assign t[169] = t[184] & t[185];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[186] & t[148];
  assign t[171] = t[8] ? t[187] : t[223];
  assign t[172] = t[188] & t[189];
  assign t[173] = t[220] ^ t[190];
  assign t[174] = ~(t[191] ^ t[35]);
  assign t[175] = t[19] ^ t[87];
  assign t[176] = t[221] ^ t[192];
  assign t[177] = ~(t[203]);
  assign t[178] = t[157] ? x[100] : x[99];
  assign t[179] = t[157] ? x[102] : x[101];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[28] ? x[104] : x[103];
  assign t[181] = t[163] ? x[106] : x[105];
  assign t[182] = t[80] ? x[108] : x[107];
  assign t[183] = t[157] ? x[110] : x[109];
  assign t[184] = ~(t[193]);
  assign t[185] = ~(t[107]);
  assign t[186] = ~(t[108]);
  assign t[187] = t[223] ^ t[194];
  assign t[188] = ~(t[169] ^ t[195]);
  assign t[189] = t[196] ^ t[193];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[163] ? x[112] : x[111];
  assign t[191] = t[123] ^ t[33];
  assign t[192] = t[80] ? x[114] : x[113];
  assign t[193] = t[148] ^ t[108];
  assign t[194] = t[80] ? x[116] : x[115];
  assign t[195] = t[147] ^ t[107];
  assign t[196] = t[107] ^ t[115];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = t[39] ^ t[40];
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[36];
  assign t[235] = t[262] ^ x[39];
  assign t[236] = t[263] ^ x[42];
  assign t[237] = t[264] ^ x[45];
  assign t[238] = t[265] ^ x[48];
  assign t[239] = t[266] ^ x[51];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[56];
  assign t[241] = t[268] ^ x[63];
  assign t[242] = t[269] ^ x[66];
  assign t[243] = t[270] ^ x[69];
  assign t[244] = t[271] ^ x[76];
  assign t[245] = t[272] ^ x[79];
  assign t[246] = t[273] ^ x[82];
  assign t[247] = t[274] ^ x[85];
  assign t[248] = t[275] ^ x[88];
  assign t[249] = t[276] ^ x[91];
  assign t[24] = t[43] ^ t[44];
  assign t[250] = t[277] ^ x[98];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = ~(t[45] ^ t[11]);
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[36];
  assign t[299] = t[353] ^ x[35];
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[39];
  assign t[301] = t[355] ^ x[38];
  assign t[302] = t[356] ^ x[42];
  assign t[303] = t[357] ^ x[41];
  assign t[304] = t[358] ^ x[45];
  assign t[305] = t[359] ^ x[44];
  assign t[306] = t[360] ^ x[48];
  assign t[307] = t[361] ^ x[47];
  assign t[308] = t[362] ^ x[51];
  assign t[309] = t[363] ^ x[50];
  assign t[30] = ~(t[199]);
  assign t[310] = t[364] ^ x[56];
  assign t[311] = t[365] ^ x[55];
  assign t[312] = t[366] ^ x[63];
  assign t[313] = t[367] ^ x[62];
  assign t[314] = t[368] ^ x[66];
  assign t[315] = t[369] ^ x[65];
  assign t[316] = t[370] ^ x[69];
  assign t[317] = t[371] ^ x[68];
  assign t[318] = t[372] ^ x[76];
  assign t[319] = t[373] ^ x[75];
  assign t[31] = ~(t[200]);
  assign t[320] = t[374] ^ x[79];
  assign t[321] = t[375] ^ x[78];
  assign t[322] = t[376] ^ x[82];
  assign t[323] = t[377] ^ x[81];
  assign t[324] = t[378] ^ x[85];
  assign t[325] = t[379] ^ x[84];
  assign t[326] = t[380] ^ x[88];
  assign t[327] = t[381] ^ x[87];
  assign t[328] = t[382] ^ x[91];
  assign t[329] = t[383] ^ x[90];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[384] ^ x[98];
  assign t[331] = t[385] ^ x[97];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = t[200] ^ t[53];
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = t[201] ^ t[54];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[34]);
  assign t[353] = (x[34]);
  assign t[354] = (x[37]);
  assign t[355] = (x[37]);
  assign t[356] = (x[40]);
  assign t[357] = (x[40]);
  assign t[358] = (x[43]);
  assign t[359] = (x[43]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[46]);
  assign t[361] = (x[46]);
  assign t[362] = (x[49]);
  assign t[363] = (x[49]);
  assign t[364] = (x[54]);
  assign t[365] = (x[54]);
  assign t[366] = (x[61]);
  assign t[367] = (x[61]);
  assign t[368] = (x[64]);
  assign t[369] = (x[64]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[67]);
  assign t[371] = (x[67]);
  assign t[372] = (x[74]);
  assign t[373] = (x[74]);
  assign t[374] = (x[77]);
  assign t[375] = (x[77]);
  assign t[376] = (x[80]);
  assign t[377] = (x[80]);
  assign t[378] = (x[83]);
  assign t[379] = (x[83]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[86]);
  assign t[381] = (x[86]);
  assign t[382] = (x[89]);
  assign t[383] = (x[89]);
  assign t[384] = (x[96]);
  assign t[385] = (x[96]);
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[8] ? t[66] : t[202];
  assign t[42] = t[67] ^ t[60];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = ~(t[72] ^ t[73]);
  assign t[46] = t[22] ^ t[74];
  assign t[47] = ~(t[75] ^ t[76]);
  assign t[48] = ~(t[77] & t[78]);
  assign t[49] = t[203] | t[79];
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[80]);
  assign t[51] = ~(t[201]);
  assign t[52] = ~(t[81] & t[204]);
  assign t[53] = t[8] ? t[82] : t[205];
  assign t[54] = t[8] ? t[83] : t[206];
  assign t[55] = t[84] & t[85];
  assign t[56] = t[86] & t[87];
  assign t[57] = ~(t[55] ^ t[88]);
  assign t[58] = t[89] ^ t[90];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] & t[94];
  assign t[61] = t[95] ? t[96] : t[207];
  assign t[62] = t[64] ^ t[97];
  assign t[63] = t[95] ? t[98] : t[208];
  assign t[64] = t[99] ^ t[100];
  assign t[65] = t[101] & t[102];
  assign t[66] = t[202] ^ t[103];
  assign t[67] = t[104] ^ t[105];
  assign t[68] = t[92] ^ t[41];
  assign t[69] = t[67] ^ t[106];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[107] ^ t[108];
  assign t[71] = t[109] & t[110];
  assign t[72] = t[111] ^ t[23];
  assign t[73] = t[112] ^ t[97];
  assign t[74] = t[113] ^ t[105];
  assign t[75] = t[34] ^ t[114];
  assign t[76] = t[115] ^ t[116];
  assign t[77] = ~(t[79] & t[117]);
  assign t[78] = ~(t[209] ^ t[118]);
  assign t[79] = ~(t[119] & t[120]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[49]);
  assign t[81] = ~(t[210]);
  assign t[82] = t[205] ^ t[121];
  assign t[83] = t[206] ^ t[122];
  assign t[84] = ~(t[90]);
  assign t[85] = ~(t[123]);
  assign t[86] = ~(t[33]);
  assign t[87] = t[210] ^ t[124];
  assign t[88] = t[19] ^ t[123];
  assign t[89] = t[123] ^ t[34];
  assign t[8] = ~(t[15]);
  assign t[90] = t[87] ^ t[33];
  assign t[91] = t[8] ? t[125] : t[211];
  assign t[92] = t[8] ? t[126] : t[212];
  assign t[93] = ~(t[59] ^ t[67]);
  assign t[94] = t[68] ^ t[127];
  assign t[95] = ~(t[15]);
  assign t[96] = t[207] ^ t[128];
  assign t[97] = t[129] & t[130];
  assign t[98] = t[208] ^ t[131];
  assign t[99] = t[132] & t[133];
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[134] & t[135];
  assign t[101] = ~(t[99] ^ t[136]);
  assign t[102] = t[137] ^ t[138];
  assign t[103] = t[80] ? x[53] : x[52];
  assign t[104] = t[139] & t[140];
  assign t[105] = t[141] & t[127];
  assign t[106] = t[142] & t[143];
  assign t[107] = t[144];
  assign t[108] = ~t[145];
  assign t[109] = ~(t[70] ^ t[146]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[147] ^ t[148];
  assign t[111] = t[147] ^ t[149];
  assign t[112] = t[150] ^ t[63];
  assign t[113] = t[91] ^ t[41];
  assign t[114] = t[35] ^ t[151];
  assign t[115] = t[152];
  assign t[116] = t[146] ^ t[71];
  assign t[117] = ~(t[153] & t[154]);
  assign t[118] = t[155] ^ t[213];
  assign t[119] = ~(t[209]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[156] & t[155];
  assign t[121] = t[157] ? x[58] : x[57];
  assign t[122] = t[157] ? x[60] : x[59];
  assign t[123] = t[8] ? t[158] : t[214];
  assign t[124] = t[8] ? t[159] : t[215];
  assign t[125] = t[211] ^ t[160];
  assign t[126] = t[212] ^ t[161];
  assign t[127] = t[8] ? t[162] : t[216];
  assign t[128] = t[163] ? x[71] : x[70];
  assign t[129] = ~(t[112] ^ t[64]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[39] ^ t[135];
  assign t[131] = t[163] ? x[73] : x[72];
  assign t[132] = ~(t[138]);
  assign t[133] = ~(t[150]);
  assign t[134] = ~(t[63]);
  assign t[135] = t[95] ? t[164] : t[217];
  assign t[136] = t[39] ^ t[150];
  assign t[137] = t[150] ^ t[61];
  assign t[138] = t[135] ^ t[63];
  assign t[139] = ~(t[165]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = ~(t[91]);
  assign t[141] = ~(t[92]);
  assign t[142] = ~(t[104] ^ t[166]);
  assign t[143] = t[113] ^ t[165];
  assign t[144] = t[8] ? t[167] : t[218];
  assign t[145] = t[8] ? t[168] : t[219];
  assign t[146] = t[169] ^ t[170];
  assign t[147] = t[108] ^ t[115];
  assign t[148] = t[171];
  assign t[149] = t[146] ^ t[172];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[95] ? t[173] : t[220];
  assign t[151] = t[174] & t[175];
  assign t[152] = t[8] ? t[176] : t[221];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[177] | t[119]);
  assign t[155] = ~(t[222]);
  assign t[156] = ~(t[213]);
  assign t[157] = ~(t[50]);
  assign t[158] = t[214] ^ t[178];
  assign t[159] = t[215] ^ t[179];
  assign t[15] = ~(t[27]);
  assign t[160] = t[28] ? x[93] : x[92];
  assign t[161] = t[28] ? x[95] : x[94];
  assign t[162] = t[216] ^ t[180];
  assign t[163] = ~(t[50]);
  assign t[164] = t[217] ^ t[181];
  assign t[165] = t[127] ^ t[92];
  assign t[166] = t[68] ^ t[91];
  assign t[167] = t[218] ^ t[182];
  assign t[168] = t[219] ^ t[183];
  assign t[169] = t[184] & t[185];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[186] & t[148];
  assign t[171] = t[8] ? t[187] : t[223];
  assign t[172] = t[188] & t[189];
  assign t[173] = t[220] ^ t[190];
  assign t[174] = ~(t[191] ^ t[35]);
  assign t[175] = t[19] ^ t[87];
  assign t[176] = t[221] ^ t[192];
  assign t[177] = ~(t[203]);
  assign t[178] = t[157] ? x[100] : x[99];
  assign t[179] = t[157] ? x[102] : x[101];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[28] ? x[104] : x[103];
  assign t[181] = t[163] ? x[106] : x[105];
  assign t[182] = t[80] ? x[108] : x[107];
  assign t[183] = t[157] ? x[110] : x[109];
  assign t[184] = ~(t[193]);
  assign t[185] = ~(t[107]);
  assign t[186] = ~(t[108]);
  assign t[187] = t[223] ^ t[194];
  assign t[188] = ~(t[169] ^ t[195]);
  assign t[189] = t[196] ^ t[193];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[163] ? x[112] : x[111];
  assign t[191] = t[123] ^ t[33];
  assign t[192] = t[80] ? x[114] : x[113];
  assign t[193] = t[148] ^ t[108];
  assign t[194] = t[80] ? x[116] : x[115];
  assign t[195] = t[147] ^ t[107];
  assign t[196] = t[107] ^ t[115];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = t[39] ^ t[40];
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[36];
  assign t[235] = t[262] ^ x[39];
  assign t[236] = t[263] ^ x[42];
  assign t[237] = t[264] ^ x[45];
  assign t[238] = t[265] ^ x[48];
  assign t[239] = t[266] ^ x[51];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[56];
  assign t[241] = t[268] ^ x[63];
  assign t[242] = t[269] ^ x[66];
  assign t[243] = t[270] ^ x[69];
  assign t[244] = t[271] ^ x[76];
  assign t[245] = t[272] ^ x[79];
  assign t[246] = t[273] ^ x[82];
  assign t[247] = t[274] ^ x[85];
  assign t[248] = t[275] ^ x[88];
  assign t[249] = t[276] ^ x[91];
  assign t[24] = t[43] ^ t[44];
  assign t[250] = t[277] ^ x[98];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = ~(t[45] ^ t[11]);
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[36];
  assign t[299] = t[353] ^ x[35];
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[39];
  assign t[301] = t[355] ^ x[38];
  assign t[302] = t[356] ^ x[42];
  assign t[303] = t[357] ^ x[41];
  assign t[304] = t[358] ^ x[45];
  assign t[305] = t[359] ^ x[44];
  assign t[306] = t[360] ^ x[48];
  assign t[307] = t[361] ^ x[47];
  assign t[308] = t[362] ^ x[51];
  assign t[309] = t[363] ^ x[50];
  assign t[30] = ~(t[199]);
  assign t[310] = t[364] ^ x[56];
  assign t[311] = t[365] ^ x[55];
  assign t[312] = t[366] ^ x[63];
  assign t[313] = t[367] ^ x[62];
  assign t[314] = t[368] ^ x[66];
  assign t[315] = t[369] ^ x[65];
  assign t[316] = t[370] ^ x[69];
  assign t[317] = t[371] ^ x[68];
  assign t[318] = t[372] ^ x[76];
  assign t[319] = t[373] ^ x[75];
  assign t[31] = ~(t[200]);
  assign t[320] = t[374] ^ x[79];
  assign t[321] = t[375] ^ x[78];
  assign t[322] = t[376] ^ x[82];
  assign t[323] = t[377] ^ x[81];
  assign t[324] = t[378] ^ x[85];
  assign t[325] = t[379] ^ x[84];
  assign t[326] = t[380] ^ x[88];
  assign t[327] = t[381] ^ x[87];
  assign t[328] = t[382] ^ x[91];
  assign t[329] = t[383] ^ x[90];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[384] ^ x[98];
  assign t[331] = t[385] ^ x[97];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = t[200] ^ t[53];
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = t[201] ^ t[54];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[34]);
  assign t[353] = (x[34]);
  assign t[354] = (x[37]);
  assign t[355] = (x[37]);
  assign t[356] = (x[40]);
  assign t[357] = (x[40]);
  assign t[358] = (x[43]);
  assign t[359] = (x[43]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[46]);
  assign t[361] = (x[46]);
  assign t[362] = (x[49]);
  assign t[363] = (x[49]);
  assign t[364] = (x[54]);
  assign t[365] = (x[54]);
  assign t[366] = (x[61]);
  assign t[367] = (x[61]);
  assign t[368] = (x[64]);
  assign t[369] = (x[64]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[67]);
  assign t[371] = (x[67]);
  assign t[372] = (x[74]);
  assign t[373] = (x[74]);
  assign t[374] = (x[77]);
  assign t[375] = (x[77]);
  assign t[376] = (x[80]);
  assign t[377] = (x[80]);
  assign t[378] = (x[83]);
  assign t[379] = (x[83]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[86]);
  assign t[381] = (x[86]);
  assign t[382] = (x[89]);
  assign t[383] = (x[89]);
  assign t[384] = (x[96]);
  assign t[385] = (x[96]);
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = t[8] ? t[66] : t[202];
  assign t[42] = t[67] ^ t[60];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = ~(t[72] ^ t[73]);
  assign t[46] = t[22] ^ t[74];
  assign t[47] = ~(t[75] ^ t[76]);
  assign t[48] = ~(t[77] & t[78]);
  assign t[49] = t[203] | t[79];
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[80]);
  assign t[51] = ~(t[201]);
  assign t[52] = ~(t[81] & t[204]);
  assign t[53] = t[8] ? t[82] : t[205];
  assign t[54] = t[8] ? t[83] : t[206];
  assign t[55] = t[84] & t[85];
  assign t[56] = t[86] & t[87];
  assign t[57] = ~(t[55] ^ t[88]);
  assign t[58] = t[89] ^ t[90];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] & t[94];
  assign t[61] = t[95] ? t[96] : t[207];
  assign t[62] = t[64] ^ t[97];
  assign t[63] = t[95] ? t[98] : t[208];
  assign t[64] = t[99] ^ t[100];
  assign t[65] = t[101] & t[102];
  assign t[66] = t[202] ^ t[103];
  assign t[67] = t[104] ^ t[105];
  assign t[68] = t[92] ^ t[41];
  assign t[69] = t[67] ^ t[106];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[107] ^ t[108];
  assign t[71] = t[109] & t[110];
  assign t[72] = t[111] ^ t[23];
  assign t[73] = t[112] ^ t[97];
  assign t[74] = t[113] ^ t[105];
  assign t[75] = t[34] ^ t[114];
  assign t[76] = t[115] ^ t[116];
  assign t[77] = ~(t[79] & t[117]);
  assign t[78] = ~(t[209] ^ t[118]);
  assign t[79] = ~(t[119] & t[120]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[49]);
  assign t[81] = ~(t[210]);
  assign t[82] = t[205] ^ t[121];
  assign t[83] = t[206] ^ t[122];
  assign t[84] = ~(t[90]);
  assign t[85] = ~(t[123]);
  assign t[86] = ~(t[33]);
  assign t[87] = t[210] ^ t[124];
  assign t[88] = t[19] ^ t[123];
  assign t[89] = t[123] ^ t[34];
  assign t[8] = ~(t[15]);
  assign t[90] = t[87] ^ t[33];
  assign t[91] = t[8] ? t[125] : t[211];
  assign t[92] = t[8] ? t[126] : t[212];
  assign t[93] = ~(t[59] ^ t[67]);
  assign t[94] = t[68] ^ t[127];
  assign t[95] = ~(t[15]);
  assign t[96] = t[207] ^ t[128];
  assign t[97] = t[129] & t[130];
  assign t[98] = t[208] ^ t[131];
  assign t[99] = t[132] & t[133];
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [116:0] x;
 output y;

 wire [383:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[87]);
  assign t[101] = ~(t[88]);
  assign t[102] = t[201] ^ t[138];
  assign t[103] = t[88] ^ t[27];
  assign t[104] = t[205] ^ t[139];
  assign t[105] = t[206] ^ t[140];
  assign t[106] = t[141] & t[142];
  assign t[107] = t[143] & t[72];
  assign t[108] = t[144];
  assign t[109] = t[9] ? t[145] : t[214];
  assign t[10] = t[195] ^ t[20];
  assign t[110] = ~(t[146] & t[147]);
  assign t[111] = t[148] ^ t[215];
  assign t[112] = ~(t[207]);
  assign t[113] = t[149] & t[148];
  assign t[114] = t[150] ^ t[65];
  assign t[115] = ~(t[151] ^ t[40]);
  assign t[116] = t[152] ^ t[153];
  assign t[117] = t[44] ^ t[108];
  assign t[118] = t[70] ^ t[30];
  assign t[119] = t[208] ^ t[154];
  assign t[11] = ~(t[196]);
  assign t[120] = t[209] ^ t[155];
  assign t[121] = t[9] ? t[156] : t[216];
  assign t[122] = t[210] ^ t[157];
  assign t[123] = t[158] & t[159];
  assign t[124] = t[160] ^ t[54];
  assign t[125] = t[161] & t[162];
  assign t[126] = t[211] ^ t[163];
  assign t[127] = t[9] ? t[164] : t[217];
  assign t[128] = t[212] ^ t[165];
  assign t[129] = t[94] ? t[166] : t[218];
  assign t[12] = ~(t[197]);
  assign t[130] = t[213] ^ t[167];
  assign t[131] = t[168] & t[169];
  assign t[132] = t[170] ? x[79] : x[78];
  assign t[133] = t[171] & t[172];
  assign t[134] = ~(t[173] ^ t[96]);
  assign t[135] = t[152] ^ t[91];
  assign t[136] = ~(t[50]);
  assign t[137] = t[102] ^ t[88];
  assign t[138] = t[9] ? t[174] : t[219];
  assign t[139] = t[76] ? x[84] : x[83];
  assign t[13] = ~(t[198]);
  assign t[140] = t[136] ? x[86] : x[85];
  assign t[141] = ~(t[175]);
  assign t[142] = ~(t[44]);
  assign t[143] = ~(t[45]);
  assign t[144] = t[9] ? t[176] : t[220];
  assign t[145] = t[214] ^ t[177];
  assign t[146] = ~(t[149] | t[148]);
  assign t[147] = ~(t[178] | t[112]);
  assign t[148] = ~(t[221]);
  assign t[149] = ~(t[215]);
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = t[87] ^ t[27];
  assign t[151] = t[179] ^ t[125];
  assign t[152] = t[129] ^ t[61];
  assign t[153] = t[96] ^ t[180];
  assign t[154] = t[32] ? x[94] : x[93];
  assign t[155] = t[76] ? x[96] : x[95];
  assign t[156] = t[216] ^ t[181];
  assign t[157] = t[32] ? x[98] : x[97];
  assign t[158] = ~(t[106] ^ t[182]);
  assign t[159] = t[117] ^ t[175];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[183] & t[184];
  assign t[161] = ~(t[179] ^ t[124]);
  assign t[162] = t[92] ^ t[84];
  assign t[163] = t[136] ? x[100] : x[99];
  assign t[164] = t[217] ^ t[185];
  assign t[165] = t[170] ? x[102] : x[101];
  assign t[166] = t[218] ^ t[186];
  assign t[167] = t[170] ? x[104] : x[103];
  assign t[168] = ~(t[160] ^ t[187]);
  assign t[169] = t[53] ^ t[188];
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = ~(t[50]);
  assign t[171] = ~(t[189]);
  assign t[172] = ~(t[89]);
  assign t[173] = t[89] ^ t[129];
  assign t[174] = t[219] ^ t[190];
  assign t[175] = t[72] ^ t[45];
  assign t[176] = t[220] ^ t[191];
  assign t[177] = t[76] ? x[106] : x[105];
  assign t[178] = ~(t[203]);
  assign t[179] = t[81] ^ t[121];
  assign t[17] = t[27] ^ t[28];
  assign t[180] = t[192] & t[193];
  assign t[181] = t[32] ? x[108] : x[107];
  assign t[182] = t[71] ^ t[44];
  assign t[183] = ~(t[188]);
  assign t[184] = ~(t[81]);
  assign t[185] = t[136] ? x[110] : x[109];
  assign t[186] = t[170] ? x[112] : x[111];
  assign t[187] = t[92] ^ t[81];
  assign t[188] = t[84] ^ t[121];
  assign t[189] = t[91] ^ t[129];
  assign t[18] = t[29] ^ t[30];
  assign t[190] = t[136] ? x[114] : x[113];
  assign t[191] = t[76] ? x[116] : x[115];
  assign t[192] = ~(t[133] ^ t[194]);
  assign t[193] = t[58] ^ t[189];
  assign t[194] = t[152] ^ t[89];
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[199]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = t[249] ^ x[4];
  assign t[223] = t[250] ^ x[7];
  assign t[224] = t[251] ^ x[10];
  assign t[225] = t[252] ^ x[13];
  assign t[226] = t[253] ^ x[18];
  assign t[227] = t[254] ^ x[21];
  assign t[228] = t[255] ^ x[24];
  assign t[229] = t[256] ^ x[27];
  assign t[22] = ~(t[33] & t[200]);
  assign t[230] = t[257] ^ x[30];
  assign t[231] = t[258] ^ x[33];
  assign t[232] = t[259] ^ x[36];
  assign t[233] = t[260] ^ x[39];
  assign t[234] = t[261] ^ x[42];
  assign t[235] = t[262] ^ x[45];
  assign t[236] = t[263] ^ x[48];
  assign t[237] = t[264] ^ x[51];
  assign t[238] = t[265] ^ x[54];
  assign t[239] = t[266] ^ x[57];
  assign t[23] = t[34] ^ t[35];
  assign t[240] = t[267] ^ x[60];
  assign t[241] = t[268] ^ x[65];
  assign t[242] = t[269] ^ x[68];
  assign t[243] = t[270] ^ x[71];
  assign t[244] = t[271] ^ x[74];
  assign t[245] = t[272] ^ x[77];
  assign t[246] = t[273] ^ x[82];
  assign t[247] = t[274] ^ x[89];
  assign t[248] = t[275] ^ x[92];
  assign t[249] = (t[276] & ~t[277]);
  assign t[24] = ~(t[36] ^ t[37]);
  assign t[250] = (t[278] & ~t[279]);
  assign t[251] = (t[280] & ~t[281]);
  assign t[252] = (t[282] & ~t[283]);
  assign t[253] = (t[284] & ~t[285]);
  assign t[254] = (t[286] & ~t[287]);
  assign t[255] = (t[288] & ~t[289]);
  assign t[256] = (t[290] & ~t[291]);
  assign t[257] = (t[292] & ~t[293]);
  assign t[258] = (t[294] & ~t[295]);
  assign t[259] = (t[296] & ~t[297]);
  assign t[25] = t[38] ^ t[37];
  assign t[260] = (t[298] & ~t[299]);
  assign t[261] = (t[300] & ~t[301]);
  assign t[262] = (t[302] & ~t[303]);
  assign t[263] = (t[304] & ~t[305]);
  assign t[264] = (t[306] & ~t[307]);
  assign t[265] = (t[308] & ~t[309]);
  assign t[266] = (t[310] & ~t[311]);
  assign t[267] = (t[312] & ~t[313]);
  assign t[268] = (t[314] & ~t[315]);
  assign t[269] = (t[316] & ~t[317]);
  assign t[26] = ~(t[39] ^ t[40]);
  assign t[270] = (t[318] & ~t[319]);
  assign t[271] = (t[320] & ~t[321]);
  assign t[272] = (t[322] & ~t[323]);
  assign t[273] = (t[324] & ~t[325]);
  assign t[274] = (t[326] & ~t[327]);
  assign t[275] = (t[328] & ~t[329]);
  assign t[276] = t[330] ^ x[4];
  assign t[277] = t[331] ^ x[3];
  assign t[278] = t[332] ^ x[7];
  assign t[279] = t[333] ^ x[6];
  assign t[27] = t[199] ^ t[41];
  assign t[280] = t[334] ^ x[10];
  assign t[281] = t[335] ^ x[9];
  assign t[282] = t[336] ^ x[13];
  assign t[283] = t[337] ^ x[12];
  assign t[284] = t[338] ^ x[18];
  assign t[285] = t[339] ^ x[17];
  assign t[286] = t[340] ^ x[21];
  assign t[287] = t[341] ^ x[20];
  assign t[288] = t[342] ^ x[24];
  assign t[289] = t[343] ^ x[23];
  assign t[28] = t[42] ^ t[43];
  assign t[290] = t[344] ^ x[27];
  assign t[291] = t[345] ^ x[26];
  assign t[292] = t[346] ^ x[30];
  assign t[293] = t[347] ^ x[29];
  assign t[294] = t[348] ^ x[33];
  assign t[295] = t[349] ^ x[32];
  assign t[296] = t[350] ^ x[36];
  assign t[297] = t[351] ^ x[35];
  assign t[298] = t[352] ^ x[39];
  assign t[299] = t[353] ^ x[38];
  assign t[29] = t[44] ^ t[45];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[42];
  assign t[301] = t[355] ^ x[41];
  assign t[302] = t[356] ^ x[45];
  assign t[303] = t[357] ^ x[44];
  assign t[304] = t[358] ^ x[48];
  assign t[305] = t[359] ^ x[47];
  assign t[306] = t[360] ^ x[51];
  assign t[307] = t[361] ^ x[50];
  assign t[308] = t[362] ^ x[54];
  assign t[309] = t[363] ^ x[53];
  assign t[30] = t[46] & t[47];
  assign t[310] = t[364] ^ x[57];
  assign t[311] = t[365] ^ x[56];
  assign t[312] = t[366] ^ x[60];
  assign t[313] = t[367] ^ x[59];
  assign t[314] = t[368] ^ x[65];
  assign t[315] = t[369] ^ x[64];
  assign t[316] = t[370] ^ x[68];
  assign t[317] = t[371] ^ x[67];
  assign t[318] = t[372] ^ x[71];
  assign t[319] = t[373] ^ x[70];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[74];
  assign t[321] = t[375] ^ x[73];
  assign t[322] = t[376] ^ x[77];
  assign t[323] = t[377] ^ x[76];
  assign t[324] = t[378] ^ x[82];
  assign t[325] = t[379] ^ x[81];
  assign t[326] = t[380] ^ x[89];
  assign t[327] = t[381] ^ x[88];
  assign t[328] = t[382] ^ x[92];
  assign t[329] = t[383] ^ x[91];
  assign t[32] = ~(t[50]);
  assign t[330] = (x[2]);
  assign t[331] = (x[2]);
  assign t[332] = (x[5]);
  assign t[333] = (x[5]);
  assign t[334] = (x[8]);
  assign t[335] = (x[8]);
  assign t[336] = (x[11]);
  assign t[337] = (x[11]);
  assign t[338] = (x[16]);
  assign t[339] = (x[16]);
  assign t[33] = ~(t[201]);
  assign t[340] = (x[19]);
  assign t[341] = (x[19]);
  assign t[342] = (x[22]);
  assign t[343] = (x[22]);
  assign t[344] = (x[25]);
  assign t[345] = (x[25]);
  assign t[346] = (x[28]);
  assign t[347] = (x[28]);
  assign t[348] = (x[31]);
  assign t[349] = (x[31]);
  assign t[34] = ~(t[51] ^ t[52]);
  assign t[350] = (x[34]);
  assign t[351] = (x[34]);
  assign t[352] = (x[37]);
  assign t[353] = (x[37]);
  assign t[354] = (x[40]);
  assign t[355] = (x[40]);
  assign t[356] = (x[43]);
  assign t[357] = (x[43]);
  assign t[358] = (x[46]);
  assign t[359] = (x[46]);
  assign t[35] = t[53] ^ t[54];
  assign t[360] = (x[49]);
  assign t[361] = (x[49]);
  assign t[362] = (x[52]);
  assign t[363] = (x[52]);
  assign t[364] = (x[55]);
  assign t[365] = (x[55]);
  assign t[366] = (x[58]);
  assign t[367] = (x[58]);
  assign t[368] = (x[63]);
  assign t[369] = (x[63]);
  assign t[36] = t[55] ^ t[56];
  assign t[370] = (x[66]);
  assign t[371] = (x[66]);
  assign t[372] = (x[69]);
  assign t[373] = (x[69]);
  assign t[374] = (x[72]);
  assign t[375] = (x[72]);
  assign t[376] = (x[75]);
  assign t[377] = (x[75]);
  assign t[378] = (x[80]);
  assign t[379] = (x[80]);
  assign t[37] = t[57] ^ t[43];
  assign t[380] = (x[87]);
  assign t[381] = (x[87]);
  assign t[382] = (x[90]);
  assign t[383] = (x[90]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[60] ^ t[18];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[9] ? t[63] : t[202];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[68];
  assign t[45] = ~t[69];
  assign t[46] = ~(t[29] ^ t[70]);
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[203] | t[75];
  assign t[4] = t[9] ? t[10] : t[195];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[71] ^ t[85];
  assign t[56] = t[82] ^ t[86];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] ^ t[61];
  assign t[59] = t[90] & t[91];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[94] ? t[95] : t[204];
  assign t[62] = t[96] ^ t[97];
  assign t[63] = t[202] ^ t[98];
  assign t[64] = t[99] & t[100];
  assign t[65] = t[101] & t[102];
  assign t[66] = ~(t[57] ^ t[42]);
  assign t[67] = t[103] ^ t[102];
  assign t[68] = t[9] ? t[104] : t[205];
  assign t[69] = t[9] ? t[105] : t[206];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[106] ^ t[107];
  assign t[71] = t[45] ^ t[108];
  assign t[72] = t[109];
  assign t[73] = ~(t[75] & t[110]);
  assign t[74] = ~(t[207] ^ t[111]);
  assign t[75] = ~(t[112] & t[113]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[17] ^ t[114];
  assign t[78] = ~(t[115] ^ t[116]);
  assign t[79] = t[117] ^ t[107];
  assign t[7] = t[15] ^ t[16];
  assign t[80] = t[108] ^ t[118];
  assign t[81] = t[9] ? t[119] : t[208];
  assign t[82] = t[9] ? t[120] : t[209];
  assign t[83] = ~(t[121]);
  assign t[84] = t[9] ? t[122] : t[210];
  assign t[85] = t[70] ^ t[123];
  assign t[86] = t[124] ^ t[125];
  assign t[87] = t[9] ? t[126] : t[211];
  assign t[88] = t[198] ^ t[127];
  assign t[89] = t[94] ? t[128] : t[212];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = ~(t[129]);
  assign t[91] = t[94] ? t[130] : t[213];
  assign t[92] = t[121] ^ t[82];
  assign t[93] = t[124] ^ t[131];
  assign t[94] = ~(t[19]);
  assign t[95] = t[204] ^ t[132];
  assign t[96] = t[133] ^ t[59];
  assign t[97] = t[134] & t[135];
  assign t[98] = t[136] ? x[62] : x[61];
  assign t[99] = ~(t[137]);
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind111(x, y);
 input [116:0] x;
 output y;

 wire [383:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[87]);
  assign t[101] = ~(t[88]);
  assign t[102] = t[201] ^ t[138];
  assign t[103] = t[88] ^ t[27];
  assign t[104] = t[205] ^ t[139];
  assign t[105] = t[206] ^ t[140];
  assign t[106] = t[141] & t[142];
  assign t[107] = t[143] & t[72];
  assign t[108] = t[144];
  assign t[109] = t[9] ? t[145] : t[214];
  assign t[10] = t[195] ^ t[20];
  assign t[110] = ~(t[146] & t[147]);
  assign t[111] = t[148] ^ t[215];
  assign t[112] = ~(t[207]);
  assign t[113] = t[149] & t[148];
  assign t[114] = t[150] ^ t[65];
  assign t[115] = ~(t[151] ^ t[40]);
  assign t[116] = t[152] ^ t[153];
  assign t[117] = t[44] ^ t[108];
  assign t[118] = t[70] ^ t[30];
  assign t[119] = t[208] ^ t[154];
  assign t[11] = ~(t[196]);
  assign t[120] = t[209] ^ t[155];
  assign t[121] = t[9] ? t[156] : t[216];
  assign t[122] = t[210] ^ t[157];
  assign t[123] = t[158] & t[159];
  assign t[124] = t[160] ^ t[54];
  assign t[125] = t[161] & t[162];
  assign t[126] = t[211] ^ t[163];
  assign t[127] = t[9] ? t[164] : t[217];
  assign t[128] = t[212] ^ t[165];
  assign t[129] = t[94] ? t[166] : t[218];
  assign t[12] = ~(t[197]);
  assign t[130] = t[213] ^ t[167];
  assign t[131] = t[168] & t[169];
  assign t[132] = t[170] ? x[79] : x[78];
  assign t[133] = t[171] & t[172];
  assign t[134] = ~(t[173] ^ t[96]);
  assign t[135] = t[152] ^ t[91];
  assign t[136] = ~(t[50]);
  assign t[137] = t[102] ^ t[88];
  assign t[138] = t[9] ? t[174] : t[219];
  assign t[139] = t[76] ? x[84] : x[83];
  assign t[13] = ~(t[198]);
  assign t[140] = t[136] ? x[86] : x[85];
  assign t[141] = ~(t[175]);
  assign t[142] = ~(t[44]);
  assign t[143] = ~(t[45]);
  assign t[144] = t[9] ? t[176] : t[220];
  assign t[145] = t[214] ^ t[177];
  assign t[146] = ~(t[149] | t[148]);
  assign t[147] = ~(t[178] | t[112]);
  assign t[148] = ~(t[221]);
  assign t[149] = ~(t[215]);
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = t[87] ^ t[27];
  assign t[151] = t[179] ^ t[125];
  assign t[152] = t[129] ^ t[61];
  assign t[153] = t[96] ^ t[180];
  assign t[154] = t[32] ? x[94] : x[93];
  assign t[155] = t[76] ? x[96] : x[95];
  assign t[156] = t[216] ^ t[181];
  assign t[157] = t[32] ? x[98] : x[97];
  assign t[158] = ~(t[106] ^ t[182]);
  assign t[159] = t[117] ^ t[175];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[183] & t[184];
  assign t[161] = ~(t[179] ^ t[124]);
  assign t[162] = t[92] ^ t[84];
  assign t[163] = t[136] ? x[100] : x[99];
  assign t[164] = t[217] ^ t[185];
  assign t[165] = t[170] ? x[102] : x[101];
  assign t[166] = t[218] ^ t[186];
  assign t[167] = t[170] ? x[104] : x[103];
  assign t[168] = ~(t[160] ^ t[187]);
  assign t[169] = t[53] ^ t[188];
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = ~(t[50]);
  assign t[171] = ~(t[189]);
  assign t[172] = ~(t[89]);
  assign t[173] = t[89] ^ t[129];
  assign t[174] = t[219] ^ t[190];
  assign t[175] = t[72] ^ t[45];
  assign t[176] = t[220] ^ t[191];
  assign t[177] = t[76] ? x[106] : x[105];
  assign t[178] = ~(t[203]);
  assign t[179] = t[81] ^ t[121];
  assign t[17] = t[27] ^ t[28];
  assign t[180] = t[192] & t[193];
  assign t[181] = t[32] ? x[108] : x[107];
  assign t[182] = t[71] ^ t[44];
  assign t[183] = ~(t[188]);
  assign t[184] = ~(t[81]);
  assign t[185] = t[136] ? x[110] : x[109];
  assign t[186] = t[170] ? x[112] : x[111];
  assign t[187] = t[92] ^ t[81];
  assign t[188] = t[84] ^ t[121];
  assign t[189] = t[91] ^ t[129];
  assign t[18] = t[29] ^ t[30];
  assign t[190] = t[136] ? x[114] : x[113];
  assign t[191] = t[76] ? x[116] : x[115];
  assign t[192] = ~(t[133] ^ t[194]);
  assign t[193] = t[58] ^ t[189];
  assign t[194] = t[152] ^ t[89];
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[199]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = t[249] ^ x[4];
  assign t[223] = t[250] ^ x[7];
  assign t[224] = t[251] ^ x[10];
  assign t[225] = t[252] ^ x[13];
  assign t[226] = t[253] ^ x[18];
  assign t[227] = t[254] ^ x[21];
  assign t[228] = t[255] ^ x[24];
  assign t[229] = t[256] ^ x[27];
  assign t[22] = ~(t[33] & t[200]);
  assign t[230] = t[257] ^ x[30];
  assign t[231] = t[258] ^ x[33];
  assign t[232] = t[259] ^ x[36];
  assign t[233] = t[260] ^ x[39];
  assign t[234] = t[261] ^ x[42];
  assign t[235] = t[262] ^ x[45];
  assign t[236] = t[263] ^ x[48];
  assign t[237] = t[264] ^ x[51];
  assign t[238] = t[265] ^ x[54];
  assign t[239] = t[266] ^ x[57];
  assign t[23] = t[34] ^ t[35];
  assign t[240] = t[267] ^ x[60];
  assign t[241] = t[268] ^ x[65];
  assign t[242] = t[269] ^ x[68];
  assign t[243] = t[270] ^ x[71];
  assign t[244] = t[271] ^ x[74];
  assign t[245] = t[272] ^ x[77];
  assign t[246] = t[273] ^ x[82];
  assign t[247] = t[274] ^ x[89];
  assign t[248] = t[275] ^ x[92];
  assign t[249] = (t[276] & ~t[277]);
  assign t[24] = ~(t[36] ^ t[37]);
  assign t[250] = (t[278] & ~t[279]);
  assign t[251] = (t[280] & ~t[281]);
  assign t[252] = (t[282] & ~t[283]);
  assign t[253] = (t[284] & ~t[285]);
  assign t[254] = (t[286] & ~t[287]);
  assign t[255] = (t[288] & ~t[289]);
  assign t[256] = (t[290] & ~t[291]);
  assign t[257] = (t[292] & ~t[293]);
  assign t[258] = (t[294] & ~t[295]);
  assign t[259] = (t[296] & ~t[297]);
  assign t[25] = t[38] ^ t[37];
  assign t[260] = (t[298] & ~t[299]);
  assign t[261] = (t[300] & ~t[301]);
  assign t[262] = (t[302] & ~t[303]);
  assign t[263] = (t[304] & ~t[305]);
  assign t[264] = (t[306] & ~t[307]);
  assign t[265] = (t[308] & ~t[309]);
  assign t[266] = (t[310] & ~t[311]);
  assign t[267] = (t[312] & ~t[313]);
  assign t[268] = (t[314] & ~t[315]);
  assign t[269] = (t[316] & ~t[317]);
  assign t[26] = ~(t[39] ^ t[40]);
  assign t[270] = (t[318] & ~t[319]);
  assign t[271] = (t[320] & ~t[321]);
  assign t[272] = (t[322] & ~t[323]);
  assign t[273] = (t[324] & ~t[325]);
  assign t[274] = (t[326] & ~t[327]);
  assign t[275] = (t[328] & ~t[329]);
  assign t[276] = t[330] ^ x[4];
  assign t[277] = t[331] ^ x[3];
  assign t[278] = t[332] ^ x[7];
  assign t[279] = t[333] ^ x[6];
  assign t[27] = t[199] ^ t[41];
  assign t[280] = t[334] ^ x[10];
  assign t[281] = t[335] ^ x[9];
  assign t[282] = t[336] ^ x[13];
  assign t[283] = t[337] ^ x[12];
  assign t[284] = t[338] ^ x[18];
  assign t[285] = t[339] ^ x[17];
  assign t[286] = t[340] ^ x[21];
  assign t[287] = t[341] ^ x[20];
  assign t[288] = t[342] ^ x[24];
  assign t[289] = t[343] ^ x[23];
  assign t[28] = t[42] ^ t[43];
  assign t[290] = t[344] ^ x[27];
  assign t[291] = t[345] ^ x[26];
  assign t[292] = t[346] ^ x[30];
  assign t[293] = t[347] ^ x[29];
  assign t[294] = t[348] ^ x[33];
  assign t[295] = t[349] ^ x[32];
  assign t[296] = t[350] ^ x[36];
  assign t[297] = t[351] ^ x[35];
  assign t[298] = t[352] ^ x[39];
  assign t[299] = t[353] ^ x[38];
  assign t[29] = t[44] ^ t[45];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[42];
  assign t[301] = t[355] ^ x[41];
  assign t[302] = t[356] ^ x[45];
  assign t[303] = t[357] ^ x[44];
  assign t[304] = t[358] ^ x[48];
  assign t[305] = t[359] ^ x[47];
  assign t[306] = t[360] ^ x[51];
  assign t[307] = t[361] ^ x[50];
  assign t[308] = t[362] ^ x[54];
  assign t[309] = t[363] ^ x[53];
  assign t[30] = t[46] & t[47];
  assign t[310] = t[364] ^ x[57];
  assign t[311] = t[365] ^ x[56];
  assign t[312] = t[366] ^ x[60];
  assign t[313] = t[367] ^ x[59];
  assign t[314] = t[368] ^ x[65];
  assign t[315] = t[369] ^ x[64];
  assign t[316] = t[370] ^ x[68];
  assign t[317] = t[371] ^ x[67];
  assign t[318] = t[372] ^ x[71];
  assign t[319] = t[373] ^ x[70];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[74];
  assign t[321] = t[375] ^ x[73];
  assign t[322] = t[376] ^ x[77];
  assign t[323] = t[377] ^ x[76];
  assign t[324] = t[378] ^ x[82];
  assign t[325] = t[379] ^ x[81];
  assign t[326] = t[380] ^ x[89];
  assign t[327] = t[381] ^ x[88];
  assign t[328] = t[382] ^ x[92];
  assign t[329] = t[383] ^ x[91];
  assign t[32] = ~(t[50]);
  assign t[330] = (x[2]);
  assign t[331] = (x[2]);
  assign t[332] = (x[5]);
  assign t[333] = (x[5]);
  assign t[334] = (x[8]);
  assign t[335] = (x[8]);
  assign t[336] = (x[11]);
  assign t[337] = (x[11]);
  assign t[338] = (x[16]);
  assign t[339] = (x[16]);
  assign t[33] = ~(t[201]);
  assign t[340] = (x[19]);
  assign t[341] = (x[19]);
  assign t[342] = (x[22]);
  assign t[343] = (x[22]);
  assign t[344] = (x[25]);
  assign t[345] = (x[25]);
  assign t[346] = (x[28]);
  assign t[347] = (x[28]);
  assign t[348] = (x[31]);
  assign t[349] = (x[31]);
  assign t[34] = ~(t[51] ^ t[52]);
  assign t[350] = (x[34]);
  assign t[351] = (x[34]);
  assign t[352] = (x[37]);
  assign t[353] = (x[37]);
  assign t[354] = (x[40]);
  assign t[355] = (x[40]);
  assign t[356] = (x[43]);
  assign t[357] = (x[43]);
  assign t[358] = (x[46]);
  assign t[359] = (x[46]);
  assign t[35] = t[53] ^ t[54];
  assign t[360] = (x[49]);
  assign t[361] = (x[49]);
  assign t[362] = (x[52]);
  assign t[363] = (x[52]);
  assign t[364] = (x[55]);
  assign t[365] = (x[55]);
  assign t[366] = (x[58]);
  assign t[367] = (x[58]);
  assign t[368] = (x[63]);
  assign t[369] = (x[63]);
  assign t[36] = t[55] ^ t[56];
  assign t[370] = (x[66]);
  assign t[371] = (x[66]);
  assign t[372] = (x[69]);
  assign t[373] = (x[69]);
  assign t[374] = (x[72]);
  assign t[375] = (x[72]);
  assign t[376] = (x[75]);
  assign t[377] = (x[75]);
  assign t[378] = (x[80]);
  assign t[379] = (x[80]);
  assign t[37] = t[57] ^ t[43];
  assign t[380] = (x[87]);
  assign t[381] = (x[87]);
  assign t[382] = (x[90]);
  assign t[383] = (x[90]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[60] ^ t[18];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[9] ? t[63] : t[202];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[68];
  assign t[45] = ~t[69];
  assign t[46] = ~(t[29] ^ t[70]);
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[203] | t[75];
  assign t[4] = t[9] ? t[10] : t[195];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[71] ^ t[85];
  assign t[56] = t[82] ^ t[86];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] ^ t[61];
  assign t[59] = t[90] & t[91];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[94] ? t[95] : t[204];
  assign t[62] = t[96] ^ t[97];
  assign t[63] = t[202] ^ t[98];
  assign t[64] = t[99] & t[100];
  assign t[65] = t[101] & t[102];
  assign t[66] = ~(t[57] ^ t[42]);
  assign t[67] = t[103] ^ t[102];
  assign t[68] = t[9] ? t[104] : t[205];
  assign t[69] = t[9] ? t[105] : t[206];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[106] ^ t[107];
  assign t[71] = t[45] ^ t[108];
  assign t[72] = t[109];
  assign t[73] = ~(t[75] & t[110]);
  assign t[74] = ~(t[207] ^ t[111]);
  assign t[75] = ~(t[112] & t[113]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[17] ^ t[114];
  assign t[78] = ~(t[115] ^ t[116]);
  assign t[79] = t[117] ^ t[107];
  assign t[7] = t[15] ^ t[16];
  assign t[80] = t[108] ^ t[118];
  assign t[81] = t[9] ? t[119] : t[208];
  assign t[82] = t[9] ? t[120] : t[209];
  assign t[83] = ~(t[121]);
  assign t[84] = t[9] ? t[122] : t[210];
  assign t[85] = t[70] ^ t[123];
  assign t[86] = t[124] ^ t[125];
  assign t[87] = t[9] ? t[126] : t[211];
  assign t[88] = t[198] ^ t[127];
  assign t[89] = t[94] ? t[128] : t[212];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = ~(t[129]);
  assign t[91] = t[94] ? t[130] : t[213];
  assign t[92] = t[121] ^ t[82];
  assign t[93] = t[124] ^ t[131];
  assign t[94] = ~(t[19]);
  assign t[95] = t[204] ^ t[132];
  assign t[96] = t[133] ^ t[59];
  assign t[97] = t[134] & t[135];
  assign t[98] = t[136] ? x[62] : x[61];
  assign t[99] = ~(t[137]);
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [116:0] x;
 output y;

 wire [378:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~t[134];
  assign t[101] = t[125] ^ t[60];
  assign t[102] = t[135] ? t[136] : t[205];
  assign t[103] = t[135] ? t[137] : t[206];
  assign t[104] = ~(t[69] ^ t[138]);
  assign t[105] = t[139] ^ t[140];
  assign t[106] = t[141] & t[142];
  assign t[107] = ~(t[106] ^ t[143]);
  assign t[108] = t[19] ^ t[144];
  assign t[109] = ~(t[145] & t[146]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[147] ^ t[207];
  assign t[111] = ~(t[203]);
  assign t[112] = t[148] & t[147];
  assign t[113] = ~(t[50]);
  assign t[114] = t[113] ? x[65] : x[64];
  assign t[115] = t[102] ^ t[121];
  assign t[116] = t[149] & t[140];
  assign t[117] = t[33] ^ t[55];
  assign t[118] = t[150] & t[151];
  assign t[119] = t[126] ^ t[152];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[153] ^ t[90];
  assign t[121] = t[135] ? t[154] : t[208];
  assign t[122] = t[138] ^ t[70];
  assign t[123] = t[27] ? t[155] : t[209];
  assign t[124] = t[27] ? t[156] : t[210];
  assign t[125] = t[157] ^ t[158];
  assign t[126] = t[87] ^ t[100];
  assign t[127] = t[159];
  assign t[128] = ~(t[153] ^ t[42]);
  assign t[129] = t[23] ^ t[96];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[28] ? x[76] : x[75];
  assign t[131] = t[76] ? x[78] : x[77];
  assign t[132] = t[8] ? t[160] : t[211];
  assign t[133] = t[8] ? t[161] : t[212];
  assign t[134] = t[27] ? t[162] : t[213];
  assign t[135] = ~(t[15]);
  assign t[136] = t[205] ^ t[163];
  assign t[137] = t[206] ^ t[164];
  assign t[138] = t[165] ^ t[116];
  assign t[139] = t[103] ^ t[121];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[135] ? t[166] : t[214];
  assign t[141] = ~(t[144]);
  assign t[142] = ~(t[33]);
  assign t[143] = t[46] ^ t[33];
  assign t[144] = t[36] ^ t[55];
  assign t[145] = ~(t[148] | t[147]);
  assign t[146] = ~(t[167] | t[111]);
  assign t[147] = ~(t[215]);
  assign t[148] = ~(t[207]);
  assign t[149] = ~(t[103]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[117] ^ t[71]);
  assign t[151] = t[46] ^ t[36];
  assign t[152] = t[125] ^ t[168];
  assign t[153] = t[132] ^ t[40];
  assign t[154] = t[208] ^ t[169];
  assign t[155] = t[209] ^ t[170];
  assign t[156] = t[210] ^ t[171];
  assign t[157] = t[172] & t[173];
  assign t[158] = t[174] & t[127];
  assign t[159] = t[27] ? t[175] : t[216];
  assign t[15] = ~(t[27]);
  assign t[160] = t[211] ^ t[176];
  assign t[161] = t[212] ^ t[177];
  assign t[162] = t[213] ^ t[178];
  assign t[163] = t[179] ? x[98] : x[97];
  assign t[164] = t[179] ? x[100] : x[99];
  assign t[165] = t[180] & t[181];
  assign t[166] = t[214] ^ t[182];
  assign t[167] = ~(t[198]);
  assign t[168] = t[183] & t[184];
  assign t[169] = t[179] ? x[102] : x[101];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[76] ? x[104] : x[103];
  assign t[171] = t[28] ? x[106] : x[105];
  assign t[172] = ~(t[185]);
  assign t[173] = ~(t[86]);
  assign t[174] = ~(t[87]);
  assign t[175] = t[216] ^ t[186];
  assign t[176] = t[76] ? x[108] : x[107];
  assign t[177] = t[28] ? x[110] : x[109];
  assign t[178] = t[76] ? x[112] : x[111];
  assign t[179] = ~(t[50]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[187]);
  assign t[181] = ~(t[102]);
  assign t[182] = t[179] ? x[114] : x[113];
  assign t[183] = ~(t[157] ^ t[188]);
  assign t[184] = t[189] ^ t[185];
  assign t[185] = t[127] ^ t[87];
  assign t[186] = t[113] ? x[116] : x[115];
  assign t[187] = t[140] ^ t[103];
  assign t[188] = t[126] ^ t[86];
  assign t[189] = t[86] ^ t[100];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] & t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = t[244] ^ x[4];
  assign t[218] = t[245] ^ x[9];
  assign t[219] = t[246] ^ x[12];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[15];
  assign t[221] = t[248] ^ x[18];
  assign t[222] = t[249] ^ x[21];
  assign t[223] = t[250] ^ x[24];
  assign t[224] = t[251] ^ x[27];
  assign t[225] = t[252] ^ x[30];
  assign t[226] = t[253] ^ x[33];
  assign t[227] = t[254] ^ x[36];
  assign t[228] = t[255] ^ x[39];
  assign t[229] = t[256] ^ x[42];
  assign t[22] = ~(t[26] ^ t[39]);
  assign t[230] = t[257] ^ x[45];
  assign t[231] = t[258] ^ x[48];
  assign t[232] = t[259] ^ x[57];
  assign t[233] = t[260] ^ x[60];
  assign t[234] = t[261] ^ x[63];
  assign t[235] = t[262] ^ x[68];
  assign t[236] = t[263] ^ x[71];
  assign t[237] = t[264] ^ x[74];
  assign t[238] = t[265] ^ x[81];
  assign t[239] = t[266] ^ x[84];
  assign t[23] = t[40] ^ t[41];
  assign t[240] = t[267] ^ x[87];
  assign t[241] = t[268] ^ x[90];
  assign t[242] = t[269] ^ x[93];
  assign t[243] = t[270] ^ x[96];
  assign t[244] = (t[271] & ~t[272]);
  assign t[245] = (t[273] & ~t[274]);
  assign t[246] = (t[275] & ~t[276]);
  assign t[247] = (t[277] & ~t[278]);
  assign t[248] = (t[279] & ~t[280]);
  assign t[249] = (t[281] & ~t[282]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[283] & ~t[284]);
  assign t[251] = (t[285] & ~t[286]);
  assign t[252] = (t[287] & ~t[288]);
  assign t[253] = (t[289] & ~t[290]);
  assign t[254] = (t[291] & ~t[292]);
  assign t[255] = (t[293] & ~t[294]);
  assign t[256] = (t[295] & ~t[296]);
  assign t[257] = (t[297] & ~t[298]);
  assign t[258] = (t[299] & ~t[300]);
  assign t[259] = (t[301] & ~t[302]);
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[260] = (t[303] & ~t[304]);
  assign t[261] = (t[305] & ~t[306]);
  assign t[262] = (t[307] & ~t[308]);
  assign t[263] = (t[309] & ~t[310]);
  assign t[264] = (t[311] & ~t[312]);
  assign t[265] = (t[313] & ~t[314]);
  assign t[266] = (t[315] & ~t[316]);
  assign t[267] = (t[317] & ~t[318]);
  assign t[268] = (t[319] & ~t[320]);
  assign t[269] = (t[321] & ~t[322]);
  assign t[26] = t[46] ^ t[47];
  assign t[270] = (t[323] & ~t[324]);
  assign t[271] = t[325] ^ x[4];
  assign t[272] = t[326] ^ x[3];
  assign t[273] = t[327] ^ x[9];
  assign t[274] = t[328] ^ x[8];
  assign t[275] = t[329] ^ x[12];
  assign t[276] = t[330] ^ x[11];
  assign t[277] = t[331] ^ x[15];
  assign t[278] = t[332] ^ x[14];
  assign t[279] = t[333] ^ x[18];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[17];
  assign t[281] = t[335] ^ x[21];
  assign t[282] = t[336] ^ x[20];
  assign t[283] = t[337] ^ x[24];
  assign t[284] = t[338] ^ x[23];
  assign t[285] = t[339] ^ x[27];
  assign t[286] = t[340] ^ x[26];
  assign t[287] = t[341] ^ x[30];
  assign t[288] = t[342] ^ x[29];
  assign t[289] = t[343] ^ x[33];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[32];
  assign t[291] = t[345] ^ x[36];
  assign t[292] = t[346] ^ x[35];
  assign t[293] = t[347] ^ x[39];
  assign t[294] = t[348] ^ x[38];
  assign t[295] = t[349] ^ x[42];
  assign t[296] = t[350] ^ x[41];
  assign t[297] = t[351] ^ x[45];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[48];
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[47];
  assign t[301] = t[355] ^ x[57];
  assign t[302] = t[356] ^ x[56];
  assign t[303] = t[357] ^ x[60];
  assign t[304] = t[358] ^ x[59];
  assign t[305] = t[359] ^ x[63];
  assign t[306] = t[360] ^ x[62];
  assign t[307] = t[361] ^ x[68];
  assign t[308] = t[362] ^ x[67];
  assign t[309] = t[363] ^ x[71];
  assign t[30] = ~(t[192]);
  assign t[310] = t[364] ^ x[70];
  assign t[311] = t[365] ^ x[74];
  assign t[312] = t[366] ^ x[73];
  assign t[313] = t[367] ^ x[81];
  assign t[314] = t[368] ^ x[80];
  assign t[315] = t[369] ^ x[84];
  assign t[316] = t[370] ^ x[83];
  assign t[317] = t[371] ^ x[87];
  assign t[318] = t[372] ^ x[86];
  assign t[319] = t[373] ^ x[90];
  assign t[31] = ~(t[193]);
  assign t[320] = t[374] ^ x[89];
  assign t[321] = t[375] ^ x[93];
  assign t[322] = t[376] ^ x[92];
  assign t[323] = t[377] ^ x[96];
  assign t[324] = t[378] ^ x[95];
  assign t[325] = (x[2]);
  assign t[326] = (x[2]);
  assign t[327] = (x[7]);
  assign t[328] = (x[7]);
  assign t[329] = (x[10]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[10]);
  assign t[331] = (x[13]);
  assign t[332] = (x[13]);
  assign t[333] = (x[16]);
  assign t[334] = (x[16]);
  assign t[335] = (x[19]);
  assign t[336] = (x[19]);
  assign t[337] = (x[22]);
  assign t[338] = (x[22]);
  assign t[339] = (x[25]);
  assign t[33] = t[8] ? t[53] : t[194];
  assign t[340] = (x[25]);
  assign t[341] = (x[28]);
  assign t[342] = (x[28]);
  assign t[343] = (x[31]);
  assign t[344] = (x[31]);
  assign t[345] = (x[34]);
  assign t[346] = (x[34]);
  assign t[347] = (x[37]);
  assign t[348] = (x[37]);
  assign t[349] = (x[40]);
  assign t[34] = t[8] ? t[54] : t[195];
  assign t[350] = (x[40]);
  assign t[351] = (x[43]);
  assign t[352] = (x[43]);
  assign t[353] = (x[46]);
  assign t[354] = (x[46]);
  assign t[355] = (x[55]);
  assign t[356] = (x[55]);
  assign t[357] = (x[58]);
  assign t[358] = (x[58]);
  assign t[359] = (x[61]);
  assign t[35] = ~(t[55]);
  assign t[360] = (x[61]);
  assign t[361] = (x[66]);
  assign t[362] = (x[66]);
  assign t[363] = (x[69]);
  assign t[364] = (x[69]);
  assign t[365] = (x[72]);
  assign t[366] = (x[72]);
  assign t[367] = (x[79]);
  assign t[368] = (x[79]);
  assign t[369] = (x[82]);
  assign t[36] = t[8] ? t[56] : t[196];
  assign t[370] = (x[82]);
  assign t[371] = (x[85]);
  assign t[372] = (x[85]);
  assign t[373] = (x[88]);
  assign t[374] = (x[88]);
  assign t[375] = (x[91]);
  assign t[376] = (x[91]);
  assign t[377] = (x[94]);
  assign t[378] = (x[94]);
  assign t[37] = ~(t[57] ^ t[58]);
  assign t[38] = t[59] ^ t[60];
  assign t[39] = t[41] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[191] ^ t[62];
  assign t[41] = t[197] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[13] ^ t[68];
  assign t[45] = t[69] ^ t[70];
  assign t[46] = t[55] ^ t[34];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[198] | t[75];
  assign t[4] = t[8] ? t[9] : t[190];
  assign t[50] = ~(t[76]);
  assign t[51] = ~(t[199]);
  assign t[52] = ~(t[77] & t[197]);
  assign t[53] = t[194] ^ t[78];
  assign t[54] = t[195] ^ t[79];
  assign t[55] = t[8] ? t[80] : t[200];
  assign t[56] = t[196] ^ t[81];
  assign t[57] = t[82] ^ t[83];
  assign t[58] = ~(t[84] ^ t[85]);
  assign t[59] = t[86] ^ t[87];
  assign t[5] = ~(t[10]);
  assign t[60] = t[88] & t[89];
  assign t[61] = t[42] ^ t[90];
  assign t[62] = t[27] ? t[91] : t[201];
  assign t[63] = t[8] ? t[92] : t[202];
  assign t[64] = t[93] & t[94];
  assign t[65] = t[95] & t[96];
  assign t[66] = ~(t[64] ^ t[97]);
  assign t[67] = t[98] ^ t[99];
  assign t[68] = t[100] ^ t[101];
  assign t[69] = t[102] ^ t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[104] & t[105];
  assign t[71] = t[106] ^ t[20];
  assign t[72] = t[107] & t[108];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[203] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[49]);
  assign t[77] = ~(t[204]);
  assign t[78] = t[113] ? x[50] : x[49];
  assign t[79] = t[113] ? x[52] : x[51];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[200] ^ t[114];
  assign t[81] = t[113] ? x[54] : x[53];
  assign t[82] = t[115] ^ t[116];
  assign t[83] = t[117] ^ t[118];
  assign t[84] = t[119] ^ t[120];
  assign t[85] = t[121] ^ t[122];
  assign t[86] = ~t[123];
  assign t[87] = t[124];
  assign t[88] = ~(t[59] ^ t[125]);
  assign t[89] = t[126] ^ t[127];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] & t[129];
  assign t[91] = t[201] ^ t[130];
  assign t[92] = t[202] ^ t[131];
  assign t[93] = ~(t[99]);
  assign t[94] = ~(t[132]);
  assign t[95] = ~(t[40]);
  assign t[96] = t[192] ^ t[133];
  assign t[97] = t[23] ^ t[132];
  assign t[98] = t[132] ^ t[41];
  assign t[99] = t[96] ^ t[40];
  assign t[9] = t[190] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [116:0] x;
 output y;

 wire [378:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~t[134];
  assign t[101] = t[125] ^ t[60];
  assign t[102] = t[135] ? t[136] : t[205];
  assign t[103] = t[135] ? t[137] : t[206];
  assign t[104] = ~(t[69] ^ t[138]);
  assign t[105] = t[139] ^ t[140];
  assign t[106] = t[141] & t[142];
  assign t[107] = ~(t[106] ^ t[143]);
  assign t[108] = t[19] ^ t[144];
  assign t[109] = ~(t[145] & t[146]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[147] ^ t[207];
  assign t[111] = ~(t[203]);
  assign t[112] = t[148] & t[147];
  assign t[113] = ~(t[50]);
  assign t[114] = t[113] ? x[65] : x[64];
  assign t[115] = t[102] ^ t[121];
  assign t[116] = t[149] & t[140];
  assign t[117] = t[33] ^ t[55];
  assign t[118] = t[150] & t[151];
  assign t[119] = t[126] ^ t[152];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[153] ^ t[90];
  assign t[121] = t[135] ? t[154] : t[208];
  assign t[122] = t[138] ^ t[70];
  assign t[123] = t[27] ? t[155] : t[209];
  assign t[124] = t[27] ? t[156] : t[210];
  assign t[125] = t[157] ^ t[158];
  assign t[126] = t[87] ^ t[100];
  assign t[127] = t[159];
  assign t[128] = ~(t[153] ^ t[42]);
  assign t[129] = t[23] ^ t[96];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[28] ? x[76] : x[75];
  assign t[131] = t[76] ? x[78] : x[77];
  assign t[132] = t[8] ? t[160] : t[211];
  assign t[133] = t[8] ? t[161] : t[212];
  assign t[134] = t[27] ? t[162] : t[213];
  assign t[135] = ~(t[15]);
  assign t[136] = t[205] ^ t[163];
  assign t[137] = t[206] ^ t[164];
  assign t[138] = t[165] ^ t[116];
  assign t[139] = t[103] ^ t[121];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[135] ? t[166] : t[214];
  assign t[141] = ~(t[144]);
  assign t[142] = ~(t[33]);
  assign t[143] = t[46] ^ t[33];
  assign t[144] = t[36] ^ t[55];
  assign t[145] = ~(t[148] | t[147]);
  assign t[146] = ~(t[167] | t[111]);
  assign t[147] = ~(t[215]);
  assign t[148] = ~(t[207]);
  assign t[149] = ~(t[103]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[117] ^ t[71]);
  assign t[151] = t[46] ^ t[36];
  assign t[152] = t[125] ^ t[168];
  assign t[153] = t[132] ^ t[40];
  assign t[154] = t[208] ^ t[169];
  assign t[155] = t[209] ^ t[170];
  assign t[156] = t[210] ^ t[171];
  assign t[157] = t[172] & t[173];
  assign t[158] = t[174] & t[127];
  assign t[159] = t[27] ? t[175] : t[216];
  assign t[15] = ~(t[27]);
  assign t[160] = t[211] ^ t[176];
  assign t[161] = t[212] ^ t[177];
  assign t[162] = t[213] ^ t[178];
  assign t[163] = t[179] ? x[98] : x[97];
  assign t[164] = t[179] ? x[100] : x[99];
  assign t[165] = t[180] & t[181];
  assign t[166] = t[214] ^ t[182];
  assign t[167] = ~(t[198]);
  assign t[168] = t[183] & t[184];
  assign t[169] = t[179] ? x[102] : x[101];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[76] ? x[104] : x[103];
  assign t[171] = t[28] ? x[106] : x[105];
  assign t[172] = ~(t[185]);
  assign t[173] = ~(t[86]);
  assign t[174] = ~(t[87]);
  assign t[175] = t[216] ^ t[186];
  assign t[176] = t[76] ? x[108] : x[107];
  assign t[177] = t[28] ? x[110] : x[109];
  assign t[178] = t[76] ? x[112] : x[111];
  assign t[179] = ~(t[50]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[187]);
  assign t[181] = ~(t[102]);
  assign t[182] = t[179] ? x[114] : x[113];
  assign t[183] = ~(t[157] ^ t[188]);
  assign t[184] = t[189] ^ t[185];
  assign t[185] = t[127] ^ t[87];
  assign t[186] = t[113] ? x[116] : x[115];
  assign t[187] = t[140] ^ t[103];
  assign t[188] = t[126] ^ t[86];
  assign t[189] = t[86] ^ t[100];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = (t[217]);
  assign t[191] = (t[218]);
  assign t[192] = (t[219]);
  assign t[193] = (t[220]);
  assign t[194] = (t[221]);
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] & t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = t[244] ^ x[4];
  assign t[218] = t[245] ^ x[9];
  assign t[219] = t[246] ^ x[12];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[247] ^ x[15];
  assign t[221] = t[248] ^ x[18];
  assign t[222] = t[249] ^ x[21];
  assign t[223] = t[250] ^ x[24];
  assign t[224] = t[251] ^ x[27];
  assign t[225] = t[252] ^ x[30];
  assign t[226] = t[253] ^ x[33];
  assign t[227] = t[254] ^ x[36];
  assign t[228] = t[255] ^ x[39];
  assign t[229] = t[256] ^ x[42];
  assign t[22] = ~(t[26] ^ t[39]);
  assign t[230] = t[257] ^ x[45];
  assign t[231] = t[258] ^ x[48];
  assign t[232] = t[259] ^ x[57];
  assign t[233] = t[260] ^ x[60];
  assign t[234] = t[261] ^ x[63];
  assign t[235] = t[262] ^ x[68];
  assign t[236] = t[263] ^ x[71];
  assign t[237] = t[264] ^ x[74];
  assign t[238] = t[265] ^ x[81];
  assign t[239] = t[266] ^ x[84];
  assign t[23] = t[40] ^ t[41];
  assign t[240] = t[267] ^ x[87];
  assign t[241] = t[268] ^ x[90];
  assign t[242] = t[269] ^ x[93];
  assign t[243] = t[270] ^ x[96];
  assign t[244] = (t[271] & ~t[272]);
  assign t[245] = (t[273] & ~t[274]);
  assign t[246] = (t[275] & ~t[276]);
  assign t[247] = (t[277] & ~t[278]);
  assign t[248] = (t[279] & ~t[280]);
  assign t[249] = (t[281] & ~t[282]);
  assign t[24] = t[42] ^ t[43];
  assign t[250] = (t[283] & ~t[284]);
  assign t[251] = (t[285] & ~t[286]);
  assign t[252] = (t[287] & ~t[288]);
  assign t[253] = (t[289] & ~t[290]);
  assign t[254] = (t[291] & ~t[292]);
  assign t[255] = (t[293] & ~t[294]);
  assign t[256] = (t[295] & ~t[296]);
  assign t[257] = (t[297] & ~t[298]);
  assign t[258] = (t[299] & ~t[300]);
  assign t[259] = (t[301] & ~t[302]);
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[260] = (t[303] & ~t[304]);
  assign t[261] = (t[305] & ~t[306]);
  assign t[262] = (t[307] & ~t[308]);
  assign t[263] = (t[309] & ~t[310]);
  assign t[264] = (t[311] & ~t[312]);
  assign t[265] = (t[313] & ~t[314]);
  assign t[266] = (t[315] & ~t[316]);
  assign t[267] = (t[317] & ~t[318]);
  assign t[268] = (t[319] & ~t[320]);
  assign t[269] = (t[321] & ~t[322]);
  assign t[26] = t[46] ^ t[47];
  assign t[270] = (t[323] & ~t[324]);
  assign t[271] = t[325] ^ x[4];
  assign t[272] = t[326] ^ x[3];
  assign t[273] = t[327] ^ x[9];
  assign t[274] = t[328] ^ x[8];
  assign t[275] = t[329] ^ x[12];
  assign t[276] = t[330] ^ x[11];
  assign t[277] = t[331] ^ x[15];
  assign t[278] = t[332] ^ x[14];
  assign t[279] = t[333] ^ x[18];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[17];
  assign t[281] = t[335] ^ x[21];
  assign t[282] = t[336] ^ x[20];
  assign t[283] = t[337] ^ x[24];
  assign t[284] = t[338] ^ x[23];
  assign t[285] = t[339] ^ x[27];
  assign t[286] = t[340] ^ x[26];
  assign t[287] = t[341] ^ x[30];
  assign t[288] = t[342] ^ x[29];
  assign t[289] = t[343] ^ x[33];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[32];
  assign t[291] = t[345] ^ x[36];
  assign t[292] = t[346] ^ x[35];
  assign t[293] = t[347] ^ x[39];
  assign t[294] = t[348] ^ x[38];
  assign t[295] = t[349] ^ x[42];
  assign t[296] = t[350] ^ x[41];
  assign t[297] = t[351] ^ x[45];
  assign t[298] = t[352] ^ x[44];
  assign t[299] = t[353] ^ x[48];
  assign t[29] = ~(t[191]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[47];
  assign t[301] = t[355] ^ x[57];
  assign t[302] = t[356] ^ x[56];
  assign t[303] = t[357] ^ x[60];
  assign t[304] = t[358] ^ x[59];
  assign t[305] = t[359] ^ x[63];
  assign t[306] = t[360] ^ x[62];
  assign t[307] = t[361] ^ x[68];
  assign t[308] = t[362] ^ x[67];
  assign t[309] = t[363] ^ x[71];
  assign t[30] = ~(t[192]);
  assign t[310] = t[364] ^ x[70];
  assign t[311] = t[365] ^ x[74];
  assign t[312] = t[366] ^ x[73];
  assign t[313] = t[367] ^ x[81];
  assign t[314] = t[368] ^ x[80];
  assign t[315] = t[369] ^ x[84];
  assign t[316] = t[370] ^ x[83];
  assign t[317] = t[371] ^ x[87];
  assign t[318] = t[372] ^ x[86];
  assign t[319] = t[373] ^ x[90];
  assign t[31] = ~(t[193]);
  assign t[320] = t[374] ^ x[89];
  assign t[321] = t[375] ^ x[93];
  assign t[322] = t[376] ^ x[92];
  assign t[323] = t[377] ^ x[96];
  assign t[324] = t[378] ^ x[95];
  assign t[325] = (x[2]);
  assign t[326] = (x[2]);
  assign t[327] = (x[7]);
  assign t[328] = (x[7]);
  assign t[329] = (x[10]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (x[10]);
  assign t[331] = (x[13]);
  assign t[332] = (x[13]);
  assign t[333] = (x[16]);
  assign t[334] = (x[16]);
  assign t[335] = (x[19]);
  assign t[336] = (x[19]);
  assign t[337] = (x[22]);
  assign t[338] = (x[22]);
  assign t[339] = (x[25]);
  assign t[33] = t[8] ? t[53] : t[194];
  assign t[340] = (x[25]);
  assign t[341] = (x[28]);
  assign t[342] = (x[28]);
  assign t[343] = (x[31]);
  assign t[344] = (x[31]);
  assign t[345] = (x[34]);
  assign t[346] = (x[34]);
  assign t[347] = (x[37]);
  assign t[348] = (x[37]);
  assign t[349] = (x[40]);
  assign t[34] = t[8] ? t[54] : t[195];
  assign t[350] = (x[40]);
  assign t[351] = (x[43]);
  assign t[352] = (x[43]);
  assign t[353] = (x[46]);
  assign t[354] = (x[46]);
  assign t[355] = (x[55]);
  assign t[356] = (x[55]);
  assign t[357] = (x[58]);
  assign t[358] = (x[58]);
  assign t[359] = (x[61]);
  assign t[35] = ~(t[55]);
  assign t[360] = (x[61]);
  assign t[361] = (x[66]);
  assign t[362] = (x[66]);
  assign t[363] = (x[69]);
  assign t[364] = (x[69]);
  assign t[365] = (x[72]);
  assign t[366] = (x[72]);
  assign t[367] = (x[79]);
  assign t[368] = (x[79]);
  assign t[369] = (x[82]);
  assign t[36] = t[8] ? t[56] : t[196];
  assign t[370] = (x[82]);
  assign t[371] = (x[85]);
  assign t[372] = (x[85]);
  assign t[373] = (x[88]);
  assign t[374] = (x[88]);
  assign t[375] = (x[91]);
  assign t[376] = (x[91]);
  assign t[377] = (x[94]);
  assign t[378] = (x[94]);
  assign t[37] = ~(t[57] ^ t[58]);
  assign t[38] = t[59] ^ t[60];
  assign t[39] = t[41] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[191] ^ t[62];
  assign t[41] = t[197] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[13] ^ t[68];
  assign t[45] = t[69] ^ t[70];
  assign t[46] = t[55] ^ t[34];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[198] | t[75];
  assign t[4] = t[8] ? t[9] : t[190];
  assign t[50] = ~(t[76]);
  assign t[51] = ~(t[199]);
  assign t[52] = ~(t[77] & t[197]);
  assign t[53] = t[194] ^ t[78];
  assign t[54] = t[195] ^ t[79];
  assign t[55] = t[8] ? t[80] : t[200];
  assign t[56] = t[196] ^ t[81];
  assign t[57] = t[82] ^ t[83];
  assign t[58] = ~(t[84] ^ t[85]);
  assign t[59] = t[86] ^ t[87];
  assign t[5] = ~(t[10]);
  assign t[60] = t[88] & t[89];
  assign t[61] = t[42] ^ t[90];
  assign t[62] = t[27] ? t[91] : t[201];
  assign t[63] = t[8] ? t[92] : t[202];
  assign t[64] = t[93] & t[94];
  assign t[65] = t[95] & t[96];
  assign t[66] = ~(t[64] ^ t[97]);
  assign t[67] = t[98] ^ t[99];
  assign t[68] = t[100] ^ t[101];
  assign t[69] = t[102] ^ t[103];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = t[104] & t[105];
  assign t[71] = t[106] ^ t[20];
  assign t[72] = t[107] & t[108];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[203] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[49]);
  assign t[77] = ~(t[204]);
  assign t[78] = t[113] ? x[50] : x[49];
  assign t[79] = t[113] ? x[52] : x[51];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[200] ^ t[114];
  assign t[81] = t[113] ? x[54] : x[53];
  assign t[82] = t[115] ^ t[116];
  assign t[83] = t[117] ^ t[118];
  assign t[84] = t[119] ^ t[120];
  assign t[85] = t[121] ^ t[122];
  assign t[86] = ~t[123];
  assign t[87] = t[124];
  assign t[88] = ~(t[59] ^ t[125]);
  assign t[89] = t[126] ^ t[127];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] & t[129];
  assign t[91] = t[201] ^ t[130];
  assign t[92] = t[202] ^ t[131];
  assign t[93] = ~(t[99]);
  assign t[94] = ~(t[132]);
  assign t[95] = ~(t[40]);
  assign t[96] = t[192] ^ t[133];
  assign t[97] = t[23] ^ t[132];
  assign t[98] = t[132] ^ t[41];
  assign t[99] = t[96] ^ t[40];
  assign t[9] = t[190] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [116:0] x;
 output y;

 wire [396:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~t[137];
  assign t[101] = t[138] ^ t[121];
  assign t[102] = t[139] & t[140];
  assign t[103] = t[218] ^ t[141];
  assign t[104] = t[142] ^ t[143];
  assign t[105] = t[42] ^ t[144];
  assign t[106] = t[145] ^ t[146];
  assign t[107] = ~t[147];
  assign t[108] = ~(t[72] ^ t[101]);
  assign t[109] = t[66] ^ t[148];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[149] & t[150];
  assign t[111] = ~(t[151] & t[152]);
  assign t[112] = t[153] ^ t[224];
  assign t[113] = ~(t[219]);
  assign t[114] = t[154] & t[153];
  assign t[115] = t[100] ^ t[155];
  assign t[116] = t[156] ^ t[157];
  assign t[117] = t[158] & t[159];
  assign t[118] = t[157] ^ t[145];
  assign t[119] = t[160] ^ t[161];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[107] ^ t[100];
  assign t[121] = t[162] & t[148];
  assign t[122] = t[163] ? x[56] : x[55];
  assign t[123] = t[163] ? x[58] : x[57];
  assign t[124] = t[164] & t[165];
  assign t[125] = t[166] & t[88];
  assign t[126] = t[221] ^ t[167];
  assign t[127] = t[222] ^ t[168];
  assign t[128] = ~(t[131]);
  assign t[129] = ~(t[96]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[37] ^ t[96];
  assign t[131] = t[98] ^ t[59];
  assign t[132] = t[79] ? x[60] : x[59];
  assign t[133] = t[96] ^ t[59];
  assign t[134] = t[223] ^ t[169];
  assign t[135] = t[8] ? t[170] : t[225];
  assign t[136] = t[27] ? t[171] : t[226];
  assign t[137] = t[27] ? t[172] : t[227];
  assign t[138] = t[173] & t[174];
  assign t[139] = ~(t[138] ^ t[175]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[120] ^ t[176];
  assign t[141] = t[163] ? x[71] : x[70];
  assign t[142] = t[156] ^ t[145];
  assign t[143] = t[177] & t[178];
  assign t[144] = t[133] ^ t[63];
  assign t[145] = t[179] ? t[180] : t[228];
  assign t[146] = t[160] ^ t[117];
  assign t[147] = t[27] ? t[181] : t[229];
  assign t[148] = t[182];
  assign t[149] = ~(t[124] ^ t[183]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[184] ^ t[185];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[186] | t[113]);
  assign t[153] = ~(t[230]);
  assign t[154] = ~(t[224]);
  assign t[155] = t[101] ^ t[73];
  assign t[156] = t[179] ? t[187] : t[231];
  assign t[157] = t[179] ? t[188] : t[232];
  assign t[158] = ~(t[116] ^ t[160]);
  assign t[159] = t[118] ^ t[178];
  assign t[15] = ~(t[27]);
  assign t[160] = t[189] ^ t[143];
  assign t[161] = t[190] & t[191];
  assign t[162] = ~(t[99]);
  assign t[163] = ~(t[49]);
  assign t[164] = ~(t[185]);
  assign t[165] = ~(t[55]);
  assign t[166] = ~(t[56]);
  assign t[167] = t[163] ? x[88] : x[87];
  assign t[168] = t[28] ? x[90] : x[89];
  assign t[169] = t[79] ? x[92] : x[91];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[225] ^ t[192];
  assign t[171] = t[226] ^ t[193];
  assign t[172] = t[227] ^ t[194];
  assign t[173] = ~(t[176]);
  assign t[174] = ~(t[107]);
  assign t[175] = t[66] ^ t[107];
  assign t[176] = t[148] ^ t[99];
  assign t[177] = ~(t[157]);
  assign t[178] = t[179] ? t[195] : t[233];
  assign t[179] = ~(t[15]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[228] ^ t[196];
  assign t[181] = t[229] ^ t[197];
  assign t[182] = t[27] ? t[198] : t[234];
  assign t[183] = t[74] ^ t[55];
  assign t[184] = t[55] ^ t[68];
  assign t[185] = t[88] ^ t[56];
  assign t[186] = ~(t[213]);
  assign t[187] = t[231] ^ t[199];
  assign t[188] = t[232] ^ t[200];
  assign t[189] = t[201] & t[202];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = ~(t[189] ^ t[203]);
  assign t[191] = t[142] ^ t[204];
  assign t[192] = t[28] ? x[100] : x[99];
  assign t[193] = t[28] ? x[102] : x[101];
  assign t[194] = t[79] ? x[104] : x[103];
  assign t[195] = t[233] ^ t[205];
  assign t[196] = t[206] ? x[106] : x[105];
  assign t[197] = t[79] ? x[108] : x[107];
  assign t[198] = t[234] ^ t[207];
  assign t[199] = t[206] ? x[110] : x[109];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[206] ? x[112] : x[111];
  assign t[201] = ~(t[204]);
  assign t[202] = ~(t[156]);
  assign t[203] = t[118] ^ t[156];
  assign t[204] = t[178] ^ t[157];
  assign t[205] = t[206] ? x[114] : x[113];
  assign t[206] = ~(t[49]);
  assign t[207] = t[163] ? x[116] : x[115];
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = t[262] ^ x[4];
  assign t[236] = t[263] ^ x[9];
  assign t[237] = t[264] ^ x[12];
  assign t[238] = t[265] ^ x[15];
  assign t[239] = t[266] ^ x[18];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[21];
  assign t[241] = t[268] ^ x[24];
  assign t[242] = t[269] ^ x[27];
  assign t[243] = t[270] ^ x[30];
  assign t[244] = t[271] ^ x[33];
  assign t[245] = t[272] ^ x[36];
  assign t[246] = t[273] ^ x[39];
  assign t[247] = t[274] ^ x[42];
  assign t[248] = t[275] ^ x[45];
  assign t[249] = t[276] ^ x[48];
  assign t[24] = ~(t[33] ^ t[43]);
  assign t[250] = t[277] ^ x[51];
  assign t[251] = t[278] ^ x[54];
  assign t[252] = t[279] ^ x[63];
  assign t[253] = t[280] ^ x[66];
  assign t[254] = t[281] ^ x[69];
  assign t[255] = t[282] ^ x[74];
  assign t[256] = t[283] ^ x[77];
  assign t[257] = t[284] ^ x[80];
  assign t[258] = t[285] ^ x[83];
  assign t[259] = t[286] ^ x[86];
  assign t[25] = t[44] ^ t[45];
  assign t[260] = t[287] ^ x[95];
  assign t[261] = t[288] ^ x[98];
  assign t[262] = (t[289] & ~t[290]);
  assign t[263] = (t[291] & ~t[292]);
  assign t[264] = (t[293] & ~t[294]);
  assign t[265] = (t[295] & ~t[296]);
  assign t[266] = (t[297] & ~t[298]);
  assign t[267] = (t[299] & ~t[300]);
  assign t[268] = (t[301] & ~t[302]);
  assign t[269] = (t[303] & ~t[304]);
  assign t[26] = ~(t[46] ^ t[22]);
  assign t[270] = (t[305] & ~t[306]);
  assign t[271] = (t[307] & ~t[308]);
  assign t[272] = (t[309] & ~t[310]);
  assign t[273] = (t[311] & ~t[312]);
  assign t[274] = (t[313] & ~t[314]);
  assign t[275] = (t[315] & ~t[316]);
  assign t[276] = (t[317] & ~t[318]);
  assign t[277] = (t[319] & ~t[320]);
  assign t[278] = (t[321] & ~t[322]);
  assign t[279] = (t[323] & ~t[324]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[325] & ~t[326]);
  assign t[281] = (t[327] & ~t[328]);
  assign t[282] = (t[329] & ~t[330]);
  assign t[283] = (t[331] & ~t[332]);
  assign t[284] = (t[333] & ~t[334]);
  assign t[285] = (t[335] & ~t[336]);
  assign t[286] = (t[337] & ~t[338]);
  assign t[287] = (t[339] & ~t[340]);
  assign t[288] = (t[341] & ~t[342]);
  assign t[289] = t[343] ^ x[4];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[3];
  assign t[291] = t[345] ^ x[9];
  assign t[292] = t[346] ^ x[8];
  assign t[293] = t[347] ^ x[12];
  assign t[294] = t[348] ^ x[11];
  assign t[295] = t[349] ^ x[15];
  assign t[296] = t[350] ^ x[14];
  assign t[297] = t[351] ^ x[18];
  assign t[298] = t[352] ^ x[17];
  assign t[299] = t[353] ^ x[21];
  assign t[29] = ~(t[209]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[20];
  assign t[301] = t[355] ^ x[24];
  assign t[302] = t[356] ^ x[23];
  assign t[303] = t[357] ^ x[27];
  assign t[304] = t[358] ^ x[26];
  assign t[305] = t[359] ^ x[30];
  assign t[306] = t[360] ^ x[29];
  assign t[307] = t[361] ^ x[33];
  assign t[308] = t[362] ^ x[32];
  assign t[309] = t[363] ^ x[36];
  assign t[30] = ~(t[210]);
  assign t[310] = t[364] ^ x[35];
  assign t[311] = t[365] ^ x[39];
  assign t[312] = t[366] ^ x[38];
  assign t[313] = t[367] ^ x[42];
  assign t[314] = t[368] ^ x[41];
  assign t[315] = t[369] ^ x[45];
  assign t[316] = t[370] ^ x[44];
  assign t[317] = t[371] ^ x[48];
  assign t[318] = t[372] ^ x[47];
  assign t[319] = t[373] ^ x[51];
  assign t[31] = ~(t[211]);
  assign t[320] = t[374] ^ x[50];
  assign t[321] = t[375] ^ x[54];
  assign t[322] = t[376] ^ x[53];
  assign t[323] = t[377] ^ x[63];
  assign t[324] = t[378] ^ x[62];
  assign t[325] = t[379] ^ x[66];
  assign t[326] = t[380] ^ x[65];
  assign t[327] = t[381] ^ x[69];
  assign t[328] = t[382] ^ x[68];
  assign t[329] = t[383] ^ x[74];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[73];
  assign t[331] = t[385] ^ x[77];
  assign t[332] = t[386] ^ x[76];
  assign t[333] = t[387] ^ x[80];
  assign t[334] = t[388] ^ x[79];
  assign t[335] = t[389] ^ x[83];
  assign t[336] = t[390] ^ x[82];
  assign t[337] = t[391] ^ x[86];
  assign t[338] = t[392] ^ x[85];
  assign t[339] = t[393] ^ x[95];
  assign t[33] = ~(t[52] ^ t[46]);
  assign t[340] = t[394] ^ x[94];
  assign t[341] = t[395] ^ x[98];
  assign t[342] = t[396] ^ x[97];
  assign t[343] = (x[2]);
  assign t[344] = (x[2]);
  assign t[345] = (x[7]);
  assign t[346] = (x[7]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[49]);
  assign t[374] = (x[49]);
  assign t[375] = (x[52]);
  assign t[376] = (x[52]);
  assign t[377] = (x[61]);
  assign t[378] = (x[61]);
  assign t[379] = (x[64]);
  assign t[37] = t[59] ^ t[39];
  assign t[380] = (x[64]);
  assign t[381] = (x[67]);
  assign t[382] = (x[67]);
  assign t[383] = (x[72]);
  assign t[384] = (x[72]);
  assign t[385] = (x[75]);
  assign t[386] = (x[75]);
  assign t[387] = (x[78]);
  assign t[388] = (x[78]);
  assign t[389] = (x[81]);
  assign t[38] = t[60] ^ t[61];
  assign t[390] = (x[81]);
  assign t[391] = (x[84]);
  assign t[392] = (x[84]);
  assign t[393] = (x[93]);
  assign t[394] = (x[93]);
  assign t[395] = (x[96]);
  assign t[396] = (x[96]);
  assign t[39] = t[212] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[60] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = ~(t[70] ^ t[71]);
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = t[213] | t[78];
  assign t[49] = ~(t[79]);
  assign t[4] = t[8] ? t[9] : t[208];
  assign t[50] = ~(t[214]);
  assign t[51] = ~(t[80] & t[212]);
  assign t[52] = ~(t[81] ^ t[82]);
  assign t[53] = t[83] ^ t[84];
  assign t[54] = ~(t[43] ^ t[22]);
  assign t[55] = t[8] ? t[85] : t[215];
  assign t[56] = t[8] ? t[86] : t[216];
  assign t[57] = ~(t[35] ^ t[87]);
  assign t[58] = t[74] ^ t[88];
  assign t[59] = t[209] ^ t[89];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[65];
  assign t[61] = t[91] & t[92];
  assign t[62] = t[8] ? t[93] : t[217];
  assign t[63] = t[94] & t[95];
  assign t[64] = t[96] ^ t[39];
  assign t[65] = t[97] & t[98];
  assign t[66] = t[99] ^ t[100];
  assign t[67] = t[101] ^ t[102];
  assign t[68] = t[8] ? t[103] : t[218];
  assign t[69] = t[87] ^ t[36];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[104] ^ t[20];
  assign t[71] = ~(t[105] ^ t[106]);
  assign t[72] = t[107] ^ t[99];
  assign t[73] = t[108] & t[109];
  assign t[74] = t[56] ^ t[68];
  assign t[75] = t[87] ^ t[110];
  assign t[76] = ~(t[78] & t[111]);
  assign t[77] = ~(t[219] ^ t[112]);
  assign t[78] = ~(t[113] & t[114]);
  assign t[79] = ~(t[48]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[220]);
  assign t[81] = t[21] ^ t[115];
  assign t[82] = t[116] ^ t[117];
  assign t[83] = t[118] ^ t[119];
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[215] ^ t[122];
  assign t[86] = t[216] ^ t[123];
  assign t[87] = t[124] ^ t[125];
  assign t[88] = t[8] ? t[126] : t[221];
  assign t[89] = t[27] ? t[127] : t[222];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] & t[129];
  assign t[91] = ~(t[90] ^ t[130]);
  assign t[92] = t[64] ^ t[131];
  assign t[93] = t[217] ^ t[132];
  assign t[94] = ~(t[133] ^ t[60]);
  assign t[95] = t[37] ^ t[98];
  assign t[96] = t[8] ? t[134] : t[223];
  assign t[97] = ~(t[59]);
  assign t[98] = t[210] ^ t[135];
  assign t[99] = t[136];
  assign t[9] = t[208] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [116:0] x;
 output y;

 wire [396:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~t[137];
  assign t[101] = t[138] ^ t[121];
  assign t[102] = t[139] & t[140];
  assign t[103] = t[218] ^ t[141];
  assign t[104] = t[142] ^ t[143];
  assign t[105] = t[42] ^ t[144];
  assign t[106] = t[145] ^ t[146];
  assign t[107] = ~t[147];
  assign t[108] = ~(t[72] ^ t[101]);
  assign t[109] = t[66] ^ t[148];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[149] & t[150];
  assign t[111] = ~(t[151] & t[152]);
  assign t[112] = t[153] ^ t[224];
  assign t[113] = ~(t[219]);
  assign t[114] = t[154] & t[153];
  assign t[115] = t[100] ^ t[155];
  assign t[116] = t[156] ^ t[157];
  assign t[117] = t[158] & t[159];
  assign t[118] = t[157] ^ t[145];
  assign t[119] = t[160] ^ t[161];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[107] ^ t[100];
  assign t[121] = t[162] & t[148];
  assign t[122] = t[163] ? x[56] : x[55];
  assign t[123] = t[163] ? x[58] : x[57];
  assign t[124] = t[164] & t[165];
  assign t[125] = t[166] & t[88];
  assign t[126] = t[221] ^ t[167];
  assign t[127] = t[222] ^ t[168];
  assign t[128] = ~(t[131]);
  assign t[129] = ~(t[96]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[37] ^ t[96];
  assign t[131] = t[98] ^ t[59];
  assign t[132] = t[79] ? x[60] : x[59];
  assign t[133] = t[96] ^ t[59];
  assign t[134] = t[223] ^ t[169];
  assign t[135] = t[8] ? t[170] : t[225];
  assign t[136] = t[27] ? t[171] : t[226];
  assign t[137] = t[27] ? t[172] : t[227];
  assign t[138] = t[173] & t[174];
  assign t[139] = ~(t[138] ^ t[175]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[120] ^ t[176];
  assign t[141] = t[163] ? x[71] : x[70];
  assign t[142] = t[156] ^ t[145];
  assign t[143] = t[177] & t[178];
  assign t[144] = t[133] ^ t[63];
  assign t[145] = t[179] ? t[180] : t[228];
  assign t[146] = t[160] ^ t[117];
  assign t[147] = t[27] ? t[181] : t[229];
  assign t[148] = t[182];
  assign t[149] = ~(t[124] ^ t[183]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[184] ^ t[185];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[186] | t[113]);
  assign t[153] = ~(t[230]);
  assign t[154] = ~(t[224]);
  assign t[155] = t[101] ^ t[73];
  assign t[156] = t[179] ? t[187] : t[231];
  assign t[157] = t[179] ? t[188] : t[232];
  assign t[158] = ~(t[116] ^ t[160]);
  assign t[159] = t[118] ^ t[178];
  assign t[15] = ~(t[27]);
  assign t[160] = t[189] ^ t[143];
  assign t[161] = t[190] & t[191];
  assign t[162] = ~(t[99]);
  assign t[163] = ~(t[49]);
  assign t[164] = ~(t[185]);
  assign t[165] = ~(t[55]);
  assign t[166] = ~(t[56]);
  assign t[167] = t[163] ? x[88] : x[87];
  assign t[168] = t[28] ? x[90] : x[89];
  assign t[169] = t[79] ? x[92] : x[91];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[225] ^ t[192];
  assign t[171] = t[226] ^ t[193];
  assign t[172] = t[227] ^ t[194];
  assign t[173] = ~(t[176]);
  assign t[174] = ~(t[107]);
  assign t[175] = t[66] ^ t[107];
  assign t[176] = t[148] ^ t[99];
  assign t[177] = ~(t[157]);
  assign t[178] = t[179] ? t[195] : t[233];
  assign t[179] = ~(t[15]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[228] ^ t[196];
  assign t[181] = t[229] ^ t[197];
  assign t[182] = t[27] ? t[198] : t[234];
  assign t[183] = t[74] ^ t[55];
  assign t[184] = t[55] ^ t[68];
  assign t[185] = t[88] ^ t[56];
  assign t[186] = ~(t[213]);
  assign t[187] = t[231] ^ t[199];
  assign t[188] = t[232] ^ t[200];
  assign t[189] = t[201] & t[202];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = ~(t[189] ^ t[203]);
  assign t[191] = t[142] ^ t[204];
  assign t[192] = t[28] ? x[100] : x[99];
  assign t[193] = t[28] ? x[102] : x[101];
  assign t[194] = t[79] ? x[104] : x[103];
  assign t[195] = t[233] ^ t[205];
  assign t[196] = t[206] ? x[106] : x[105];
  assign t[197] = t[79] ? x[108] : x[107];
  assign t[198] = t[234] ^ t[207];
  assign t[199] = t[206] ? x[110] : x[109];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[206] ? x[112] : x[111];
  assign t[201] = ~(t[204]);
  assign t[202] = ~(t[156]);
  assign t[203] = t[118] ^ t[156];
  assign t[204] = t[178] ^ t[157];
  assign t[205] = t[206] ? x[114] : x[113];
  assign t[206] = ~(t[49]);
  assign t[207] = t[163] ? x[116] : x[115];
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[39] ^ t[40];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = t[262] ^ x[4];
  assign t[236] = t[263] ^ x[9];
  assign t[237] = t[264] ^ x[12];
  assign t[238] = t[265] ^ x[15];
  assign t[239] = t[266] ^ x[18];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[21];
  assign t[241] = t[268] ^ x[24];
  assign t[242] = t[269] ^ x[27];
  assign t[243] = t[270] ^ x[30];
  assign t[244] = t[271] ^ x[33];
  assign t[245] = t[272] ^ x[36];
  assign t[246] = t[273] ^ x[39];
  assign t[247] = t[274] ^ x[42];
  assign t[248] = t[275] ^ x[45];
  assign t[249] = t[276] ^ x[48];
  assign t[24] = ~(t[33] ^ t[43]);
  assign t[250] = t[277] ^ x[51];
  assign t[251] = t[278] ^ x[54];
  assign t[252] = t[279] ^ x[63];
  assign t[253] = t[280] ^ x[66];
  assign t[254] = t[281] ^ x[69];
  assign t[255] = t[282] ^ x[74];
  assign t[256] = t[283] ^ x[77];
  assign t[257] = t[284] ^ x[80];
  assign t[258] = t[285] ^ x[83];
  assign t[259] = t[286] ^ x[86];
  assign t[25] = t[44] ^ t[45];
  assign t[260] = t[287] ^ x[95];
  assign t[261] = t[288] ^ x[98];
  assign t[262] = (t[289] & ~t[290]);
  assign t[263] = (t[291] & ~t[292]);
  assign t[264] = (t[293] & ~t[294]);
  assign t[265] = (t[295] & ~t[296]);
  assign t[266] = (t[297] & ~t[298]);
  assign t[267] = (t[299] & ~t[300]);
  assign t[268] = (t[301] & ~t[302]);
  assign t[269] = (t[303] & ~t[304]);
  assign t[26] = ~(t[46] ^ t[22]);
  assign t[270] = (t[305] & ~t[306]);
  assign t[271] = (t[307] & ~t[308]);
  assign t[272] = (t[309] & ~t[310]);
  assign t[273] = (t[311] & ~t[312]);
  assign t[274] = (t[313] & ~t[314]);
  assign t[275] = (t[315] & ~t[316]);
  assign t[276] = (t[317] & ~t[318]);
  assign t[277] = (t[319] & ~t[320]);
  assign t[278] = (t[321] & ~t[322]);
  assign t[279] = (t[323] & ~t[324]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[325] & ~t[326]);
  assign t[281] = (t[327] & ~t[328]);
  assign t[282] = (t[329] & ~t[330]);
  assign t[283] = (t[331] & ~t[332]);
  assign t[284] = (t[333] & ~t[334]);
  assign t[285] = (t[335] & ~t[336]);
  assign t[286] = (t[337] & ~t[338]);
  assign t[287] = (t[339] & ~t[340]);
  assign t[288] = (t[341] & ~t[342]);
  assign t[289] = t[343] ^ x[4];
  assign t[28] = ~(t[49]);
  assign t[290] = t[344] ^ x[3];
  assign t[291] = t[345] ^ x[9];
  assign t[292] = t[346] ^ x[8];
  assign t[293] = t[347] ^ x[12];
  assign t[294] = t[348] ^ x[11];
  assign t[295] = t[349] ^ x[15];
  assign t[296] = t[350] ^ x[14];
  assign t[297] = t[351] ^ x[18];
  assign t[298] = t[352] ^ x[17];
  assign t[299] = t[353] ^ x[21];
  assign t[29] = ~(t[209]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[20];
  assign t[301] = t[355] ^ x[24];
  assign t[302] = t[356] ^ x[23];
  assign t[303] = t[357] ^ x[27];
  assign t[304] = t[358] ^ x[26];
  assign t[305] = t[359] ^ x[30];
  assign t[306] = t[360] ^ x[29];
  assign t[307] = t[361] ^ x[33];
  assign t[308] = t[362] ^ x[32];
  assign t[309] = t[363] ^ x[36];
  assign t[30] = ~(t[210]);
  assign t[310] = t[364] ^ x[35];
  assign t[311] = t[365] ^ x[39];
  assign t[312] = t[366] ^ x[38];
  assign t[313] = t[367] ^ x[42];
  assign t[314] = t[368] ^ x[41];
  assign t[315] = t[369] ^ x[45];
  assign t[316] = t[370] ^ x[44];
  assign t[317] = t[371] ^ x[48];
  assign t[318] = t[372] ^ x[47];
  assign t[319] = t[373] ^ x[51];
  assign t[31] = ~(t[211]);
  assign t[320] = t[374] ^ x[50];
  assign t[321] = t[375] ^ x[54];
  assign t[322] = t[376] ^ x[53];
  assign t[323] = t[377] ^ x[63];
  assign t[324] = t[378] ^ x[62];
  assign t[325] = t[379] ^ x[66];
  assign t[326] = t[380] ^ x[65];
  assign t[327] = t[381] ^ x[69];
  assign t[328] = t[382] ^ x[68];
  assign t[329] = t[383] ^ x[74];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[73];
  assign t[331] = t[385] ^ x[77];
  assign t[332] = t[386] ^ x[76];
  assign t[333] = t[387] ^ x[80];
  assign t[334] = t[388] ^ x[79];
  assign t[335] = t[389] ^ x[83];
  assign t[336] = t[390] ^ x[82];
  assign t[337] = t[391] ^ x[86];
  assign t[338] = t[392] ^ x[85];
  assign t[339] = t[393] ^ x[95];
  assign t[33] = ~(t[52] ^ t[46]);
  assign t[340] = t[394] ^ x[94];
  assign t[341] = t[395] ^ x[98];
  assign t[342] = t[396] ^ x[97];
  assign t[343] = (x[2]);
  assign t[344] = (x[2]);
  assign t[345] = (x[7]);
  assign t[346] = (x[7]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[49]);
  assign t[374] = (x[49]);
  assign t[375] = (x[52]);
  assign t[376] = (x[52]);
  assign t[377] = (x[61]);
  assign t[378] = (x[61]);
  assign t[379] = (x[64]);
  assign t[37] = t[59] ^ t[39];
  assign t[380] = (x[64]);
  assign t[381] = (x[67]);
  assign t[382] = (x[67]);
  assign t[383] = (x[72]);
  assign t[384] = (x[72]);
  assign t[385] = (x[75]);
  assign t[386] = (x[75]);
  assign t[387] = (x[78]);
  assign t[388] = (x[78]);
  assign t[389] = (x[81]);
  assign t[38] = t[60] ^ t[61];
  assign t[390] = (x[81]);
  assign t[391] = (x[84]);
  assign t[392] = (x[84]);
  assign t[393] = (x[93]);
  assign t[394] = (x[93]);
  assign t[395] = (x[96]);
  assign t[396] = (x[96]);
  assign t[39] = t[212] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[60] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66] ^ t[67];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = ~(t[70] ^ t[71]);
  assign t[45] = t[72] ^ t[73];
  assign t[46] = t[74] ^ t[75];
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = t[213] | t[78];
  assign t[49] = ~(t[79]);
  assign t[4] = t[8] ? t[9] : t[208];
  assign t[50] = ~(t[214]);
  assign t[51] = ~(t[80] & t[212]);
  assign t[52] = ~(t[81] ^ t[82]);
  assign t[53] = t[83] ^ t[84];
  assign t[54] = ~(t[43] ^ t[22]);
  assign t[55] = t[8] ? t[85] : t[215];
  assign t[56] = t[8] ? t[86] : t[216];
  assign t[57] = ~(t[35] ^ t[87]);
  assign t[58] = t[74] ^ t[88];
  assign t[59] = t[209] ^ t[89];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[65];
  assign t[61] = t[91] & t[92];
  assign t[62] = t[8] ? t[93] : t[217];
  assign t[63] = t[94] & t[95];
  assign t[64] = t[96] ^ t[39];
  assign t[65] = t[97] & t[98];
  assign t[66] = t[99] ^ t[100];
  assign t[67] = t[101] ^ t[102];
  assign t[68] = t[8] ? t[103] : t[218];
  assign t[69] = t[87] ^ t[36];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[104] ^ t[20];
  assign t[71] = ~(t[105] ^ t[106]);
  assign t[72] = t[107] ^ t[99];
  assign t[73] = t[108] & t[109];
  assign t[74] = t[56] ^ t[68];
  assign t[75] = t[87] ^ t[110];
  assign t[76] = ~(t[78] & t[111]);
  assign t[77] = ~(t[219] ^ t[112]);
  assign t[78] = ~(t[113] & t[114]);
  assign t[79] = ~(t[48]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[220]);
  assign t[81] = t[21] ^ t[115];
  assign t[82] = t[116] ^ t[117];
  assign t[83] = t[118] ^ t[119];
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[215] ^ t[122];
  assign t[86] = t[216] ^ t[123];
  assign t[87] = t[124] ^ t[125];
  assign t[88] = t[8] ? t[126] : t[221];
  assign t[89] = t[27] ? t[127] : t[222];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] & t[129];
  assign t[91] = ~(t[90] ^ t[130]);
  assign t[92] = t[64] ^ t[131];
  assign t[93] = t[217] ^ t[132];
  assign t[94] = ~(t[133] ^ t[60]);
  assign t[95] = t[37] ^ t[98];
  assign t[96] = t[8] ? t[134] : t[223];
  assign t[97] = ~(t[59]);
  assign t[98] = t[210] ^ t[135];
  assign t[99] = t[136];
  assign t[9] = t[208] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind116(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[133] & t[134];
  assign t[101] = ~(t[99] ^ t[135]);
  assign t[102] = t[136] ^ t[137];
  assign t[103] = t[208] ^ t[138];
  assign t[104] = t[139] & t[140];
  assign t[105] = t[141] & t[126];
  assign t[106] = t[142] & t[143];
  assign t[107] = t[8] ? t[144] : t[212];
  assign t[108] = t[198] ^ t[145];
  assign t[109] = ~(t[70] ^ t[146]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[147] ^ t[148];
  assign t[111] = t[147] ^ t[149];
  assign t[112] = t[150] ^ t[63];
  assign t[113] = t[91] ^ t[41];
  assign t[114] = t[35] ^ t[151];
  assign t[115] = t[205] ^ t[152];
  assign t[116] = t[146] ^ t[71];
  assign t[117] = ~(t[153] & t[154]);
  assign t[118] = t[155] ^ t[213];
  assign t[119] = ~(t[209]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[156] & t[155];
  assign t[121] = ~(t[50]);
  assign t[122] = t[8] ? t[157] : t[214];
  assign t[123] = t[211] ^ t[158];
  assign t[124] = t[27] ? t[159] : t[215];
  assign t[125] = t[27] ? t[160] : t[216];
  assign t[126] = t[161];
  assign t[127] = t[162] ? x[69] : x[68];
  assign t[128] = ~(t[112] ^ t[64]);
  assign t[129] = t[39] ^ t[134];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[162] ? x[71] : x[70];
  assign t[131] = ~(t[137]);
  assign t[132] = ~(t[150]);
  assign t[133] = ~(t[63]);
  assign t[134] = t[95] ? t[163] : t[217];
  assign t[135] = t[39] ^ t[150];
  assign t[136] = t[150] ^ t[61];
  assign t[137] = t[134] ^ t[63];
  assign t[138] = t[80] ? x[76] : x[75];
  assign t[139] = ~(t[164]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = ~(t[91]);
  assign t[141] = ~(t[92]);
  assign t[142] = ~(t[104] ^ t[165]);
  assign t[143] = t[113] ^ t[164];
  assign t[144] = t[212] ^ t[166];
  assign t[145] = t[27] ? t[167] : t[218];
  assign t[146] = t[168] ^ t[169];
  assign t[147] = t[108] ^ t[115];
  assign t[148] = t[199] ^ t[170];
  assign t[149] = t[146] ^ t[171];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[95] ? t[172] : t[219];
  assign t[151] = t[173] & t[174];
  assign t[152] = t[8] ? t[175] : t[220];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[176] | t[119]);
  assign t[155] = ~(t[221]);
  assign t[156] = ~(t[213]);
  assign t[157] = t[214] ^ t[177];
  assign t[158] = t[121] ? x[90] : x[89];
  assign t[159] = t[215] ^ t[178];
  assign t[15] = ~(t[27]);
  assign t[160] = t[216] ^ t[179];
  assign t[161] = t[27] ? t[180] : t[222];
  assign t[162] = ~(t[50]);
  assign t[163] = t[217] ^ t[181];
  assign t[164] = t[126] ^ t[92];
  assign t[165] = t[68] ^ t[91];
  assign t[166] = t[80] ? x[95] : x[94];
  assign t[167] = t[218] ^ t[182];
  assign t[168] = t[183] & t[184];
  assign t[169] = t[185] & t[148];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[8] ? t[186] : t[223];
  assign t[171] = t[187] & t[188];
  assign t[172] = t[219] ^ t[189];
  assign t[173] = ~(t[190] ^ t[35]);
  assign t[174] = t[19] ^ t[87];
  assign t[175] = t[220] ^ t[191];
  assign t[176] = ~(t[203]);
  assign t[177] = t[121] ? x[100] : x[99];
  assign t[178] = t[80] ? x[102] : x[101];
  assign t[179] = t[28] ? x[104] : x[103];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[222] ^ t[192];
  assign t[181] = t[162] ? x[106] : x[105];
  assign t[182] = t[28] ? x[108] : x[107];
  assign t[183] = ~(t[193]);
  assign t[184] = ~(t[107]);
  assign t[185] = ~(t[108]);
  assign t[186] = t[223] ^ t[194];
  assign t[187] = ~(t[168] ^ t[195]);
  assign t[188] = t[196] ^ t[193];
  assign t[189] = t[162] ? x[110] : x[109];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[122] ^ t[33];
  assign t[191] = t[80] ? x[112] : x[111];
  assign t[192] = t[121] ? x[114] : x[113];
  assign t[193] = t[148] ^ t[108];
  assign t[194] = t[28] ? x[116] : x[115];
  assign t[195] = t[147] ^ t[107];
  assign t[196] = t[107] ^ t[115];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = t[39] ^ t[40];
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[36];
  assign t[235] = t[262] ^ x[39];
  assign t[236] = t[263] ^ x[42];
  assign t[237] = t[264] ^ x[45];
  assign t[238] = t[265] ^ x[52];
  assign t[239] = t[266] ^ x[55];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[58];
  assign t[241] = t[268] ^ x[61];
  assign t[242] = t[269] ^ x[64];
  assign t[243] = t[270] ^ x[67];
  assign t[244] = t[271] ^ x[74];
  assign t[245] = t[272] ^ x[79];
  assign t[246] = t[273] ^ x[82];
  assign t[247] = t[274] ^ x[85];
  assign t[248] = t[275] ^ x[88];
  assign t[249] = t[276] ^ x[93];
  assign t[24] = t[43] ^ t[44];
  assign t[250] = t[277] ^ x[98];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = ~(t[45] ^ t[11]);
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[36];
  assign t[299] = t[353] ^ x[35];
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[39];
  assign t[301] = t[355] ^ x[38];
  assign t[302] = t[356] ^ x[42];
  assign t[303] = t[357] ^ x[41];
  assign t[304] = t[358] ^ x[45];
  assign t[305] = t[359] ^ x[44];
  assign t[306] = t[360] ^ x[52];
  assign t[307] = t[361] ^ x[51];
  assign t[308] = t[362] ^ x[55];
  assign t[309] = t[363] ^ x[54];
  assign t[30] = ~(t[199]);
  assign t[310] = t[364] ^ x[58];
  assign t[311] = t[365] ^ x[57];
  assign t[312] = t[366] ^ x[61];
  assign t[313] = t[367] ^ x[60];
  assign t[314] = t[368] ^ x[64];
  assign t[315] = t[369] ^ x[63];
  assign t[316] = t[370] ^ x[67];
  assign t[317] = t[371] ^ x[66];
  assign t[318] = t[372] ^ x[74];
  assign t[319] = t[373] ^ x[73];
  assign t[31] = ~(t[200]);
  assign t[320] = t[374] ^ x[79];
  assign t[321] = t[375] ^ x[78];
  assign t[322] = t[376] ^ x[82];
  assign t[323] = t[377] ^ x[81];
  assign t[324] = t[378] ^ x[85];
  assign t[325] = t[379] ^ x[84];
  assign t[326] = t[380] ^ x[88];
  assign t[327] = t[381] ^ x[87];
  assign t[328] = t[382] ^ x[93];
  assign t[329] = t[383] ^ x[92];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[384] ^ x[98];
  assign t[331] = t[385] ^ x[97];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = t[8] ? t[53] : t[201];
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = t[8] ? t[54] : t[202];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[34]);
  assign t[353] = (x[34]);
  assign t[354] = (x[37]);
  assign t[355] = (x[37]);
  assign t[356] = (x[40]);
  assign t[357] = (x[40]);
  assign t[358] = (x[43]);
  assign t[359] = (x[43]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[50]);
  assign t[361] = (x[50]);
  assign t[362] = (x[53]);
  assign t[363] = (x[53]);
  assign t[364] = (x[56]);
  assign t[365] = (x[56]);
  assign t[366] = (x[59]);
  assign t[367] = (x[59]);
  assign t[368] = (x[62]);
  assign t[369] = (x[62]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[65]);
  assign t[371] = (x[65]);
  assign t[372] = (x[72]);
  assign t[373] = (x[72]);
  assign t[374] = (x[77]);
  assign t[375] = (x[77]);
  assign t[376] = (x[80]);
  assign t[377] = (x[80]);
  assign t[378] = (x[83]);
  assign t[379] = (x[83]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[86]);
  assign t[381] = (x[86]);
  assign t[382] = (x[91]);
  assign t[383] = (x[91]);
  assign t[384] = (x[96]);
  assign t[385] = (x[96]);
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = ~t[66];
  assign t[42] = t[67] ^ t[60];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = ~(t[72] ^ t[73]);
  assign t[46] = t[22] ^ t[74];
  assign t[47] = ~(t[75] ^ t[76]);
  assign t[48] = ~(t[77] & t[78]);
  assign t[49] = t[203] | t[79];
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[80]);
  assign t[51] = ~(t[204]);
  assign t[52] = ~(t[81] & t[205]);
  assign t[53] = t[201] ^ t[82];
  assign t[54] = t[202] ^ t[83];
  assign t[55] = t[84] & t[85];
  assign t[56] = t[86] & t[87];
  assign t[57] = ~(t[55] ^ t[88]);
  assign t[58] = t[89] ^ t[90];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] & t[94];
  assign t[61] = t[95] ? t[96] : t[206];
  assign t[62] = t[64] ^ t[97];
  assign t[63] = t[95] ? t[98] : t[207];
  assign t[64] = t[99] ^ t[100];
  assign t[65] = t[101] & t[102];
  assign t[66] = t[27] ? t[103] : t[208];
  assign t[67] = t[104] ^ t[105];
  assign t[68] = t[92] ^ t[41];
  assign t[69] = t[67] ^ t[106];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[107] ^ t[108];
  assign t[71] = t[109] & t[110];
  assign t[72] = t[111] ^ t[23];
  assign t[73] = t[112] ^ t[97];
  assign t[74] = t[113] ^ t[105];
  assign t[75] = t[34] ^ t[114];
  assign t[76] = t[115] ^ t[116];
  assign t[77] = ~(t[79] & t[117]);
  assign t[78] = ~(t[209] ^ t[118]);
  assign t[79] = ~(t[119] & t[120]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[49]);
  assign t[81] = ~(t[210]);
  assign t[82] = t[121] ? x[47] : x[46];
  assign t[83] = t[121] ? x[49] : x[48];
  assign t[84] = ~(t[90]);
  assign t[85] = ~(t[122]);
  assign t[86] = ~(t[33]);
  assign t[87] = t[8] ? t[123] : t[211];
  assign t[88] = t[19] ^ t[122];
  assign t[89] = t[122] ^ t[34];
  assign t[8] = ~(t[15]);
  assign t[90] = t[87] ^ t[33];
  assign t[91] = ~t[124];
  assign t[92] = t[125];
  assign t[93] = ~(t[59] ^ t[67]);
  assign t[94] = t[68] ^ t[126];
  assign t[95] = ~(t[15]);
  assign t[96] = t[206] ^ t[127];
  assign t[97] = t[128] & t[129];
  assign t[98] = t[207] ^ t[130];
  assign t[99] = t[131] & t[132];
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [116:0] x;
 output y;

 wire [385:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[133] & t[134];
  assign t[101] = ~(t[99] ^ t[135]);
  assign t[102] = t[136] ^ t[137];
  assign t[103] = t[208] ^ t[138];
  assign t[104] = t[139] & t[140];
  assign t[105] = t[141] & t[126];
  assign t[106] = t[142] & t[143];
  assign t[107] = t[8] ? t[144] : t[212];
  assign t[108] = t[198] ^ t[145];
  assign t[109] = ~(t[70] ^ t[146]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[147] ^ t[148];
  assign t[111] = t[147] ^ t[149];
  assign t[112] = t[150] ^ t[63];
  assign t[113] = t[91] ^ t[41];
  assign t[114] = t[35] ^ t[151];
  assign t[115] = t[205] ^ t[152];
  assign t[116] = t[146] ^ t[71];
  assign t[117] = ~(t[153] & t[154]);
  assign t[118] = t[155] ^ t[213];
  assign t[119] = ~(t[209]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[156] & t[155];
  assign t[121] = ~(t[50]);
  assign t[122] = t[8] ? t[157] : t[214];
  assign t[123] = t[211] ^ t[158];
  assign t[124] = t[27] ? t[159] : t[215];
  assign t[125] = t[27] ? t[160] : t[216];
  assign t[126] = t[161];
  assign t[127] = t[162] ? x[69] : x[68];
  assign t[128] = ~(t[112] ^ t[64]);
  assign t[129] = t[39] ^ t[134];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[162] ? x[71] : x[70];
  assign t[131] = ~(t[137]);
  assign t[132] = ~(t[150]);
  assign t[133] = ~(t[63]);
  assign t[134] = t[95] ? t[163] : t[217];
  assign t[135] = t[39] ^ t[150];
  assign t[136] = t[150] ^ t[61];
  assign t[137] = t[134] ^ t[63];
  assign t[138] = t[80] ? x[76] : x[75];
  assign t[139] = ~(t[164]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = ~(t[91]);
  assign t[141] = ~(t[92]);
  assign t[142] = ~(t[104] ^ t[165]);
  assign t[143] = t[113] ^ t[164];
  assign t[144] = t[212] ^ t[166];
  assign t[145] = t[27] ? t[167] : t[218];
  assign t[146] = t[168] ^ t[169];
  assign t[147] = t[108] ^ t[115];
  assign t[148] = t[199] ^ t[170];
  assign t[149] = t[146] ^ t[171];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[95] ? t[172] : t[219];
  assign t[151] = t[173] & t[174];
  assign t[152] = t[8] ? t[175] : t[220];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[176] | t[119]);
  assign t[155] = ~(t[221]);
  assign t[156] = ~(t[213]);
  assign t[157] = t[214] ^ t[177];
  assign t[158] = t[121] ? x[90] : x[89];
  assign t[159] = t[215] ^ t[178];
  assign t[15] = ~(t[27]);
  assign t[160] = t[216] ^ t[179];
  assign t[161] = t[27] ? t[180] : t[222];
  assign t[162] = ~(t[50]);
  assign t[163] = t[217] ^ t[181];
  assign t[164] = t[126] ^ t[92];
  assign t[165] = t[68] ^ t[91];
  assign t[166] = t[80] ? x[95] : x[94];
  assign t[167] = t[218] ^ t[182];
  assign t[168] = t[183] & t[184];
  assign t[169] = t[185] & t[148];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[8] ? t[186] : t[223];
  assign t[171] = t[187] & t[188];
  assign t[172] = t[219] ^ t[189];
  assign t[173] = ~(t[190] ^ t[35]);
  assign t[174] = t[19] ^ t[87];
  assign t[175] = t[220] ^ t[191];
  assign t[176] = ~(t[203]);
  assign t[177] = t[121] ? x[100] : x[99];
  assign t[178] = t[80] ? x[102] : x[101];
  assign t[179] = t[28] ? x[104] : x[103];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[222] ^ t[192];
  assign t[181] = t[162] ? x[106] : x[105];
  assign t[182] = t[28] ? x[108] : x[107];
  assign t[183] = ~(t[193]);
  assign t[184] = ~(t[107]);
  assign t[185] = ~(t[108]);
  assign t[186] = t[223] ^ t[194];
  assign t[187] = ~(t[168] ^ t[195]);
  assign t[188] = t[196] ^ t[193];
  assign t[189] = t[162] ? x[110] : x[109];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[122] ^ t[33];
  assign t[191] = t[80] ? x[112] : x[111];
  assign t[192] = t[121] ? x[114] : x[113];
  assign t[193] = t[148] ^ t[108];
  assign t[194] = t[28] ? x[116] : x[115];
  assign t[195] = t[147] ^ t[107];
  assign t[196] = t[107] ^ t[115];
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[35] ^ t[36];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[38]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = t[251] ^ x[4];
  assign t[225] = t[252] ^ x[9];
  assign t[226] = t[253] ^ x[12];
  assign t[227] = t[254] ^ x[15];
  assign t[228] = t[255] ^ x[18];
  assign t[229] = t[256] ^ x[21];
  assign t[22] = t[39] ^ t[40];
  assign t[230] = t[257] ^ x[24];
  assign t[231] = t[258] ^ x[27];
  assign t[232] = t[259] ^ x[30];
  assign t[233] = t[260] ^ x[33];
  assign t[234] = t[261] ^ x[36];
  assign t[235] = t[262] ^ x[39];
  assign t[236] = t[263] ^ x[42];
  assign t[237] = t[264] ^ x[45];
  assign t[238] = t[265] ^ x[52];
  assign t[239] = t[266] ^ x[55];
  assign t[23] = t[41] ^ t[42];
  assign t[240] = t[267] ^ x[58];
  assign t[241] = t[268] ^ x[61];
  assign t[242] = t[269] ^ x[64];
  assign t[243] = t[270] ^ x[67];
  assign t[244] = t[271] ^ x[74];
  assign t[245] = t[272] ^ x[79];
  assign t[246] = t[273] ^ x[82];
  assign t[247] = t[274] ^ x[85];
  assign t[248] = t[275] ^ x[88];
  assign t[249] = t[276] ^ x[93];
  assign t[24] = t[43] ^ t[44];
  assign t[250] = t[277] ^ x[98];
  assign t[251] = (t[278] & ~t[279]);
  assign t[252] = (t[280] & ~t[281]);
  assign t[253] = (t[282] & ~t[283]);
  assign t[254] = (t[284] & ~t[285]);
  assign t[255] = (t[286] & ~t[287]);
  assign t[256] = (t[288] & ~t[289]);
  assign t[257] = (t[290] & ~t[291]);
  assign t[258] = (t[292] & ~t[293]);
  assign t[259] = (t[294] & ~t[295]);
  assign t[25] = ~(t[45] ^ t[11]);
  assign t[260] = (t[296] & ~t[297]);
  assign t[261] = (t[298] & ~t[299]);
  assign t[262] = (t[300] & ~t[301]);
  assign t[263] = (t[302] & ~t[303]);
  assign t[264] = (t[304] & ~t[305]);
  assign t[265] = (t[306] & ~t[307]);
  assign t[266] = (t[308] & ~t[309]);
  assign t[267] = (t[310] & ~t[311]);
  assign t[268] = (t[312] & ~t[313]);
  assign t[269] = (t[314] & ~t[315]);
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[270] = (t[316] & ~t[317]);
  assign t[271] = (t[318] & ~t[319]);
  assign t[272] = (t[320] & ~t[321]);
  assign t[273] = (t[322] & ~t[323]);
  assign t[274] = (t[324] & ~t[325]);
  assign t[275] = (t[326] & ~t[327]);
  assign t[276] = (t[328] & ~t[329]);
  assign t[277] = (t[330] & ~t[331]);
  assign t[278] = t[332] ^ x[4];
  assign t[279] = t[333] ^ x[3];
  assign t[27] = ~(t[48] & t[49]);
  assign t[280] = t[334] ^ x[9];
  assign t[281] = t[335] ^ x[8];
  assign t[282] = t[336] ^ x[12];
  assign t[283] = t[337] ^ x[11];
  assign t[284] = t[338] ^ x[15];
  assign t[285] = t[339] ^ x[14];
  assign t[286] = t[340] ^ x[18];
  assign t[287] = t[341] ^ x[17];
  assign t[288] = t[342] ^ x[21];
  assign t[289] = t[343] ^ x[20];
  assign t[28] = ~(t[50]);
  assign t[290] = t[344] ^ x[24];
  assign t[291] = t[345] ^ x[23];
  assign t[292] = t[346] ^ x[27];
  assign t[293] = t[347] ^ x[26];
  assign t[294] = t[348] ^ x[30];
  assign t[295] = t[349] ^ x[29];
  assign t[296] = t[350] ^ x[33];
  assign t[297] = t[351] ^ x[32];
  assign t[298] = t[352] ^ x[36];
  assign t[299] = t[353] ^ x[35];
  assign t[29] = ~(t[198]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[39];
  assign t[301] = t[355] ^ x[38];
  assign t[302] = t[356] ^ x[42];
  assign t[303] = t[357] ^ x[41];
  assign t[304] = t[358] ^ x[45];
  assign t[305] = t[359] ^ x[44];
  assign t[306] = t[360] ^ x[52];
  assign t[307] = t[361] ^ x[51];
  assign t[308] = t[362] ^ x[55];
  assign t[309] = t[363] ^ x[54];
  assign t[30] = ~(t[199]);
  assign t[310] = t[364] ^ x[58];
  assign t[311] = t[365] ^ x[57];
  assign t[312] = t[366] ^ x[61];
  assign t[313] = t[367] ^ x[60];
  assign t[314] = t[368] ^ x[64];
  assign t[315] = t[369] ^ x[63];
  assign t[316] = t[370] ^ x[67];
  assign t[317] = t[371] ^ x[66];
  assign t[318] = t[372] ^ x[74];
  assign t[319] = t[373] ^ x[73];
  assign t[31] = ~(t[200]);
  assign t[320] = t[374] ^ x[79];
  assign t[321] = t[375] ^ x[78];
  assign t[322] = t[376] ^ x[82];
  assign t[323] = t[377] ^ x[81];
  assign t[324] = t[378] ^ x[85];
  assign t[325] = t[379] ^ x[84];
  assign t[326] = t[380] ^ x[88];
  assign t[327] = t[381] ^ x[87];
  assign t[328] = t[382] ^ x[93];
  assign t[329] = t[383] ^ x[92];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[384] ^ x[98];
  assign t[331] = t[385] ^ x[97];
  assign t[332] = (x[2]);
  assign t[333] = (x[2]);
  assign t[334] = (x[7]);
  assign t[335] = (x[7]);
  assign t[336] = (x[10]);
  assign t[337] = (x[10]);
  assign t[338] = (x[13]);
  assign t[339] = (x[13]);
  assign t[33] = t[8] ? t[53] : t[201];
  assign t[340] = (x[16]);
  assign t[341] = (x[16]);
  assign t[342] = (x[19]);
  assign t[343] = (x[19]);
  assign t[344] = (x[22]);
  assign t[345] = (x[22]);
  assign t[346] = (x[25]);
  assign t[347] = (x[25]);
  assign t[348] = (x[28]);
  assign t[349] = (x[28]);
  assign t[34] = t[8] ? t[54] : t[202];
  assign t[350] = (x[31]);
  assign t[351] = (x[31]);
  assign t[352] = (x[34]);
  assign t[353] = (x[34]);
  assign t[354] = (x[37]);
  assign t[355] = (x[37]);
  assign t[356] = (x[40]);
  assign t[357] = (x[40]);
  assign t[358] = (x[43]);
  assign t[359] = (x[43]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[50]);
  assign t[361] = (x[50]);
  assign t[362] = (x[53]);
  assign t[363] = (x[53]);
  assign t[364] = (x[56]);
  assign t[365] = (x[56]);
  assign t[366] = (x[59]);
  assign t[367] = (x[59]);
  assign t[368] = (x[62]);
  assign t[369] = (x[62]);
  assign t[36] = t[57] & t[58];
  assign t[370] = (x[65]);
  assign t[371] = (x[65]);
  assign t[372] = (x[72]);
  assign t[373] = (x[72]);
  assign t[374] = (x[77]);
  assign t[375] = (x[77]);
  assign t[376] = (x[80]);
  assign t[377] = (x[80]);
  assign t[378] = (x[83]);
  assign t[379] = (x[83]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[86]);
  assign t[381] = (x[86]);
  assign t[382] = (x[91]);
  assign t[383] = (x[91]);
  assign t[384] = (x[96]);
  assign t[385] = (x[96]);
  assign t[38] = t[61] ^ t[62];
  assign t[39] = t[63] ^ t[61];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[64] ^ t[65];
  assign t[41] = ~t[66];
  assign t[42] = t[67] ^ t[60];
  assign t[43] = t[68] ^ t[69];
  assign t[44] = t[70] ^ t[71];
  assign t[45] = ~(t[72] ^ t[73]);
  assign t[46] = t[22] ^ t[74];
  assign t[47] = ~(t[75] ^ t[76]);
  assign t[48] = ~(t[77] & t[78]);
  assign t[49] = t[203] | t[79];
  assign t[4] = t[8] ? t[9] : t[197];
  assign t[50] = ~(t[80]);
  assign t[51] = ~(t[204]);
  assign t[52] = ~(t[81] & t[205]);
  assign t[53] = t[201] ^ t[82];
  assign t[54] = t[202] ^ t[83];
  assign t[55] = t[84] & t[85];
  assign t[56] = t[86] & t[87];
  assign t[57] = ~(t[55] ^ t[88]);
  assign t[58] = t[89] ^ t[90];
  assign t[59] = t[91] ^ t[92];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] & t[94];
  assign t[61] = t[95] ? t[96] : t[206];
  assign t[62] = t[64] ^ t[97];
  assign t[63] = t[95] ? t[98] : t[207];
  assign t[64] = t[99] ^ t[100];
  assign t[65] = t[101] & t[102];
  assign t[66] = t[27] ? t[103] : t[208];
  assign t[67] = t[104] ^ t[105];
  assign t[68] = t[92] ^ t[41];
  assign t[69] = t[67] ^ t[106];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[107] ^ t[108];
  assign t[71] = t[109] & t[110];
  assign t[72] = t[111] ^ t[23];
  assign t[73] = t[112] ^ t[97];
  assign t[74] = t[113] ^ t[105];
  assign t[75] = t[34] ^ t[114];
  assign t[76] = t[115] ^ t[116];
  assign t[77] = ~(t[79] & t[117]);
  assign t[78] = ~(t[209] ^ t[118]);
  assign t[79] = ~(t[119] & t[120]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[49]);
  assign t[81] = ~(t[210]);
  assign t[82] = t[121] ? x[47] : x[46];
  assign t[83] = t[121] ? x[49] : x[48];
  assign t[84] = ~(t[90]);
  assign t[85] = ~(t[122]);
  assign t[86] = ~(t[33]);
  assign t[87] = t[8] ? t[123] : t[211];
  assign t[88] = t[19] ^ t[122];
  assign t[89] = t[122] ^ t[34];
  assign t[8] = ~(t[15]);
  assign t[90] = t[87] ^ t[33];
  assign t[91] = ~t[124];
  assign t[92] = t[125];
  assign t[93] = ~(t[59] ^ t[67]);
  assign t[94] = t[68] ^ t[126];
  assign t[95] = ~(t[15]);
  assign t[96] = t[206] ^ t[127];
  assign t[97] = t[128] & t[129];
  assign t[98] = t[207] ^ t[130];
  assign t[99] = t[131] & t[132];
  assign t[9] = t[197] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [116:0] x;
 output y;

 wire [383:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[87]);
  assign t[101] = ~(t[88]);
  assign t[102] = t[9] ? t[137] : t[212];
  assign t[103] = t[88] ^ t[27];
  assign t[104] = t[76] ? x[61] : x[60];
  assign t[105] = t[206] ^ t[138];
  assign t[106] = t[139] & t[140];
  assign t[107] = t[141] & t[72];
  assign t[108] = t[200] ^ t[142];
  assign t[109] = t[9] ? t[143] : t[213];
  assign t[10] = t[195] ^ t[20];
  assign t[110] = ~(t[144] & t[145]);
  assign t[111] = t[146] ^ t[214];
  assign t[112] = ~(t[207]);
  assign t[113] = t[147] & t[146];
  assign t[114] = t[148] ^ t[65];
  assign t[115] = ~(t[149] ^ t[40]);
  assign t[116] = t[150] ^ t[151];
  assign t[117] = t[44] ^ t[108];
  assign t[118] = t[70] ^ t[30];
  assign t[119] = t[31] ? t[152] : t[215];
  assign t[11] = ~(t[196]);
  assign t[120] = t[31] ? t[153] : t[216];
  assign t[121] = t[154];
  assign t[122] = t[31] ? t[155] : t[217];
  assign t[123] = t[156] & t[157];
  assign t[124] = t[158] ^ t[54];
  assign t[125] = t[159] & t[160];
  assign t[126] = t[208] ^ t[161];
  assign t[127] = t[209] ^ t[162];
  assign t[128] = t[210] ^ t[163];
  assign t[129] = t[94] ? t[164] : t[218];
  assign t[12] = ~(t[197]);
  assign t[130] = t[211] ^ t[165];
  assign t[131] = t[166] & t[167];
  assign t[132] = t[168] ? x[81] : x[80];
  assign t[133] = t[169] & t[170];
  assign t[134] = ~(t[171] ^ t[96]);
  assign t[135] = t[150] ^ t[91];
  assign t[136] = t[102] ^ t[88];
  assign t[137] = t[212] ^ t[172];
  assign t[138] = t[32] ? x[83] : x[82];
  assign t[139] = ~(t[173]);
  assign t[13] = ~(t[198]);
  assign t[140] = ~(t[44]);
  assign t[141] = ~(t[45]);
  assign t[142] = t[9] ? t[174] : t[219];
  assign t[143] = t[213] ^ t[175];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[176] | t[112]);
  assign t[146] = ~(t[220]);
  assign t[147] = ~(t[214]);
  assign t[148] = t[87] ^ t[27];
  assign t[149] = t[177] ^ t[125];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = t[129] ^ t[61];
  assign t[151] = t[96] ^ t[178];
  assign t[152] = t[215] ^ t[179];
  assign t[153] = t[216] ^ t[180];
  assign t[154] = t[31] ? t[181] : t[221];
  assign t[155] = t[217] ^ t[182];
  assign t[156] = ~(t[106] ^ t[183]);
  assign t[157] = t[117] ^ t[173];
  assign t[158] = t[184] & t[185];
  assign t[159] = ~(t[177] ^ t[124]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[92] ^ t[84];
  assign t[161] = t[98] ? x[94] : x[93];
  assign t[162] = t[98] ? x[96] : x[95];
  assign t[163] = t[168] ? x[98] : x[97];
  assign t[164] = t[218] ^ t[186];
  assign t[165] = t[168] ? x[100] : x[99];
  assign t[166] = ~(t[158] ^ t[187]);
  assign t[167] = t[53] ^ t[188];
  assign t[168] = ~(t[50]);
  assign t[169] = ~(t[189]);
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = ~(t[89]);
  assign t[171] = t[89] ^ t[129];
  assign t[172] = t[98] ? x[102] : x[101];
  assign t[173] = t[72] ^ t[45];
  assign t[174] = t[219] ^ t[190];
  assign t[175] = t[32] ? x[104] : x[103];
  assign t[176] = ~(t[204]);
  assign t[177] = t[81] ^ t[121];
  assign t[178] = t[191] & t[192];
  assign t[179] = t[76] ? x[106] : x[105];
  assign t[17] = t[27] ^ t[28];
  assign t[180] = t[76] ? x[108] : x[107];
  assign t[181] = t[221] ^ t[193];
  assign t[182] = t[98] ? x[110] : x[109];
  assign t[183] = t[71] ^ t[44];
  assign t[184] = ~(t[188]);
  assign t[185] = ~(t[81]);
  assign t[186] = t[168] ? x[112] : x[111];
  assign t[187] = t[92] ^ t[81];
  assign t[188] = t[84] ^ t[121];
  assign t[189] = t[91] ^ t[129];
  assign t[18] = t[29] ^ t[30];
  assign t[190] = t[76] ? x[114] : x[113];
  assign t[191] = ~(t[133] ^ t[194]);
  assign t[192] = t[58] ^ t[189];
  assign t[193] = t[32] ? x[116] : x[115];
  assign t[194] = t[150] ^ t[89];
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[199]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = t[249] ^ x[4];
  assign t[223] = t[250] ^ x[7];
  assign t[224] = t[251] ^ x[10];
  assign t[225] = t[252] ^ x[13];
  assign t[226] = t[253] ^ x[18];
  assign t[227] = t[254] ^ x[21];
  assign t[228] = t[255] ^ x[24];
  assign t[229] = t[256] ^ x[27];
  assign t[22] = ~(t[33] & t[200]);
  assign t[230] = t[257] ^ x[30];
  assign t[231] = t[258] ^ x[33];
  assign t[232] = t[259] ^ x[36];
  assign t[233] = t[260] ^ x[41];
  assign t[234] = t[261] ^ x[44];
  assign t[235] = t[262] ^ x[47];
  assign t[236] = t[263] ^ x[50];
  assign t[237] = t[264] ^ x[53];
  assign t[238] = t[265] ^ x[56];
  assign t[239] = t[266] ^ x[59];
  assign t[23] = t[34] ^ t[35];
  assign t[240] = t[267] ^ x[64];
  assign t[241] = t[268] ^ x[67];
  assign t[242] = t[269] ^ x[70];
  assign t[243] = t[270] ^ x[73];
  assign t[244] = t[271] ^ x[76];
  assign t[245] = t[272] ^ x[79];
  assign t[246] = t[273] ^ x[86];
  assign t[247] = t[274] ^ x[89];
  assign t[248] = t[275] ^ x[92];
  assign t[249] = (t[276] & ~t[277]);
  assign t[24] = ~(t[36] ^ t[37]);
  assign t[250] = (t[278] & ~t[279]);
  assign t[251] = (t[280] & ~t[281]);
  assign t[252] = (t[282] & ~t[283]);
  assign t[253] = (t[284] & ~t[285]);
  assign t[254] = (t[286] & ~t[287]);
  assign t[255] = (t[288] & ~t[289]);
  assign t[256] = (t[290] & ~t[291]);
  assign t[257] = (t[292] & ~t[293]);
  assign t[258] = (t[294] & ~t[295]);
  assign t[259] = (t[296] & ~t[297]);
  assign t[25] = t[38] ^ t[37];
  assign t[260] = (t[298] & ~t[299]);
  assign t[261] = (t[300] & ~t[301]);
  assign t[262] = (t[302] & ~t[303]);
  assign t[263] = (t[304] & ~t[305]);
  assign t[264] = (t[306] & ~t[307]);
  assign t[265] = (t[308] & ~t[309]);
  assign t[266] = (t[310] & ~t[311]);
  assign t[267] = (t[312] & ~t[313]);
  assign t[268] = (t[314] & ~t[315]);
  assign t[269] = (t[316] & ~t[317]);
  assign t[26] = ~(t[39] ^ t[40]);
  assign t[270] = (t[318] & ~t[319]);
  assign t[271] = (t[320] & ~t[321]);
  assign t[272] = (t[322] & ~t[323]);
  assign t[273] = (t[324] & ~t[325]);
  assign t[274] = (t[326] & ~t[327]);
  assign t[275] = (t[328] & ~t[329]);
  assign t[276] = t[330] ^ x[4];
  assign t[277] = t[331] ^ x[3];
  assign t[278] = t[332] ^ x[7];
  assign t[279] = t[333] ^ x[6];
  assign t[27] = t[9] ? t[41] : t[201];
  assign t[280] = t[334] ^ x[10];
  assign t[281] = t[335] ^ x[9];
  assign t[282] = t[336] ^ x[13];
  assign t[283] = t[337] ^ x[12];
  assign t[284] = t[338] ^ x[18];
  assign t[285] = t[339] ^ x[17];
  assign t[286] = t[340] ^ x[21];
  assign t[287] = t[341] ^ x[20];
  assign t[288] = t[342] ^ x[24];
  assign t[289] = t[343] ^ x[23];
  assign t[28] = t[42] ^ t[43];
  assign t[290] = t[344] ^ x[27];
  assign t[291] = t[345] ^ x[26];
  assign t[292] = t[346] ^ x[30];
  assign t[293] = t[347] ^ x[29];
  assign t[294] = t[348] ^ x[33];
  assign t[295] = t[349] ^ x[32];
  assign t[296] = t[350] ^ x[36];
  assign t[297] = t[351] ^ x[35];
  assign t[298] = t[352] ^ x[41];
  assign t[299] = t[353] ^ x[40];
  assign t[29] = t[44] ^ t[45];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[44];
  assign t[301] = t[355] ^ x[43];
  assign t[302] = t[356] ^ x[47];
  assign t[303] = t[357] ^ x[46];
  assign t[304] = t[358] ^ x[50];
  assign t[305] = t[359] ^ x[49];
  assign t[306] = t[360] ^ x[53];
  assign t[307] = t[361] ^ x[52];
  assign t[308] = t[362] ^ x[56];
  assign t[309] = t[363] ^ x[55];
  assign t[30] = t[46] & t[47];
  assign t[310] = t[364] ^ x[59];
  assign t[311] = t[365] ^ x[58];
  assign t[312] = t[366] ^ x[64];
  assign t[313] = t[367] ^ x[63];
  assign t[314] = t[368] ^ x[67];
  assign t[315] = t[369] ^ x[66];
  assign t[316] = t[370] ^ x[70];
  assign t[317] = t[371] ^ x[69];
  assign t[318] = t[372] ^ x[73];
  assign t[319] = t[373] ^ x[72];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[76];
  assign t[321] = t[375] ^ x[75];
  assign t[322] = t[376] ^ x[79];
  assign t[323] = t[377] ^ x[78];
  assign t[324] = t[378] ^ x[86];
  assign t[325] = t[379] ^ x[85];
  assign t[326] = t[380] ^ x[89];
  assign t[327] = t[381] ^ x[88];
  assign t[328] = t[382] ^ x[92];
  assign t[329] = t[383] ^ x[91];
  assign t[32] = ~(t[50]);
  assign t[330] = (x[2]);
  assign t[331] = (x[2]);
  assign t[332] = (x[5]);
  assign t[333] = (x[5]);
  assign t[334] = (x[8]);
  assign t[335] = (x[8]);
  assign t[336] = (x[11]);
  assign t[337] = (x[11]);
  assign t[338] = (x[16]);
  assign t[339] = (x[16]);
  assign t[33] = ~(t[202]);
  assign t[340] = (x[19]);
  assign t[341] = (x[19]);
  assign t[342] = (x[22]);
  assign t[343] = (x[22]);
  assign t[344] = (x[25]);
  assign t[345] = (x[25]);
  assign t[346] = (x[28]);
  assign t[347] = (x[28]);
  assign t[348] = (x[31]);
  assign t[349] = (x[31]);
  assign t[34] = ~(t[51] ^ t[52]);
  assign t[350] = (x[34]);
  assign t[351] = (x[34]);
  assign t[352] = (x[39]);
  assign t[353] = (x[39]);
  assign t[354] = (x[42]);
  assign t[355] = (x[42]);
  assign t[356] = (x[45]);
  assign t[357] = (x[45]);
  assign t[358] = (x[48]);
  assign t[359] = (x[48]);
  assign t[35] = t[53] ^ t[54];
  assign t[360] = (x[51]);
  assign t[361] = (x[51]);
  assign t[362] = (x[54]);
  assign t[363] = (x[54]);
  assign t[364] = (x[57]);
  assign t[365] = (x[57]);
  assign t[366] = (x[62]);
  assign t[367] = (x[62]);
  assign t[368] = (x[65]);
  assign t[369] = (x[65]);
  assign t[36] = t[55] ^ t[56];
  assign t[370] = (x[68]);
  assign t[371] = (x[68]);
  assign t[372] = (x[71]);
  assign t[373] = (x[71]);
  assign t[374] = (x[74]);
  assign t[375] = (x[74]);
  assign t[376] = (x[77]);
  assign t[377] = (x[77]);
  assign t[378] = (x[84]);
  assign t[379] = (x[84]);
  assign t[37] = t[57] ^ t[43];
  assign t[380] = (x[87]);
  assign t[381] = (x[87]);
  assign t[382] = (x[90]);
  assign t[383] = (x[90]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[60] ^ t[18];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[201] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[9] ? t[68] : t[203];
  assign t[45] = t[196] ^ t[69];
  assign t[46] = ~(t[29] ^ t[70]);
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[204] | t[75];
  assign t[4] = t[9] ? t[10] : t[195];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[71] ^ t[85];
  assign t[56] = t[82] ^ t[86];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] ^ t[61];
  assign t[59] = t[90] & t[91];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[94] ? t[95] : t[205];
  assign t[62] = t[96] ^ t[97];
  assign t[63] = t[98] ? x[38] : x[37];
  assign t[64] = t[99] & t[100];
  assign t[65] = t[101] & t[102];
  assign t[66] = ~(t[57] ^ t[42]);
  assign t[67] = t[103] ^ t[102];
  assign t[68] = t[203] ^ t[104];
  assign t[69] = t[31] ? t[105] : t[206];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[106] ^ t[107];
  assign t[71] = t[45] ^ t[108];
  assign t[72] = t[197] ^ t[109];
  assign t[73] = ~(t[75] & t[110]);
  assign t[74] = ~(t[207] ^ t[111]);
  assign t[75] = ~(t[112] & t[113]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[17] ^ t[114];
  assign t[78] = ~(t[115] ^ t[116]);
  assign t[79] = t[117] ^ t[107];
  assign t[7] = t[15] ^ t[16];
  assign t[80] = t[108] ^ t[118];
  assign t[81] = ~t[119];
  assign t[82] = ~t[120];
  assign t[83] = ~(t[121]);
  assign t[84] = t[122];
  assign t[85] = t[70] ^ t[123];
  assign t[86] = t[124] ^ t[125];
  assign t[87] = t[9] ? t[126] : t[208];
  assign t[88] = t[9] ? t[127] : t[209];
  assign t[89] = t[94] ? t[128] : t[210];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = ~(t[129]);
  assign t[91] = t[94] ? t[130] : t[211];
  assign t[92] = t[121] ^ t[82];
  assign t[93] = t[124] ^ t[131];
  assign t[94] = ~(t[19]);
  assign t[95] = t[205] ^ t[132];
  assign t[96] = t[133] ^ t[59];
  assign t[97] = t[134] & t[135];
  assign t[98] = ~(t[50]);
  assign t[99] = ~(t[136]);
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [116:0] x;
 output y;

 wire [383:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = ~(t[87]);
  assign t[101] = ~(t[88]);
  assign t[102] = t[9] ? t[137] : t[212];
  assign t[103] = t[88] ^ t[27];
  assign t[104] = t[76] ? x[61] : x[60];
  assign t[105] = t[206] ^ t[138];
  assign t[106] = t[139] & t[140];
  assign t[107] = t[141] & t[72];
  assign t[108] = t[200] ^ t[142];
  assign t[109] = t[9] ? t[143] : t[213];
  assign t[10] = t[195] ^ t[20];
  assign t[110] = ~(t[144] & t[145]);
  assign t[111] = t[146] ^ t[214];
  assign t[112] = ~(t[207]);
  assign t[113] = t[147] & t[146];
  assign t[114] = t[148] ^ t[65];
  assign t[115] = ~(t[149] ^ t[40]);
  assign t[116] = t[150] ^ t[151];
  assign t[117] = t[44] ^ t[108];
  assign t[118] = t[70] ^ t[30];
  assign t[119] = t[31] ? t[152] : t[215];
  assign t[11] = ~(t[196]);
  assign t[120] = t[31] ? t[153] : t[216];
  assign t[121] = t[154];
  assign t[122] = t[31] ? t[155] : t[217];
  assign t[123] = t[156] & t[157];
  assign t[124] = t[158] ^ t[54];
  assign t[125] = t[159] & t[160];
  assign t[126] = t[208] ^ t[161];
  assign t[127] = t[209] ^ t[162];
  assign t[128] = t[210] ^ t[163];
  assign t[129] = t[94] ? t[164] : t[218];
  assign t[12] = ~(t[197]);
  assign t[130] = t[211] ^ t[165];
  assign t[131] = t[166] & t[167];
  assign t[132] = t[168] ? x[81] : x[80];
  assign t[133] = t[169] & t[170];
  assign t[134] = ~(t[171] ^ t[96]);
  assign t[135] = t[150] ^ t[91];
  assign t[136] = t[102] ^ t[88];
  assign t[137] = t[212] ^ t[172];
  assign t[138] = t[32] ? x[83] : x[82];
  assign t[139] = ~(t[173]);
  assign t[13] = ~(t[198]);
  assign t[140] = ~(t[44]);
  assign t[141] = ~(t[45]);
  assign t[142] = t[9] ? t[174] : t[219];
  assign t[143] = t[213] ^ t[175];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[176] | t[112]);
  assign t[146] = ~(t[220]);
  assign t[147] = ~(t[214]);
  assign t[148] = t[87] ^ t[27];
  assign t[149] = t[177] ^ t[125];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = t[129] ^ t[61];
  assign t[151] = t[96] ^ t[178];
  assign t[152] = t[215] ^ t[179];
  assign t[153] = t[216] ^ t[180];
  assign t[154] = t[31] ? t[181] : t[221];
  assign t[155] = t[217] ^ t[182];
  assign t[156] = ~(t[106] ^ t[183]);
  assign t[157] = t[117] ^ t[173];
  assign t[158] = t[184] & t[185];
  assign t[159] = ~(t[177] ^ t[124]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[92] ^ t[84];
  assign t[161] = t[98] ? x[94] : x[93];
  assign t[162] = t[98] ? x[96] : x[95];
  assign t[163] = t[168] ? x[98] : x[97];
  assign t[164] = t[218] ^ t[186];
  assign t[165] = t[168] ? x[100] : x[99];
  assign t[166] = ~(t[158] ^ t[187]);
  assign t[167] = t[53] ^ t[188];
  assign t[168] = ~(t[50]);
  assign t[169] = ~(t[189]);
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = ~(t[89]);
  assign t[171] = t[89] ^ t[129];
  assign t[172] = t[98] ? x[102] : x[101];
  assign t[173] = t[72] ^ t[45];
  assign t[174] = t[219] ^ t[190];
  assign t[175] = t[32] ? x[104] : x[103];
  assign t[176] = ~(t[204]);
  assign t[177] = t[81] ^ t[121];
  assign t[178] = t[191] & t[192];
  assign t[179] = t[76] ? x[106] : x[105];
  assign t[17] = t[27] ^ t[28];
  assign t[180] = t[76] ? x[108] : x[107];
  assign t[181] = t[221] ^ t[193];
  assign t[182] = t[98] ? x[110] : x[109];
  assign t[183] = t[71] ^ t[44];
  assign t[184] = ~(t[188]);
  assign t[185] = ~(t[81]);
  assign t[186] = t[168] ? x[112] : x[111];
  assign t[187] = t[92] ^ t[81];
  assign t[188] = t[84] ^ t[121];
  assign t[189] = t[91] ^ t[129];
  assign t[18] = t[29] ^ t[30];
  assign t[190] = t[76] ? x[114] : x[113];
  assign t[191] = ~(t[133] ^ t[194]);
  assign t[192] = t[58] ^ t[189];
  assign t[193] = t[32] ? x[116] : x[115];
  assign t[194] = t[150] ^ t[89];
  assign t[195] = (t[222]);
  assign t[196] = (t[223]);
  assign t[197] = (t[224]);
  assign t[198] = (t[225]);
  assign t[199] = (t[226]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = (t[227]);
  assign t[201] = (t[228]);
  assign t[202] = (t[229]);
  assign t[203] = (t[230]);
  assign t[204] = (t[231]);
  assign t[205] = (t[232]);
  assign t[206] = (t[233]);
  assign t[207] = (t[234]);
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[199]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = t[249] ^ x[4];
  assign t[223] = t[250] ^ x[7];
  assign t[224] = t[251] ^ x[10];
  assign t[225] = t[252] ^ x[13];
  assign t[226] = t[253] ^ x[18];
  assign t[227] = t[254] ^ x[21];
  assign t[228] = t[255] ^ x[24];
  assign t[229] = t[256] ^ x[27];
  assign t[22] = ~(t[33] & t[200]);
  assign t[230] = t[257] ^ x[30];
  assign t[231] = t[258] ^ x[33];
  assign t[232] = t[259] ^ x[36];
  assign t[233] = t[260] ^ x[41];
  assign t[234] = t[261] ^ x[44];
  assign t[235] = t[262] ^ x[47];
  assign t[236] = t[263] ^ x[50];
  assign t[237] = t[264] ^ x[53];
  assign t[238] = t[265] ^ x[56];
  assign t[239] = t[266] ^ x[59];
  assign t[23] = t[34] ^ t[35];
  assign t[240] = t[267] ^ x[64];
  assign t[241] = t[268] ^ x[67];
  assign t[242] = t[269] ^ x[70];
  assign t[243] = t[270] ^ x[73];
  assign t[244] = t[271] ^ x[76];
  assign t[245] = t[272] ^ x[79];
  assign t[246] = t[273] ^ x[86];
  assign t[247] = t[274] ^ x[89];
  assign t[248] = t[275] ^ x[92];
  assign t[249] = (t[276] & ~t[277]);
  assign t[24] = ~(t[36] ^ t[37]);
  assign t[250] = (t[278] & ~t[279]);
  assign t[251] = (t[280] & ~t[281]);
  assign t[252] = (t[282] & ~t[283]);
  assign t[253] = (t[284] & ~t[285]);
  assign t[254] = (t[286] & ~t[287]);
  assign t[255] = (t[288] & ~t[289]);
  assign t[256] = (t[290] & ~t[291]);
  assign t[257] = (t[292] & ~t[293]);
  assign t[258] = (t[294] & ~t[295]);
  assign t[259] = (t[296] & ~t[297]);
  assign t[25] = t[38] ^ t[37];
  assign t[260] = (t[298] & ~t[299]);
  assign t[261] = (t[300] & ~t[301]);
  assign t[262] = (t[302] & ~t[303]);
  assign t[263] = (t[304] & ~t[305]);
  assign t[264] = (t[306] & ~t[307]);
  assign t[265] = (t[308] & ~t[309]);
  assign t[266] = (t[310] & ~t[311]);
  assign t[267] = (t[312] & ~t[313]);
  assign t[268] = (t[314] & ~t[315]);
  assign t[269] = (t[316] & ~t[317]);
  assign t[26] = ~(t[39] ^ t[40]);
  assign t[270] = (t[318] & ~t[319]);
  assign t[271] = (t[320] & ~t[321]);
  assign t[272] = (t[322] & ~t[323]);
  assign t[273] = (t[324] & ~t[325]);
  assign t[274] = (t[326] & ~t[327]);
  assign t[275] = (t[328] & ~t[329]);
  assign t[276] = t[330] ^ x[4];
  assign t[277] = t[331] ^ x[3];
  assign t[278] = t[332] ^ x[7];
  assign t[279] = t[333] ^ x[6];
  assign t[27] = t[9] ? t[41] : t[201];
  assign t[280] = t[334] ^ x[10];
  assign t[281] = t[335] ^ x[9];
  assign t[282] = t[336] ^ x[13];
  assign t[283] = t[337] ^ x[12];
  assign t[284] = t[338] ^ x[18];
  assign t[285] = t[339] ^ x[17];
  assign t[286] = t[340] ^ x[21];
  assign t[287] = t[341] ^ x[20];
  assign t[288] = t[342] ^ x[24];
  assign t[289] = t[343] ^ x[23];
  assign t[28] = t[42] ^ t[43];
  assign t[290] = t[344] ^ x[27];
  assign t[291] = t[345] ^ x[26];
  assign t[292] = t[346] ^ x[30];
  assign t[293] = t[347] ^ x[29];
  assign t[294] = t[348] ^ x[33];
  assign t[295] = t[349] ^ x[32];
  assign t[296] = t[350] ^ x[36];
  assign t[297] = t[351] ^ x[35];
  assign t[298] = t[352] ^ x[41];
  assign t[299] = t[353] ^ x[40];
  assign t[29] = t[44] ^ t[45];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[44];
  assign t[301] = t[355] ^ x[43];
  assign t[302] = t[356] ^ x[47];
  assign t[303] = t[357] ^ x[46];
  assign t[304] = t[358] ^ x[50];
  assign t[305] = t[359] ^ x[49];
  assign t[306] = t[360] ^ x[53];
  assign t[307] = t[361] ^ x[52];
  assign t[308] = t[362] ^ x[56];
  assign t[309] = t[363] ^ x[55];
  assign t[30] = t[46] & t[47];
  assign t[310] = t[364] ^ x[59];
  assign t[311] = t[365] ^ x[58];
  assign t[312] = t[366] ^ x[64];
  assign t[313] = t[367] ^ x[63];
  assign t[314] = t[368] ^ x[67];
  assign t[315] = t[369] ^ x[66];
  assign t[316] = t[370] ^ x[70];
  assign t[317] = t[371] ^ x[69];
  assign t[318] = t[372] ^ x[73];
  assign t[319] = t[373] ^ x[72];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[76];
  assign t[321] = t[375] ^ x[75];
  assign t[322] = t[376] ^ x[79];
  assign t[323] = t[377] ^ x[78];
  assign t[324] = t[378] ^ x[86];
  assign t[325] = t[379] ^ x[85];
  assign t[326] = t[380] ^ x[89];
  assign t[327] = t[381] ^ x[88];
  assign t[328] = t[382] ^ x[92];
  assign t[329] = t[383] ^ x[91];
  assign t[32] = ~(t[50]);
  assign t[330] = (x[2]);
  assign t[331] = (x[2]);
  assign t[332] = (x[5]);
  assign t[333] = (x[5]);
  assign t[334] = (x[8]);
  assign t[335] = (x[8]);
  assign t[336] = (x[11]);
  assign t[337] = (x[11]);
  assign t[338] = (x[16]);
  assign t[339] = (x[16]);
  assign t[33] = ~(t[202]);
  assign t[340] = (x[19]);
  assign t[341] = (x[19]);
  assign t[342] = (x[22]);
  assign t[343] = (x[22]);
  assign t[344] = (x[25]);
  assign t[345] = (x[25]);
  assign t[346] = (x[28]);
  assign t[347] = (x[28]);
  assign t[348] = (x[31]);
  assign t[349] = (x[31]);
  assign t[34] = ~(t[51] ^ t[52]);
  assign t[350] = (x[34]);
  assign t[351] = (x[34]);
  assign t[352] = (x[39]);
  assign t[353] = (x[39]);
  assign t[354] = (x[42]);
  assign t[355] = (x[42]);
  assign t[356] = (x[45]);
  assign t[357] = (x[45]);
  assign t[358] = (x[48]);
  assign t[359] = (x[48]);
  assign t[35] = t[53] ^ t[54];
  assign t[360] = (x[51]);
  assign t[361] = (x[51]);
  assign t[362] = (x[54]);
  assign t[363] = (x[54]);
  assign t[364] = (x[57]);
  assign t[365] = (x[57]);
  assign t[366] = (x[62]);
  assign t[367] = (x[62]);
  assign t[368] = (x[65]);
  assign t[369] = (x[65]);
  assign t[36] = t[55] ^ t[56];
  assign t[370] = (x[68]);
  assign t[371] = (x[68]);
  assign t[372] = (x[71]);
  assign t[373] = (x[71]);
  assign t[374] = (x[74]);
  assign t[375] = (x[74]);
  assign t[376] = (x[77]);
  assign t[377] = (x[77]);
  assign t[378] = (x[84]);
  assign t[379] = (x[84]);
  assign t[37] = t[57] ^ t[43];
  assign t[380] = (x[87]);
  assign t[381] = (x[87]);
  assign t[382] = (x[90]);
  assign t[383] = (x[90]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = t[60] ^ t[18];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[201] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[9] ? t[68] : t[203];
  assign t[45] = t[196] ^ t[69];
  assign t[46] = ~(t[29] ^ t[70]);
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[204] | t[75];
  assign t[4] = t[9] ? t[10] : t[195];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] & t[84];
  assign t[55] = t[71] ^ t[85];
  assign t[56] = t[82] ^ t[86];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] ^ t[61];
  assign t[59] = t[90] & t[91];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = t[94] ? t[95] : t[205];
  assign t[62] = t[96] ^ t[97];
  assign t[63] = t[98] ? x[38] : x[37];
  assign t[64] = t[99] & t[100];
  assign t[65] = t[101] & t[102];
  assign t[66] = ~(t[57] ^ t[42]);
  assign t[67] = t[103] ^ t[102];
  assign t[68] = t[203] ^ t[104];
  assign t[69] = t[31] ? t[105] : t[206];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[106] ^ t[107];
  assign t[71] = t[45] ^ t[108];
  assign t[72] = t[197] ^ t[109];
  assign t[73] = ~(t[75] & t[110]);
  assign t[74] = ~(t[207] ^ t[111]);
  assign t[75] = ~(t[112] & t[113]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[17] ^ t[114];
  assign t[78] = ~(t[115] ^ t[116]);
  assign t[79] = t[117] ^ t[107];
  assign t[7] = t[15] ^ t[16];
  assign t[80] = t[108] ^ t[118];
  assign t[81] = ~t[119];
  assign t[82] = ~t[120];
  assign t[83] = ~(t[121]);
  assign t[84] = t[122];
  assign t[85] = t[70] ^ t[123];
  assign t[86] = t[124] ^ t[125];
  assign t[87] = t[9] ? t[126] : t[208];
  assign t[88] = t[9] ? t[127] : t[209];
  assign t[89] = t[94] ? t[128] : t[210];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = ~(t[129]);
  assign t[91] = t[94] ? t[130] : t[211];
  assign t[92] = t[121] ^ t[82];
  assign t[93] = t[124] ^ t[131];
  assign t[94] = ~(t[19]);
  assign t[95] = t[205] ^ t[132];
  assign t[96] = t[133] ^ t[59];
  assign t[97] = t[134] & t[135];
  assign t[98] = ~(t[50]);
  assign t[99] = ~(t[136]);
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[31] ? t[143] : t[226];
  assign t[101] = t[144] ? x[56] : x[55];
  assign t[102] = ~(t[114] ^ t[56]);
  assign t[103] = t[36] ^ t[124];
  assign t[104] = t[32] ? x[58] : x[57];
  assign t[105] = t[145] & t[146];
  assign t[106] = t[147] & t[148];
  assign t[107] = ~(t[91] ^ t[71]);
  assign t[108] = t[149] ^ t[148];
  assign t[109] = ~(t[150] & t[151]);
  assign t[10] = t[210] ^ t[20];
  assign t[110] = t[152] ^ t[227];
  assign t[111] = ~(t[222]);
  assign t[112] = t[153] & t[152];
  assign t[113] = t[154] ^ t[61];
  assign t[114] = t[155] ^ t[55];
  assign t[115] = t[119] ^ t[156];
  assign t[116] = t[62] ^ t[157];
  assign t[117] = t[31] ? t[158] : t[228];
  assign t[118] = t[159] ^ t[43];
  assign t[119] = t[81] ^ t[65];
  assign t[11] = ~(t[211]);
  assign t[120] = t[144] ? x[66] : x[65];
  assign t[121] = ~(t[127]);
  assign t[122] = ~(t[155]);
  assign t[123] = ~(t[55]);
  assign t[124] = t[9] ? t[160] : t[229];
  assign t[125] = t[36] ^ t[155];
  assign t[126] = t[155] ^ t[44];
  assign t[127] = t[124] ^ t[55];
  assign t[128] = ~(t[161] ^ t[162]);
  assign t[129] = t[163] ^ t[164];
  assign t[12] = ~(t[212]);
  assign t[130] = t[9] ? t[165] : t[230];
  assign t[131] = t[9] ? t[166] : t[231];
  assign t[132] = t[223] ^ t[167];
  assign t[133] = t[224] ^ t[168];
  assign t[134] = ~(t[139]);
  assign t[135] = ~(t[154]);
  assign t[136] = ~(t[60]);
  assign t[137] = t[169];
  assign t[138] = t[40] ^ t[154];
  assign t[139] = t[137] ^ t[60];
  assign t[13] = ~(t[213]);
  assign t[140] = t[144] ? x[77] : x[76];
  assign t[141] = ~(t[19]);
  assign t[142] = t[225] ^ t[170];
  assign t[143] = t[226] ^ t[171];
  assign t[144] = ~(t[50]);
  assign t[145] = ~(t[172]);
  assign t[146] = ~(t[130]);
  assign t[147] = ~(t[131]);
  assign t[148] = t[9] ? t[173] : t[232];
  assign t[149] = t[131] ^ t[46];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = ~(t[153] | t[152]);
  assign t[151] = ~(t[174] | t[111]);
  assign t[152] = ~(t[233]);
  assign t[153] = ~(t[227]);
  assign t[154] = ~t[175];
  assign t[155] = t[9] ? t[176] : t[234];
  assign t[156] = t[118] ^ t[177];
  assign t[157] = t[178] & t[179];
  assign t[158] = t[228] ^ t[180];
  assign t[159] = t[181] & t[182];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[229] ^ t[183];
  assign t[161] = t[184] ^ t[185];
  assign t[162] = ~(t[186] ^ t[30]);
  assign t[163] = t[149] ^ t[187];
  assign t[164] = t[65] ^ t[188];
  assign t[165] = t[230] ^ t[189];
  assign t[166] = t[231] ^ t[190];
  assign t[167] = t[191] ? x[88] : x[87];
  assign t[168] = t[76] ? x[90] : x[89];
  assign t[169] = t[31] ? t[192] : t[235];
  assign t[16] = t[25] ^ t[26];
  assign t[170] = t[191] ? x[95] : x[94];
  assign t[171] = t[76] ? x[97] : x[96];
  assign t[172] = t[148] ^ t[131];
  assign t[173] = t[232] ^ t[193];
  assign t[174] = ~(t[219]);
  assign t[175] = t[31] ? t[194] : t[236];
  assign t[176] = t[234] ^ t[195];
  assign t[177] = t[196] & t[197];
  assign t[178] = ~(t[198] ^ t[62]);
  assign t[179] = t[40] ^ t[137];
  assign t[17] = t[27] ^ t[28];
  assign t[180] = t[144] ? x[102] : x[101];
  assign t[181] = ~(t[199]);
  assign t[182] = ~(t[64]);
  assign t[183] = t[144] ? x[104] : x[103];
  assign t[184] = t[29] ^ t[200];
  assign t[185] = ~(t[201] ^ t[27]);
  assign t[186] = t[202] ^ t[106];
  assign t[187] = t[71] ^ t[203];
  assign t[188] = t[118] ^ t[54];
  assign t[189] = t[32] ? x[106] : x[105];
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[190] = t[32] ? x[108] : x[107];
  assign t[191] = ~(t[50]);
  assign t[192] = t[235] ^ t[204];
  assign t[193] = t[32] ? x[110] : x[109];
  assign t[194] = t[236] ^ t[205];
  assign t[195] = t[144] ? x[112] : x[111];
  assign t[196] = ~(t[159] ^ t[206]);
  assign t[197] = t[42] ^ t[199];
  assign t[198] = t[154] ^ t[60];
  assign t[199] = t[67] ^ t[81];
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[126] ^ t[86];
  assign t[201] = ~(t[35] ^ t[80]);
  assign t[202] = t[130] ^ t[46];
  assign t[203] = t[207] & t[208];
  assign t[204] = t[191] ? x[114] : x[113];
  assign t[205] = t[76] ? x[116] : x[115];
  assign t[206] = t[119] ^ t[64];
  assign t[207] = ~(t[105] ^ t[209]);
  assign t[208] = t[202] ^ t[172];
  assign t[209] = t[149] ^ t[130];
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[214]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[33] & t[215]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[7];
  assign t[239] = t[266] ^ x[10];
  assign t[23] = t[34] ^ t[35];
  assign t[240] = t[267] ^ x[13];
  assign t[241] = t[268] ^ x[18];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = ~(t[25] ^ t[30]);
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[51];
  assign t[253] = t[280] ^ x[54];
  assign t[254] = t[281] ^ x[61];
  assign t[255] = t[282] ^ x[64];
  assign t[256] = t[283] ^ x[69];
  assign t[257] = t[284] ^ x[72];
  assign t[258] = t[285] ^ x[75];
  assign t[259] = t[286] ^ x[80];
  assign t[25] = t[36] ^ t[37];
  assign t[260] = t[287] ^ x[83];
  assign t[261] = t[288] ^ x[86];
  assign t[262] = t[289] ^ x[93];
  assign t[263] = t[290] ^ x[100];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = t[42] ^ t[43];
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[7];
  assign t[294] = t[348] ^ x[6];
  assign t[295] = t[349] ^ x[10];
  assign t[296] = t[350] ^ x[9];
  assign t[297] = t[351] ^ x[13];
  assign t[298] = t[352] ^ x[12];
  assign t[299] = t[353] ^ x[18];
  assign t[29] = t[44] ^ t[45];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[17];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = t[46] ^ t[47];
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[51];
  assign t[322] = t[376] ^ x[50];
  assign t[323] = t[377] ^ x[54];
  assign t[324] = t[378] ^ x[53];
  assign t[325] = t[379] ^ x[61];
  assign t[326] = t[380] ^ x[60];
  assign t[327] = t[381] ^ x[64];
  assign t[328] = t[382] ^ x[63];
  assign t[329] = t[383] ^ x[69];
  assign t[32] = ~(t[50]);
  assign t[330] = t[384] ^ x[68];
  assign t[331] = t[385] ^ x[72];
  assign t[332] = t[386] ^ x[71];
  assign t[333] = t[387] ^ x[75];
  assign t[334] = t[388] ^ x[74];
  assign t[335] = t[389] ^ x[80];
  assign t[336] = t[390] ^ x[79];
  assign t[337] = t[391] ^ x[83];
  assign t[338] = t[392] ^ x[82];
  assign t[339] = t[393] ^ x[86];
  assign t[33] = ~(t[216]);
  assign t[340] = t[394] ^ x[85];
  assign t[341] = t[395] ^ x[93];
  assign t[342] = t[396] ^ x[92];
  assign t[343] = t[397] ^ x[100];
  assign t[344] = t[398] ^ x[99];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[5]);
  assign t[348] = (x[5]);
  assign t[349] = (x[8]);
  assign t[34] = ~(t[51] ^ t[52]);
  assign t[350] = (x[8]);
  assign t[351] = (x[11]);
  assign t[352] = (x[11]);
  assign t[353] = (x[16]);
  assign t[354] = (x[16]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = t[53] ^ t[54];
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = t[55] ^ t[44];
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[49]);
  assign t[376] = (x[49]);
  assign t[377] = (x[52]);
  assign t[378] = (x[52]);
  assign t[379] = (x[59]);
  assign t[37] = t[56] ^ t[57];
  assign t[380] = (x[59]);
  assign t[381] = (x[62]);
  assign t[382] = (x[62]);
  assign t[383] = (x[67]);
  assign t[384] = (x[67]);
  assign t[385] = (x[70]);
  assign t[386] = (x[70]);
  assign t[387] = (x[73]);
  assign t[388] = (x[73]);
  assign t[389] = (x[78]);
  assign t[38] = t[58] ^ t[34];
  assign t[390] = (x[78]);
  assign t[391] = (x[81]);
  assign t[392] = (x[81]);
  assign t[393] = (x[84]);
  assign t[394] = (x[84]);
  assign t[395] = (x[91]);
  assign t[396] = (x[91]);
  assign t[397] = (x[98]);
  assign t[398] = (x[98]);
  assign t[39] = ~(t[29] ^ t[59]);
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[9] ? t[68] : t[217];
  assign t[45] = t[56] ^ t[69];
  assign t[46] = t[9] ? t[70] : t[218];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[219] | t[75];
  assign t[4] = t[9] ? t[10] : t[210];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[64] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = t[9] ? t[84] : t[220];
  assign t[56] = t[85] ^ t[86];
  assign t[57] = t[87] & t[88];
  assign t[58] = ~(t[89] ^ t[90]);
  assign t[59] = t[91] ^ t[72];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[92];
  assign t[61] = t[93];
  assign t[62] = t[94] ^ t[95];
  assign t[63] = t[96] & t[97];
  assign t[64] = t[31] ? t[98] : t[221];
  assign t[65] = t[214] ^ t[99];
  assign t[66] = ~(t[81]);
  assign t[67] = t[216] ^ t[100];
  assign t[68] = t[217] ^ t[101];
  assign t[69] = t[102] & t[103];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[218] ^ t[104];
  assign t[71] = t[105] ^ t[106];
  assign t[72] = t[107] & t[108];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[222] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[113] ^ t[95];
  assign t[78] = t[114] ^ t[69];
  assign t[79] = t[115] ^ t[59];
  assign t[7] = ~(t[15] ^ t[16]);
  assign t[80] = t[61] ^ t[116];
  assign t[81] = t[213] ^ t[117];
  assign t[82] = ~(t[53] ^ t[118]);
  assign t[83] = t[119] ^ t[67];
  assign t[84] = t[220] ^ t[120];
  assign t[85] = t[121] & t[122];
  assign t[86] = t[123] & t[124];
  assign t[87] = ~(t[85] ^ t[125]);
  assign t[88] = t[126] ^ t[127];
  assign t[89] = t[128] ^ t[28];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = ~(t[129] ^ t[78]);
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[31] ? t[132] : t[223];
  assign t[93] = t[31] ? t[133] : t[224];
  assign t[94] = t[134] & t[135];
  assign t[95] = t[136] & t[137];
  assign t[96] = ~(t[94] ^ t[138]);
  assign t[97] = t[113] ^ t[139];
  assign t[98] = t[221] ^ t[140];
  assign t[99] = t[141] ? t[142] : t[225];
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind121(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[31] ? t[143] : t[226];
  assign t[101] = t[144] ? x[56] : x[55];
  assign t[102] = ~(t[114] ^ t[56]);
  assign t[103] = t[36] ^ t[124];
  assign t[104] = t[32] ? x[58] : x[57];
  assign t[105] = t[145] & t[146];
  assign t[106] = t[147] & t[148];
  assign t[107] = ~(t[91] ^ t[71]);
  assign t[108] = t[149] ^ t[148];
  assign t[109] = ~(t[150] & t[151]);
  assign t[10] = t[210] ^ t[20];
  assign t[110] = t[152] ^ t[227];
  assign t[111] = ~(t[222]);
  assign t[112] = t[153] & t[152];
  assign t[113] = t[154] ^ t[61];
  assign t[114] = t[155] ^ t[55];
  assign t[115] = t[119] ^ t[156];
  assign t[116] = t[62] ^ t[157];
  assign t[117] = t[31] ? t[158] : t[228];
  assign t[118] = t[159] ^ t[43];
  assign t[119] = t[81] ^ t[65];
  assign t[11] = ~(t[211]);
  assign t[120] = t[144] ? x[66] : x[65];
  assign t[121] = ~(t[127]);
  assign t[122] = ~(t[155]);
  assign t[123] = ~(t[55]);
  assign t[124] = t[9] ? t[160] : t[229];
  assign t[125] = t[36] ^ t[155];
  assign t[126] = t[155] ^ t[44];
  assign t[127] = t[124] ^ t[55];
  assign t[128] = ~(t[161] ^ t[162]);
  assign t[129] = t[163] ^ t[164];
  assign t[12] = ~(t[212]);
  assign t[130] = t[9] ? t[165] : t[230];
  assign t[131] = t[9] ? t[166] : t[231];
  assign t[132] = t[223] ^ t[167];
  assign t[133] = t[224] ^ t[168];
  assign t[134] = ~(t[139]);
  assign t[135] = ~(t[154]);
  assign t[136] = ~(t[60]);
  assign t[137] = t[169];
  assign t[138] = t[40] ^ t[154];
  assign t[139] = t[137] ^ t[60];
  assign t[13] = ~(t[213]);
  assign t[140] = t[144] ? x[77] : x[76];
  assign t[141] = ~(t[19]);
  assign t[142] = t[225] ^ t[170];
  assign t[143] = t[226] ^ t[171];
  assign t[144] = ~(t[50]);
  assign t[145] = ~(t[172]);
  assign t[146] = ~(t[130]);
  assign t[147] = ~(t[131]);
  assign t[148] = t[9] ? t[173] : t[232];
  assign t[149] = t[131] ^ t[46];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = ~(t[153] | t[152]);
  assign t[151] = ~(t[174] | t[111]);
  assign t[152] = ~(t[233]);
  assign t[153] = ~(t[227]);
  assign t[154] = ~t[175];
  assign t[155] = t[9] ? t[176] : t[234];
  assign t[156] = t[118] ^ t[177];
  assign t[157] = t[178] & t[179];
  assign t[158] = t[228] ^ t[180];
  assign t[159] = t[181] & t[182];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[229] ^ t[183];
  assign t[161] = t[184] ^ t[185];
  assign t[162] = ~(t[186] ^ t[30]);
  assign t[163] = t[149] ^ t[187];
  assign t[164] = t[65] ^ t[188];
  assign t[165] = t[230] ^ t[189];
  assign t[166] = t[231] ^ t[190];
  assign t[167] = t[191] ? x[88] : x[87];
  assign t[168] = t[76] ? x[90] : x[89];
  assign t[169] = t[31] ? t[192] : t[235];
  assign t[16] = t[25] ^ t[26];
  assign t[170] = t[191] ? x[95] : x[94];
  assign t[171] = t[76] ? x[97] : x[96];
  assign t[172] = t[148] ^ t[131];
  assign t[173] = t[232] ^ t[193];
  assign t[174] = ~(t[219]);
  assign t[175] = t[31] ? t[194] : t[236];
  assign t[176] = t[234] ^ t[195];
  assign t[177] = t[196] & t[197];
  assign t[178] = ~(t[198] ^ t[62]);
  assign t[179] = t[40] ^ t[137];
  assign t[17] = t[27] ^ t[28];
  assign t[180] = t[144] ? x[102] : x[101];
  assign t[181] = ~(t[199]);
  assign t[182] = ~(t[64]);
  assign t[183] = t[144] ? x[104] : x[103];
  assign t[184] = t[29] ^ t[200];
  assign t[185] = ~(t[201] ^ t[27]);
  assign t[186] = t[202] ^ t[106];
  assign t[187] = t[71] ^ t[203];
  assign t[188] = t[118] ^ t[54];
  assign t[189] = t[32] ? x[106] : x[105];
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[190] = t[32] ? x[108] : x[107];
  assign t[191] = ~(t[50]);
  assign t[192] = t[235] ^ t[204];
  assign t[193] = t[32] ? x[110] : x[109];
  assign t[194] = t[236] ^ t[205];
  assign t[195] = t[144] ? x[112] : x[111];
  assign t[196] = ~(t[159] ^ t[206]);
  assign t[197] = t[42] ^ t[199];
  assign t[198] = t[154] ^ t[60];
  assign t[199] = t[67] ^ t[81];
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[126] ^ t[86];
  assign t[201] = ~(t[35] ^ t[80]);
  assign t[202] = t[130] ^ t[46];
  assign t[203] = t[207] & t[208];
  assign t[204] = t[191] ? x[114] : x[113];
  assign t[205] = t[76] ? x[116] : x[115];
  assign t[206] = t[119] ^ t[64];
  assign t[207] = ~(t[105] ^ t[209]);
  assign t[208] = t[202] ^ t[172];
  assign t[209] = t[149] ^ t[130];
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[214]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[33] & t[215]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[7];
  assign t[239] = t[266] ^ x[10];
  assign t[23] = t[34] ^ t[35];
  assign t[240] = t[267] ^ x[13];
  assign t[241] = t[268] ^ x[18];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = ~(t[25] ^ t[30]);
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[51];
  assign t[253] = t[280] ^ x[54];
  assign t[254] = t[281] ^ x[61];
  assign t[255] = t[282] ^ x[64];
  assign t[256] = t[283] ^ x[69];
  assign t[257] = t[284] ^ x[72];
  assign t[258] = t[285] ^ x[75];
  assign t[259] = t[286] ^ x[80];
  assign t[25] = t[36] ^ t[37];
  assign t[260] = t[287] ^ x[83];
  assign t[261] = t[288] ^ x[86];
  assign t[262] = t[289] ^ x[93];
  assign t[263] = t[290] ^ x[100];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = t[42] ^ t[43];
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[7];
  assign t[294] = t[348] ^ x[6];
  assign t[295] = t[349] ^ x[10];
  assign t[296] = t[350] ^ x[9];
  assign t[297] = t[351] ^ x[13];
  assign t[298] = t[352] ^ x[12];
  assign t[299] = t[353] ^ x[18];
  assign t[29] = t[44] ^ t[45];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[17];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = t[46] ^ t[47];
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[51];
  assign t[322] = t[376] ^ x[50];
  assign t[323] = t[377] ^ x[54];
  assign t[324] = t[378] ^ x[53];
  assign t[325] = t[379] ^ x[61];
  assign t[326] = t[380] ^ x[60];
  assign t[327] = t[381] ^ x[64];
  assign t[328] = t[382] ^ x[63];
  assign t[329] = t[383] ^ x[69];
  assign t[32] = ~(t[50]);
  assign t[330] = t[384] ^ x[68];
  assign t[331] = t[385] ^ x[72];
  assign t[332] = t[386] ^ x[71];
  assign t[333] = t[387] ^ x[75];
  assign t[334] = t[388] ^ x[74];
  assign t[335] = t[389] ^ x[80];
  assign t[336] = t[390] ^ x[79];
  assign t[337] = t[391] ^ x[83];
  assign t[338] = t[392] ^ x[82];
  assign t[339] = t[393] ^ x[86];
  assign t[33] = ~(t[216]);
  assign t[340] = t[394] ^ x[85];
  assign t[341] = t[395] ^ x[93];
  assign t[342] = t[396] ^ x[92];
  assign t[343] = t[397] ^ x[100];
  assign t[344] = t[398] ^ x[99];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[5]);
  assign t[348] = (x[5]);
  assign t[349] = (x[8]);
  assign t[34] = ~(t[51] ^ t[52]);
  assign t[350] = (x[8]);
  assign t[351] = (x[11]);
  assign t[352] = (x[11]);
  assign t[353] = (x[16]);
  assign t[354] = (x[16]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = t[53] ^ t[54];
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = t[55] ^ t[44];
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[49]);
  assign t[376] = (x[49]);
  assign t[377] = (x[52]);
  assign t[378] = (x[52]);
  assign t[379] = (x[59]);
  assign t[37] = t[56] ^ t[57];
  assign t[380] = (x[59]);
  assign t[381] = (x[62]);
  assign t[382] = (x[62]);
  assign t[383] = (x[67]);
  assign t[384] = (x[67]);
  assign t[385] = (x[70]);
  assign t[386] = (x[70]);
  assign t[387] = (x[73]);
  assign t[388] = (x[73]);
  assign t[389] = (x[78]);
  assign t[38] = t[58] ^ t[34];
  assign t[390] = (x[78]);
  assign t[391] = (x[81]);
  assign t[392] = (x[81]);
  assign t[393] = (x[84]);
  assign t[394] = (x[84]);
  assign t[395] = (x[91]);
  assign t[396] = (x[91]);
  assign t[397] = (x[98]);
  assign t[398] = (x[98]);
  assign t[39] = ~(t[29] ^ t[59]);
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = t[9] ? t[68] : t[217];
  assign t[45] = t[56] ^ t[69];
  assign t[46] = t[9] ? t[70] : t[218];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[219] | t[75];
  assign t[4] = t[9] ? t[10] : t[210];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[64] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = t[9] ? t[84] : t[220];
  assign t[56] = t[85] ^ t[86];
  assign t[57] = t[87] & t[88];
  assign t[58] = ~(t[89] ^ t[90]);
  assign t[59] = t[91] ^ t[72];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[92];
  assign t[61] = t[93];
  assign t[62] = t[94] ^ t[95];
  assign t[63] = t[96] & t[97];
  assign t[64] = t[31] ? t[98] : t[221];
  assign t[65] = t[214] ^ t[99];
  assign t[66] = ~(t[81]);
  assign t[67] = t[216] ^ t[100];
  assign t[68] = t[217] ^ t[101];
  assign t[69] = t[102] & t[103];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[218] ^ t[104];
  assign t[71] = t[105] ^ t[106];
  assign t[72] = t[107] & t[108];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[222] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[113] ^ t[95];
  assign t[78] = t[114] ^ t[69];
  assign t[79] = t[115] ^ t[59];
  assign t[7] = ~(t[15] ^ t[16]);
  assign t[80] = t[61] ^ t[116];
  assign t[81] = t[213] ^ t[117];
  assign t[82] = ~(t[53] ^ t[118]);
  assign t[83] = t[119] ^ t[67];
  assign t[84] = t[220] ^ t[120];
  assign t[85] = t[121] & t[122];
  assign t[86] = t[123] & t[124];
  assign t[87] = ~(t[85] ^ t[125]);
  assign t[88] = t[126] ^ t[127];
  assign t[89] = t[128] ^ t[28];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = ~(t[129] ^ t[78]);
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[31] ? t[132] : t[223];
  assign t[93] = t[31] ? t[133] : t[224];
  assign t[94] = t[134] & t[135];
  assign t[95] = t[136] & t[137];
  assign t[96] = ~(t[94] ^ t[138]);
  assign t[97] = t[113] ^ t[139];
  assign t[98] = t[221] ^ t[140];
  assign t[99] = t[141] ? t[142] : t[225];
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [116:0] x;
 output y;

 wire [407:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[142] ^ t[143];
  assign t[101] = t[128] ^ t[59];
  assign t[102] = t[43] ^ t[84];
  assign t[103] = t[144] ^ t[145];
  assign t[104] = t[31] ? t[146] : t[233];
  assign t[105] = ~(t[69] ^ t[96]);
  assign t[106] = t[64] ^ t[147];
  assign t[107] = t[228] ^ t[148];
  assign t[108] = t[149] ^ t[63];
  assign t[109] = t[150] & t[151];
  assign t[10] = t[219] ^ t[20];
  assign t[110] = ~(t[152] & t[153]);
  assign t[111] = t[154] ^ t[234];
  assign t[112] = ~(t[229]);
  assign t[113] = t[155] & t[154];
  assign t[114] = t[9] ? t[156] : t[235];
  assign t[115] = ~(t[81]);
  assign t[116] = t[9] ? t[157] : t[236];
  assign t[117] = t[9] ? t[158] : t[237];
  assign t[118] = t[159] & t[160];
  assign t[119] = t[230] ^ t[161];
  assign t[11] = ~(t[220]);
  assign t[120] = ~(t[86] ^ t[162]);
  assign t[121] = t[77] ^ t[163];
  assign t[122] = t[26] ^ t[164];
  assign t[123] = ~(t[98] ^ t[101]);
  assign t[124] = t[91] ^ t[117];
  assign t[125] = ~(t[50]);
  assign t[126] = ~(t[163]);
  assign t[127] = ~(t[114]);
  assign t[128] = t[114] ^ t[81];
  assign t[129] = t[165] ^ t[144];
  assign t[12] = ~(t[221]);
  assign t[130] = t[166] ^ t[167];
  assign t[131] = t[231] ^ t[168];
  assign t[132] = t[232] ^ t[169];
  assign t[133] = t[31] ? t[170] : t[238];
  assign t[134] = t[171] ? t[172] : t[239];
  assign t[135] = t[173] & t[174];
  assign t[136] = t[175] & t[147];
  assign t[137] = ~(t[135] ^ t[176]);
  assign t[138] = t[177] ^ t[178];
  assign t[139] = t[95] ^ t[179];
  assign t[13] = ~(t[222]);
  assign t[140] = t[180] ^ t[165];
  assign t[141] = t[181] & t[182];
  assign t[142] = t[180] ^ t[144];
  assign t[143] = t[183] & t[184];
  assign t[144] = t[185];
  assign t[145] = t[166] ^ t[141];
  assign t[146] = t[233] ^ t[186];
  assign t[147] = t[225] ^ t[187];
  assign t[148] = t[32] ? x[70] : x[69];
  assign t[149] = t[188] & t[189];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = ~(t[124] ^ t[108]);
  assign t[151] = t[79] ^ t[93];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[190] | t[112]);
  assign t[154] = ~(t[240]);
  assign t[155] = ~(t[234]);
  assign t[156] = t[235] ^ t[191];
  assign t[157] = t[236] ^ t[192];
  assign t[158] = t[237] ^ t[193];
  assign t[159] = ~(t[149] ^ t[194]);
  assign t[15] = t[23] ^ t[24];
  assign t[160] = t[62] ^ t[195];
  assign t[161] = t[125] ? x[75] : x[74];
  assign t[162] = t[53] ^ t[114];
  assign t[163] = t[116] ^ t[81];
  assign t[164] = t[177] ^ t[136];
  assign t[165] = t[196];
  assign t[166] = t[197] ^ t[143];
  assign t[167] = t[198] & t[199];
  assign t[168] = t[32] ? x[77] : x[76];
  assign t[169] = t[32] ? x[79] : x[78];
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = t[238] ^ t[200];
  assign t[171] = ~(t[19]);
  assign t[172] = t[239] ^ t[201];
  assign t[173] = ~(t[178]);
  assign t[174] = ~(t[104]);
  assign t[175] = ~(t[94]);
  assign t[176] = t[64] ^ t[104];
  assign t[177] = t[104] ^ t[95];
  assign t[178] = t[147] ^ t[94];
  assign t[179] = t[96] ^ t[70];
  assign t[17] = ~(t[27] ^ t[28]);
  assign t[180] = ~t[202];
  assign t[181] = ~(t[140] ^ t[166]);
  assign t[182] = t[129] ^ t[184];
  assign t[183] = ~(t[165]);
  assign t[184] = t[203];
  assign t[185] = t[31] ? t[204] : t[241];
  assign t[186] = t[125] ? x[84] : x[83];
  assign t[187] = t[31] ? t[205] : t[242];
  assign t[188] = ~(t[195]);
  assign t[189] = ~(t[91]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[190] = ~(t[227]);
  assign t[191] = t[125] ? x[89] : x[88];
  assign t[192] = t[125] ? x[91] : x[90];
  assign t[193] = t[32] ? x[93] : x[92];
  assign t[194] = t[79] ^ t[91];
  assign t[195] = t[93] ^ t[117];
  assign t[196] = t[31] ? t[206] : t[243];
  assign t[197] = t[207] & t[208];
  assign t[198] = ~(t[197] ^ t[209]);
  assign t[199] = t[142] ^ t[210];
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[125] ? x[98] : x[97];
  assign t[201] = t[211] ? x[100] : x[99];
  assign t[202] = t[31] ? t[212] : t[244];
  assign t[203] = t[31] ? t[213] : t[245];
  assign t[204] = t[241] ^ t[214];
  assign t[205] = t[242] ^ t[215];
  assign t[206] = t[243] ^ t[216];
  assign t[207] = ~(t[210]);
  assign t[208] = ~(t[180]);
  assign t[209] = t[129] ^ t[180];
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = t[184] ^ t[165];
  assign t[211] = ~(t[50]);
  assign t[212] = t[244] ^ t[217];
  assign t[213] = t[245] ^ t[218];
  assign t[214] = t[76] ? x[108] : x[107];
  assign t[215] = t[76] ? x[110] : x[109];
  assign t[216] = t[211] ? x[112] : x[111];
  assign t[217] = t[76] ? x[114] : x[113];
  assign t[218] = t[211] ? x[116] : x[115];
  assign t[219] = (t[246]);
  assign t[21] = ~(t[223]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[33] & t[224]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = (t[266]);
  assign t[23] = ~(t[34] ^ t[35]);
  assign t[240] = (t[267]);
  assign t[241] = (t[268]);
  assign t[242] = (t[269]);
  assign t[243] = (t[270]);
  assign t[244] = (t[271]);
  assign t[245] = (t[272]);
  assign t[246] = t[273] ^ x[4];
  assign t[247] = t[274] ^ x[7];
  assign t[248] = t[275] ^ x[10];
  assign t[249] = t[276] ^ x[13];
  assign t[24] = t[36] ^ t[37];
  assign t[250] = t[277] ^ x[18];
  assign t[251] = t[278] ^ x[21];
  assign t[252] = t[279] ^ x[24];
  assign t[253] = t[280] ^ x[27];
  assign t[254] = t[281] ^ x[30];
  assign t[255] = t[282] ^ x[33];
  assign t[256] = t[283] ^ x[36];
  assign t[257] = t[284] ^ x[39];
  assign t[258] = t[285] ^ x[44];
  assign t[259] = t[286] ^ x[47];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[287] ^ x[50];
  assign t[261] = t[288] ^ x[53];
  assign t[262] = t[289] ^ x[56];
  assign t[263] = t[290] ^ x[59];
  assign t[264] = t[291] ^ x[62];
  assign t[265] = t[292] ^ x[65];
  assign t[266] = t[293] ^ x[68];
  assign t[267] = t[294] ^ x[73];
  assign t[268] = t[295] ^ x[82];
  assign t[269] = t[296] ^ x[87];
  assign t[26] = ~(t[40] ^ t[41]);
  assign t[270] = t[297] ^ x[96];
  assign t[271] = t[298] ^ x[103];
  assign t[272] = t[299] ^ x[106];
  assign t[273] = (t[300] & ~t[301]);
  assign t[274] = (t[302] & ~t[303]);
  assign t[275] = (t[304] & ~t[305]);
  assign t[276] = (t[306] & ~t[307]);
  assign t[277] = (t[308] & ~t[309]);
  assign t[278] = (t[310] & ~t[311]);
  assign t[279] = (t[312] & ~t[313]);
  assign t[27] = t[42] ^ t[43];
  assign t[280] = (t[314] & ~t[315]);
  assign t[281] = (t[316] & ~t[317]);
  assign t[282] = (t[318] & ~t[319]);
  assign t[283] = (t[320] & ~t[321]);
  assign t[284] = (t[322] & ~t[323]);
  assign t[285] = (t[324] & ~t[325]);
  assign t[286] = (t[326] & ~t[327]);
  assign t[287] = (t[328] & ~t[329]);
  assign t[288] = (t[330] & ~t[331]);
  assign t[289] = (t[332] & ~t[333]);
  assign t[28] = ~(t[44] ^ t[25]);
  assign t[290] = (t[334] & ~t[335]);
  assign t[291] = (t[336] & ~t[337]);
  assign t[292] = (t[338] & ~t[339]);
  assign t[293] = (t[340] & ~t[341]);
  assign t[294] = (t[342] & ~t[343]);
  assign t[295] = (t[344] & ~t[345]);
  assign t[296] = (t[346] & ~t[347]);
  assign t[297] = (t[348] & ~t[349]);
  assign t[298] = (t[350] & ~t[351]);
  assign t[299] = (t[352] & ~t[353]);
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[4];
  assign t[301] = t[355] ^ x[3];
  assign t[302] = t[356] ^ x[7];
  assign t[303] = t[357] ^ x[6];
  assign t[304] = t[358] ^ x[10];
  assign t[305] = t[359] ^ x[9];
  assign t[306] = t[360] ^ x[13];
  assign t[307] = t[361] ^ x[12];
  assign t[308] = t[362] ^ x[18];
  assign t[309] = t[363] ^ x[17];
  assign t[30] = ~(t[36] ^ t[47]);
  assign t[310] = t[364] ^ x[21];
  assign t[311] = t[365] ^ x[20];
  assign t[312] = t[366] ^ x[24];
  assign t[313] = t[367] ^ x[23];
  assign t[314] = t[368] ^ x[27];
  assign t[315] = t[369] ^ x[26];
  assign t[316] = t[370] ^ x[30];
  assign t[317] = t[371] ^ x[29];
  assign t[318] = t[372] ^ x[33];
  assign t[319] = t[373] ^ x[32];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[36];
  assign t[321] = t[375] ^ x[35];
  assign t[322] = t[376] ^ x[39];
  assign t[323] = t[377] ^ x[38];
  assign t[324] = t[378] ^ x[44];
  assign t[325] = t[379] ^ x[43];
  assign t[326] = t[380] ^ x[47];
  assign t[327] = t[381] ^ x[46];
  assign t[328] = t[382] ^ x[50];
  assign t[329] = t[383] ^ x[49];
  assign t[32] = ~(t[50]);
  assign t[330] = t[384] ^ x[53];
  assign t[331] = t[385] ^ x[52];
  assign t[332] = t[386] ^ x[56];
  assign t[333] = t[387] ^ x[55];
  assign t[334] = t[388] ^ x[59];
  assign t[335] = t[389] ^ x[58];
  assign t[336] = t[390] ^ x[62];
  assign t[337] = t[391] ^ x[61];
  assign t[338] = t[392] ^ x[65];
  assign t[339] = t[393] ^ x[64];
  assign t[33] = ~(t[225]);
  assign t[340] = t[394] ^ x[68];
  assign t[341] = t[395] ^ x[67];
  assign t[342] = t[396] ^ x[73];
  assign t[343] = t[397] ^ x[72];
  assign t[344] = t[398] ^ x[82];
  assign t[345] = t[399] ^ x[81];
  assign t[346] = t[400] ^ x[87];
  assign t[347] = t[401] ^ x[86];
  assign t[348] = t[402] ^ x[96];
  assign t[349] = t[403] ^ x[95];
  assign t[34] = t[51] ^ t[18];
  assign t[350] = t[404] ^ x[103];
  assign t[351] = t[405] ^ x[102];
  assign t[352] = t[406] ^ x[106];
  assign t[353] = t[407] ^ x[105];
  assign t[354] = (x[2]);
  assign t[355] = (x[2]);
  assign t[356] = (x[5]);
  assign t[357] = (x[5]);
  assign t[358] = (x[8]);
  assign t[359] = (x[8]);
  assign t[35] = ~(t[52] ^ t[44]);
  assign t[360] = (x[11]);
  assign t[361] = (x[11]);
  assign t[362] = (x[16]);
  assign t[363] = (x[16]);
  assign t[364] = (x[19]);
  assign t[365] = (x[19]);
  assign t[366] = (x[22]);
  assign t[367] = (x[22]);
  assign t[368] = (x[25]);
  assign t[369] = (x[25]);
  assign t[36] = t[53] ^ t[54];
  assign t[370] = (x[28]);
  assign t[371] = (x[28]);
  assign t[372] = (x[31]);
  assign t[373] = (x[31]);
  assign t[374] = (x[34]);
  assign t[375] = (x[34]);
  assign t[376] = (x[37]);
  assign t[377] = (x[37]);
  assign t[378] = (x[42]);
  assign t[379] = (x[42]);
  assign t[37] = ~(t[55] ^ t[56]);
  assign t[380] = (x[45]);
  assign t[381] = (x[45]);
  assign t[382] = (x[48]);
  assign t[383] = (x[48]);
  assign t[384] = (x[51]);
  assign t[385] = (x[51]);
  assign t[386] = (x[54]);
  assign t[387] = (x[54]);
  assign t[388] = (x[57]);
  assign t[389] = (x[57]);
  assign t[38] = t[9] ? t[57] : t[226];
  assign t[390] = (x[60]);
  assign t[391] = (x[60]);
  assign t[392] = (x[63]);
  assign t[393] = (x[63]);
  assign t[394] = (x[66]);
  assign t[395] = (x[66]);
  assign t[396] = (x[71]);
  assign t[397] = (x[71]);
  assign t[398] = (x[80]);
  assign t[399] = (x[80]);
  assign t[39] = t[58] ^ t[59];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[400] = (x[85]);
  assign t[401] = (x[85]);
  assign t[402] = (x[94]);
  assign t[403] = (x[94]);
  assign t[404] = (x[101]);
  assign t[405] = (x[101]);
  assign t[406] = (x[104]);
  assign t[407] = (x[104]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[42] ^ t[47]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] ^ t[36]);
  assign t[45] = ~(t[67] ^ t[68]);
  assign t[46] = t[69] ^ t[70];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[227] | t[75];
  assign t[4] = t[9] ? t[10] : t[219];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] ^ t[38];
  assign t[54] = t[58] ^ t[82];
  assign t[55] = t[83] ^ t[45];
  assign t[56] = ~(t[25] ^ t[84]);
  assign t[57] = t[226] ^ t[85];
  assign t[58] = t[86] ^ t[78];
  assign t[59] = t[87] & t[88];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[25] ^ t[51];
  assign t[61] = ~(t[89] ^ t[90]);
  assign t[62] = t[91] ^ t[71];
  assign t[63] = t[92] & t[93];
  assign t[64] = t[94] ^ t[95];
  assign t[65] = t[96] ^ t[97];
  assign t[66] = ~(t[98] ^ t[99]);
  assign t[67] = t[100] ^ t[101];
  assign t[68] = ~(t[102] ^ t[103]);
  assign t[69] = t[104] ^ t[94];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[105] & t[106];
  assign t[71] = t[9] ? t[107] : t[228];
  assign t[72] = t[108] ^ t[109];
  assign t[73] = ~(t[75] & t[110]);
  assign t[74] = ~(t[229] ^ t[111]);
  assign t[75] = ~(t[112] & t[113]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[114] ^ t[38];
  assign t[78] = t[115] & t[116];
  assign t[79] = t[117] ^ t[71];
  assign t[7] = ~(t[15] ^ t[16]);
  assign t[80] = t[108] ^ t[118];
  assign t[81] = t[9] ? t[119] : t[230];
  assign t[82] = t[120] & t[121];
  assign t[83] = ~(t[122] ^ t[123]);
  assign t[84] = t[124] ^ t[109];
  assign t[85] = t[125] ? x[41] : x[40];
  assign t[86] = t[126] & t[127];
  assign t[87] = ~(t[128] ^ t[58]);
  assign t[88] = t[53] ^ t[116];
  assign t[89] = ~(t[46] ^ t[103]);
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[9] ? t[131] : t[231];
  assign t[92] = ~(t[117]);
  assign t[93] = t[9] ? t[132] : t[232];
  assign t[94] = t[222] ^ t[133];
  assign t[95] = t[223] ^ t[134];
  assign t[96] = t[135] ^ t[136];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[52] ^ t[139];
  assign t[99] = t[140] ^ t[141];
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [116:0] x;
 output y;

 wire [407:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[142] ^ t[143];
  assign t[101] = t[128] ^ t[59];
  assign t[102] = t[43] ^ t[84];
  assign t[103] = t[144] ^ t[145];
  assign t[104] = t[31] ? t[146] : t[233];
  assign t[105] = ~(t[69] ^ t[96]);
  assign t[106] = t[64] ^ t[147];
  assign t[107] = t[228] ^ t[148];
  assign t[108] = t[149] ^ t[63];
  assign t[109] = t[150] & t[151];
  assign t[10] = t[219] ^ t[20];
  assign t[110] = ~(t[152] & t[153]);
  assign t[111] = t[154] ^ t[234];
  assign t[112] = ~(t[229]);
  assign t[113] = t[155] & t[154];
  assign t[114] = t[9] ? t[156] : t[235];
  assign t[115] = ~(t[81]);
  assign t[116] = t[9] ? t[157] : t[236];
  assign t[117] = t[9] ? t[158] : t[237];
  assign t[118] = t[159] & t[160];
  assign t[119] = t[230] ^ t[161];
  assign t[11] = ~(t[220]);
  assign t[120] = ~(t[86] ^ t[162]);
  assign t[121] = t[77] ^ t[163];
  assign t[122] = t[26] ^ t[164];
  assign t[123] = ~(t[98] ^ t[101]);
  assign t[124] = t[91] ^ t[117];
  assign t[125] = ~(t[50]);
  assign t[126] = ~(t[163]);
  assign t[127] = ~(t[114]);
  assign t[128] = t[114] ^ t[81];
  assign t[129] = t[165] ^ t[144];
  assign t[12] = ~(t[221]);
  assign t[130] = t[166] ^ t[167];
  assign t[131] = t[231] ^ t[168];
  assign t[132] = t[232] ^ t[169];
  assign t[133] = t[31] ? t[170] : t[238];
  assign t[134] = t[171] ? t[172] : t[239];
  assign t[135] = t[173] & t[174];
  assign t[136] = t[175] & t[147];
  assign t[137] = ~(t[135] ^ t[176]);
  assign t[138] = t[177] ^ t[178];
  assign t[139] = t[95] ^ t[179];
  assign t[13] = ~(t[222]);
  assign t[140] = t[180] ^ t[165];
  assign t[141] = t[181] & t[182];
  assign t[142] = t[180] ^ t[144];
  assign t[143] = t[183] & t[184];
  assign t[144] = t[185];
  assign t[145] = t[166] ^ t[141];
  assign t[146] = t[233] ^ t[186];
  assign t[147] = t[225] ^ t[187];
  assign t[148] = t[32] ? x[70] : x[69];
  assign t[149] = t[188] & t[189];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = ~(t[124] ^ t[108]);
  assign t[151] = t[79] ^ t[93];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[190] | t[112]);
  assign t[154] = ~(t[240]);
  assign t[155] = ~(t[234]);
  assign t[156] = t[235] ^ t[191];
  assign t[157] = t[236] ^ t[192];
  assign t[158] = t[237] ^ t[193];
  assign t[159] = ~(t[149] ^ t[194]);
  assign t[15] = t[23] ^ t[24];
  assign t[160] = t[62] ^ t[195];
  assign t[161] = t[125] ? x[75] : x[74];
  assign t[162] = t[53] ^ t[114];
  assign t[163] = t[116] ^ t[81];
  assign t[164] = t[177] ^ t[136];
  assign t[165] = t[196];
  assign t[166] = t[197] ^ t[143];
  assign t[167] = t[198] & t[199];
  assign t[168] = t[32] ? x[77] : x[76];
  assign t[169] = t[32] ? x[79] : x[78];
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = t[238] ^ t[200];
  assign t[171] = ~(t[19]);
  assign t[172] = t[239] ^ t[201];
  assign t[173] = ~(t[178]);
  assign t[174] = ~(t[104]);
  assign t[175] = ~(t[94]);
  assign t[176] = t[64] ^ t[104];
  assign t[177] = t[104] ^ t[95];
  assign t[178] = t[147] ^ t[94];
  assign t[179] = t[96] ^ t[70];
  assign t[17] = ~(t[27] ^ t[28]);
  assign t[180] = ~t[202];
  assign t[181] = ~(t[140] ^ t[166]);
  assign t[182] = t[129] ^ t[184];
  assign t[183] = ~(t[165]);
  assign t[184] = t[203];
  assign t[185] = t[31] ? t[204] : t[241];
  assign t[186] = t[125] ? x[84] : x[83];
  assign t[187] = t[31] ? t[205] : t[242];
  assign t[188] = ~(t[195]);
  assign t[189] = ~(t[91]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[190] = ~(t[227]);
  assign t[191] = t[125] ? x[89] : x[88];
  assign t[192] = t[125] ? x[91] : x[90];
  assign t[193] = t[32] ? x[93] : x[92];
  assign t[194] = t[79] ^ t[91];
  assign t[195] = t[93] ^ t[117];
  assign t[196] = t[31] ? t[206] : t[243];
  assign t[197] = t[207] & t[208];
  assign t[198] = ~(t[197] ^ t[209]);
  assign t[199] = t[142] ^ t[210];
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[125] ? x[98] : x[97];
  assign t[201] = t[211] ? x[100] : x[99];
  assign t[202] = t[31] ? t[212] : t[244];
  assign t[203] = t[31] ? t[213] : t[245];
  assign t[204] = t[241] ^ t[214];
  assign t[205] = t[242] ^ t[215];
  assign t[206] = t[243] ^ t[216];
  assign t[207] = ~(t[210]);
  assign t[208] = ~(t[180]);
  assign t[209] = t[129] ^ t[180];
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = t[184] ^ t[165];
  assign t[211] = ~(t[50]);
  assign t[212] = t[244] ^ t[217];
  assign t[213] = t[245] ^ t[218];
  assign t[214] = t[76] ? x[108] : x[107];
  assign t[215] = t[76] ? x[110] : x[109];
  assign t[216] = t[211] ? x[112] : x[111];
  assign t[217] = t[76] ? x[114] : x[113];
  assign t[218] = t[211] ? x[116] : x[115];
  assign t[219] = (t[246]);
  assign t[21] = ~(t[223]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[33] & t[224]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = (t[266]);
  assign t[23] = ~(t[34] ^ t[35]);
  assign t[240] = (t[267]);
  assign t[241] = (t[268]);
  assign t[242] = (t[269]);
  assign t[243] = (t[270]);
  assign t[244] = (t[271]);
  assign t[245] = (t[272]);
  assign t[246] = t[273] ^ x[4];
  assign t[247] = t[274] ^ x[7];
  assign t[248] = t[275] ^ x[10];
  assign t[249] = t[276] ^ x[13];
  assign t[24] = t[36] ^ t[37];
  assign t[250] = t[277] ^ x[18];
  assign t[251] = t[278] ^ x[21];
  assign t[252] = t[279] ^ x[24];
  assign t[253] = t[280] ^ x[27];
  assign t[254] = t[281] ^ x[30];
  assign t[255] = t[282] ^ x[33];
  assign t[256] = t[283] ^ x[36];
  assign t[257] = t[284] ^ x[39];
  assign t[258] = t[285] ^ x[44];
  assign t[259] = t[286] ^ x[47];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[287] ^ x[50];
  assign t[261] = t[288] ^ x[53];
  assign t[262] = t[289] ^ x[56];
  assign t[263] = t[290] ^ x[59];
  assign t[264] = t[291] ^ x[62];
  assign t[265] = t[292] ^ x[65];
  assign t[266] = t[293] ^ x[68];
  assign t[267] = t[294] ^ x[73];
  assign t[268] = t[295] ^ x[82];
  assign t[269] = t[296] ^ x[87];
  assign t[26] = ~(t[40] ^ t[41]);
  assign t[270] = t[297] ^ x[96];
  assign t[271] = t[298] ^ x[103];
  assign t[272] = t[299] ^ x[106];
  assign t[273] = (t[300] & ~t[301]);
  assign t[274] = (t[302] & ~t[303]);
  assign t[275] = (t[304] & ~t[305]);
  assign t[276] = (t[306] & ~t[307]);
  assign t[277] = (t[308] & ~t[309]);
  assign t[278] = (t[310] & ~t[311]);
  assign t[279] = (t[312] & ~t[313]);
  assign t[27] = t[42] ^ t[43];
  assign t[280] = (t[314] & ~t[315]);
  assign t[281] = (t[316] & ~t[317]);
  assign t[282] = (t[318] & ~t[319]);
  assign t[283] = (t[320] & ~t[321]);
  assign t[284] = (t[322] & ~t[323]);
  assign t[285] = (t[324] & ~t[325]);
  assign t[286] = (t[326] & ~t[327]);
  assign t[287] = (t[328] & ~t[329]);
  assign t[288] = (t[330] & ~t[331]);
  assign t[289] = (t[332] & ~t[333]);
  assign t[28] = ~(t[44] ^ t[25]);
  assign t[290] = (t[334] & ~t[335]);
  assign t[291] = (t[336] & ~t[337]);
  assign t[292] = (t[338] & ~t[339]);
  assign t[293] = (t[340] & ~t[341]);
  assign t[294] = (t[342] & ~t[343]);
  assign t[295] = (t[344] & ~t[345]);
  assign t[296] = (t[346] & ~t[347]);
  assign t[297] = (t[348] & ~t[349]);
  assign t[298] = (t[350] & ~t[351]);
  assign t[299] = (t[352] & ~t[353]);
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[4];
  assign t[301] = t[355] ^ x[3];
  assign t[302] = t[356] ^ x[7];
  assign t[303] = t[357] ^ x[6];
  assign t[304] = t[358] ^ x[10];
  assign t[305] = t[359] ^ x[9];
  assign t[306] = t[360] ^ x[13];
  assign t[307] = t[361] ^ x[12];
  assign t[308] = t[362] ^ x[18];
  assign t[309] = t[363] ^ x[17];
  assign t[30] = ~(t[36] ^ t[47]);
  assign t[310] = t[364] ^ x[21];
  assign t[311] = t[365] ^ x[20];
  assign t[312] = t[366] ^ x[24];
  assign t[313] = t[367] ^ x[23];
  assign t[314] = t[368] ^ x[27];
  assign t[315] = t[369] ^ x[26];
  assign t[316] = t[370] ^ x[30];
  assign t[317] = t[371] ^ x[29];
  assign t[318] = t[372] ^ x[33];
  assign t[319] = t[373] ^ x[32];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[36];
  assign t[321] = t[375] ^ x[35];
  assign t[322] = t[376] ^ x[39];
  assign t[323] = t[377] ^ x[38];
  assign t[324] = t[378] ^ x[44];
  assign t[325] = t[379] ^ x[43];
  assign t[326] = t[380] ^ x[47];
  assign t[327] = t[381] ^ x[46];
  assign t[328] = t[382] ^ x[50];
  assign t[329] = t[383] ^ x[49];
  assign t[32] = ~(t[50]);
  assign t[330] = t[384] ^ x[53];
  assign t[331] = t[385] ^ x[52];
  assign t[332] = t[386] ^ x[56];
  assign t[333] = t[387] ^ x[55];
  assign t[334] = t[388] ^ x[59];
  assign t[335] = t[389] ^ x[58];
  assign t[336] = t[390] ^ x[62];
  assign t[337] = t[391] ^ x[61];
  assign t[338] = t[392] ^ x[65];
  assign t[339] = t[393] ^ x[64];
  assign t[33] = ~(t[225]);
  assign t[340] = t[394] ^ x[68];
  assign t[341] = t[395] ^ x[67];
  assign t[342] = t[396] ^ x[73];
  assign t[343] = t[397] ^ x[72];
  assign t[344] = t[398] ^ x[82];
  assign t[345] = t[399] ^ x[81];
  assign t[346] = t[400] ^ x[87];
  assign t[347] = t[401] ^ x[86];
  assign t[348] = t[402] ^ x[96];
  assign t[349] = t[403] ^ x[95];
  assign t[34] = t[51] ^ t[18];
  assign t[350] = t[404] ^ x[103];
  assign t[351] = t[405] ^ x[102];
  assign t[352] = t[406] ^ x[106];
  assign t[353] = t[407] ^ x[105];
  assign t[354] = (x[2]);
  assign t[355] = (x[2]);
  assign t[356] = (x[5]);
  assign t[357] = (x[5]);
  assign t[358] = (x[8]);
  assign t[359] = (x[8]);
  assign t[35] = ~(t[52] ^ t[44]);
  assign t[360] = (x[11]);
  assign t[361] = (x[11]);
  assign t[362] = (x[16]);
  assign t[363] = (x[16]);
  assign t[364] = (x[19]);
  assign t[365] = (x[19]);
  assign t[366] = (x[22]);
  assign t[367] = (x[22]);
  assign t[368] = (x[25]);
  assign t[369] = (x[25]);
  assign t[36] = t[53] ^ t[54];
  assign t[370] = (x[28]);
  assign t[371] = (x[28]);
  assign t[372] = (x[31]);
  assign t[373] = (x[31]);
  assign t[374] = (x[34]);
  assign t[375] = (x[34]);
  assign t[376] = (x[37]);
  assign t[377] = (x[37]);
  assign t[378] = (x[42]);
  assign t[379] = (x[42]);
  assign t[37] = ~(t[55] ^ t[56]);
  assign t[380] = (x[45]);
  assign t[381] = (x[45]);
  assign t[382] = (x[48]);
  assign t[383] = (x[48]);
  assign t[384] = (x[51]);
  assign t[385] = (x[51]);
  assign t[386] = (x[54]);
  assign t[387] = (x[54]);
  assign t[388] = (x[57]);
  assign t[389] = (x[57]);
  assign t[38] = t[9] ? t[57] : t[226];
  assign t[390] = (x[60]);
  assign t[391] = (x[60]);
  assign t[392] = (x[63]);
  assign t[393] = (x[63]);
  assign t[394] = (x[66]);
  assign t[395] = (x[66]);
  assign t[396] = (x[71]);
  assign t[397] = (x[71]);
  assign t[398] = (x[80]);
  assign t[399] = (x[80]);
  assign t[39] = t[58] ^ t[59];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[400] = (x[85]);
  assign t[401] = (x[85]);
  assign t[402] = (x[94]);
  assign t[403] = (x[94]);
  assign t[404] = (x[101]);
  assign t[405] = (x[101]);
  assign t[406] = (x[104]);
  assign t[407] = (x[104]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[42] ^ t[47]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] ^ t[36]);
  assign t[45] = ~(t[67] ^ t[68]);
  assign t[46] = t[69] ^ t[70];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[227] | t[75];
  assign t[4] = t[9] ? t[10] : t[219];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] ^ t[38];
  assign t[54] = t[58] ^ t[82];
  assign t[55] = t[83] ^ t[45];
  assign t[56] = ~(t[25] ^ t[84]);
  assign t[57] = t[226] ^ t[85];
  assign t[58] = t[86] ^ t[78];
  assign t[59] = t[87] & t[88];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[25] ^ t[51];
  assign t[61] = ~(t[89] ^ t[90]);
  assign t[62] = t[91] ^ t[71];
  assign t[63] = t[92] & t[93];
  assign t[64] = t[94] ^ t[95];
  assign t[65] = t[96] ^ t[97];
  assign t[66] = ~(t[98] ^ t[99]);
  assign t[67] = t[100] ^ t[101];
  assign t[68] = ~(t[102] ^ t[103]);
  assign t[69] = t[104] ^ t[94];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[105] & t[106];
  assign t[71] = t[9] ? t[107] : t[228];
  assign t[72] = t[108] ^ t[109];
  assign t[73] = ~(t[75] & t[110]);
  assign t[74] = ~(t[229] ^ t[111]);
  assign t[75] = ~(t[112] & t[113]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[114] ^ t[38];
  assign t[78] = t[115] & t[116];
  assign t[79] = t[117] ^ t[71];
  assign t[7] = ~(t[15] ^ t[16]);
  assign t[80] = t[108] ^ t[118];
  assign t[81] = t[9] ? t[119] : t[230];
  assign t[82] = t[120] & t[121];
  assign t[83] = ~(t[122] ^ t[123]);
  assign t[84] = t[124] ^ t[109];
  assign t[85] = t[125] ? x[41] : x[40];
  assign t[86] = t[126] & t[127];
  assign t[87] = ~(t[128] ^ t[58]);
  assign t[88] = t[53] ^ t[116];
  assign t[89] = ~(t[46] ^ t[103]);
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[9] ? t[131] : t[231];
  assign t[92] = ~(t[117]);
  assign t[93] = t[9] ? t[132] : t[232];
  assign t[94] = t[222] ^ t[133];
  assign t[95] = t[223] ^ t[134];
  assign t[96] = t[135] ^ t[136];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[52] ^ t[139];
  assign t[99] = t[140] ^ t[141];
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[85] ^ t[111];
  assign t[101] = t[120] ^ t[138];
  assign t[102] = t[139] ^ t[140];
  assign t[103] = t[141] ^ t[134];
  assign t[104] = t[107] ? t[142] : t[226];
  assign t[105] = t[143] ^ t[110];
  assign t[106] = t[144] & t[145];
  assign t[107] = ~(t[146]);
  assign t[108] = t[220] ^ t[147];
  assign t[109] = t[124] ^ t[71];
  assign t[10] = t[210] ^ t[21];
  assign t[110] = t[148] & t[149];
  assign t[111] = t[107] ? t[150] : t[227];
  assign t[112] = t[120] ^ t[58];
  assign t[113] = t[151] ^ t[122];
  assign t[114] = ~(t[214]);
  assign t[115] = t[9] ? t[152] : t[228];
  assign t[116] = t[153];
  assign t[117] = t[9] ? t[154] : t[229];
  assign t[118] = t[222] ^ t[155];
  assign t[119] = t[223] ^ t[156];
  assign t[11] = ~(t[211]);
  assign t[120] = t[157] ^ t[158];
  assign t[121] = t[107] ? t[159] : t[230];
  assign t[122] = t[213] ^ t[160];
  assign t[123] = t[161] & t[162];
  assign t[124] = t[107] ? t[163] : t[231];
  assign t[125] = ~(t[90] ^ t[105]);
  assign t[126] = t[69] ^ t[149];
  assign t[127] = t[224] ^ t[164];
  assign t[128] = t[165] & t[166];
  assign t[129] = ~(t[137] ^ t[93]);
  assign t[12] = ~(t[212]);
  assign t[130] = t[139] ^ t[83];
  assign t[131] = ~(t[146]);
  assign t[132] = t[225] ^ t[167];
  assign t[133] = t[168] & t[169];
  assign t[134] = t[170] & t[171];
  assign t[135] = ~(t[113] ^ t[96]);
  assign t[136] = t[88] ^ t[171];
  assign t[137] = t[81] ^ t[116];
  assign t[138] = t[172] & t[173];
  assign t[139] = t[116] ^ t[61];
  assign t[13] = ~(t[213]);
  assign t[140] = t[93] ^ t[174];
  assign t[141] = t[151] ^ t[63];
  assign t[142] = t[226] ^ t[175];
  assign t[143] = t[176] & t[177];
  assign t[144] = ~(t[143] ^ t[178]);
  assign t[145] = t[109] ^ t[179];
  assign t[146] = ~(t[9]);
  assign t[147] = t[35] ? x[71] : x[70];
  assign t[148] = ~(t[104]);
  assign t[149] = t[107] ? t[180] : t[232];
  assign t[14] = ~(t[22] | t[23]);
  assign t[150] = t[227] ^ t[181];
  assign t[151] = t[9] ? t[182] : t[233];
  assign t[152] = t[228] ^ t[183];
  assign t[153] = t[9] ? t[184] : t[234];
  assign t[154] = t[229] ^ t[185];
  assign t[155] = t[186] ? x[82] : x[81];
  assign t[156] = t[186] ? x[84] : x[83];
  assign t[157] = t[187] & t[188];
  assign t[158] = t[189] & t[121];
  assign t[159] = t[230] ^ t[190];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = t[9] ? t[191] : t[235];
  assign t[161] = ~(t[133] ^ t[192]);
  assign t[162] = t[141] ^ t[193];
  assign t[163] = t[231] ^ t[194];
  assign t[164] = t[80] ? x[89] : x[88];
  assign t[165] = ~(t[195]);
  assign t[166] = ~(t[81]);
  assign t[167] = t[196] ? x[91] : x[90];
  assign t[168] = ~(t[193]);
  assign t[169] = ~(t[151]);
  assign t[16] = ~(t[26] ^ t[27]);
  assign t[170] = ~(t[122]);
  assign t[171] = t[218] ^ t[197];
  assign t[172] = ~(t[157] ^ t[198]);
  assign t[173] = t[199] ^ t[200];
  assign t[174] = t[201] & t[202];
  assign t[175] = t[35] ? x[93] : x[92];
  assign t[176] = ~(t[179]);
  assign t[177] = ~(t[124]);
  assign t[178] = t[69] ^ t[124];
  assign t[179] = t[149] ^ t[104];
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[180] = t[232] ^ t[203];
  assign t[181] = t[186] ? x[95] : x[94];
  assign t[182] = t[233] ^ t[204];
  assign t[183] = t[80] ? x[97] : x[96];
  assign t[184] = t[234] ^ t[205];
  assign t[185] = t[196] ? x[99] : x[98];
  assign t[186] = ~(t[54]);
  assign t[187] = ~(t[200]);
  assign t[188] = ~(t[84]);
  assign t[189] = ~(t[85]);
  assign t[18] = ~(t[30] ^ t[31]);
  assign t[190] = t[186] ? x[101] : x[100];
  assign t[191] = t[235] ^ t[206];
  assign t[192] = t[88] ^ t[151];
  assign t[193] = t[171] ^ t[122];
  assign t[194] = t[35] ? x[103] : x[102];
  assign t[195] = t[83] ^ t[116];
  assign t[196] = ~(t[54]);
  assign t[197] = t[9] ? t[207] : t[236];
  assign t[198] = t[100] ^ t[84];
  assign t[199] = t[84] ^ t[111];
  assign t[19] = ~(t[32] & t[33]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[121] ^ t[85];
  assign t[201] = ~(t[128] ^ t[208]);
  assign t[202] = t[55] ^ t[195];
  assign t[203] = t[35] ? x[108] : x[107];
  assign t[204] = t[186] ? x[110] : x[109];
  assign t[205] = t[196] ? x[112] : x[111];
  assign t[206] = t[186] ? x[114] : x[113];
  assign t[207] = t[236] ^ t[209];
  assign t[208] = t[139] ^ t[81];
  assign t[209] = t[80] ? x[116] : x[115];
  assign t[20] = t[214] | t[34];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[35] ? x[18] : x[17];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[215]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[7];
  assign t[239] = t[266] ^ x[10];
  assign t[23] = ~(t[36] & t[216]);
  assign t[240] = t[267] ^ x[13];
  assign t[241] = t[268] ^ x[16];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = t[37] ^ t[38];
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[51];
  assign t[253] = t[280] ^ x[54];
  assign t[254] = t[281] ^ x[57];
  assign t[255] = t[282] ^ x[60];
  assign t[256] = t[283] ^ x[63];
  assign t[257] = t[284] ^ x[66];
  assign t[258] = t[285] ^ x[69];
  assign t[259] = t[286] ^ x[74];
  assign t[25] = ~(t[39] ^ t[40]);
  assign t[260] = t[287] ^ x[77];
  assign t[261] = t[288] ^ x[80];
  assign t[262] = t[289] ^ x[87];
  assign t[263] = t[290] ^ x[106];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = ~(t[41] ^ t[39]);
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = t[42] ^ t[43];
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = t[27] ^ t[38];
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[7];
  assign t[294] = t[348] ^ x[6];
  assign t[295] = t[349] ^ x[10];
  assign t[296] = t[350] ^ x[9];
  assign t[297] = t[351] ^ x[13];
  assign t[298] = t[352] ^ x[12];
  assign t[299] = t[353] ^ x[16];
  assign t[29] = ~(t[44] ^ t[45]);
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[15];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = ~(t[46] ^ t[47]);
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[48] ^ t[49]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[51];
  assign t[322] = t[376] ^ x[50];
  assign t[323] = t[377] ^ x[54];
  assign t[324] = t[378] ^ x[53];
  assign t[325] = t[379] ^ x[57];
  assign t[326] = t[380] ^ x[56];
  assign t[327] = t[381] ^ x[60];
  assign t[328] = t[382] ^ x[59];
  assign t[329] = t[383] ^ x[63];
  assign t[32] = ~(t[34] & t[50]);
  assign t[330] = t[384] ^ x[62];
  assign t[331] = t[385] ^ x[66];
  assign t[332] = t[386] ^ x[65];
  assign t[333] = t[387] ^ x[69];
  assign t[334] = t[388] ^ x[68];
  assign t[335] = t[389] ^ x[74];
  assign t[336] = t[390] ^ x[73];
  assign t[337] = t[391] ^ x[77];
  assign t[338] = t[392] ^ x[76];
  assign t[339] = t[393] ^ x[80];
  assign t[33] = ~(t[217] ^ t[51]);
  assign t[340] = t[394] ^ x[79];
  assign t[341] = t[395] ^ x[87];
  assign t[342] = t[396] ^ x[86];
  assign t[343] = t[397] ^ x[106];
  assign t[344] = t[398] ^ x[105];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[5]);
  assign t[348] = (x[5]);
  assign t[349] = (x[8]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[8]);
  assign t[351] = (x[11]);
  assign t[352] = (x[11]);
  assign t[353] = (x[14]);
  assign t[354] = (x[14]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = ~(t[54]);
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = ~(t[218]);
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[49]);
  assign t[376] = (x[49]);
  assign t[377] = (x[52]);
  assign t[378] = (x[52]);
  assign t[379] = (x[55]);
  assign t[37] = t[55] ^ t[56];
  assign t[380] = (x[55]);
  assign t[381] = (x[58]);
  assign t[382] = (x[58]);
  assign t[383] = (x[61]);
  assign t[384] = (x[61]);
  assign t[385] = (x[64]);
  assign t[386] = (x[64]);
  assign t[387] = (x[67]);
  assign t[388] = (x[67]);
  assign t[389] = (x[72]);
  assign t[38] = t[57] ^ t[58];
  assign t[390] = (x[72]);
  assign t[391] = (x[75]);
  assign t[392] = (x[75]);
  assign t[393] = (x[78]);
  assign t[394] = (x[78]);
  assign t[395] = (x[85]);
  assign t[396] = (x[85]);
  assign t[397] = (x[104]);
  assign t[398] = (x[104]);
  assign t[39] = t[59] ^ t[60];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = ~(t[65] ^ t[66]);
  assign t[43] = ~(t[67] ^ t[68]);
  assign t[44] = t[69] ^ t[70];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = t[73] ^ t[59];
  assign t[47] = ~(t[42] ^ t[74]);
  assign t[48] = t[15] ^ t[75];
  assign t[49] = ~(t[66] ^ t[45]);
  assign t[4] = t[9] ? t[10] : t[210];
  assign t[50] = ~(t[76] & t[77]);
  assign t[51] = t[78] ^ t[219];
  assign t[52] = ~(t[217]);
  assign t[53] = t[79] & t[78];
  assign t[54] = ~(t[80]);
  assign t[55] = t[81] ^ t[61];
  assign t[56] = t[82] & t[83];
  assign t[57] = t[84] ^ t[85];
  assign t[58] = t[86] & t[87];
  assign t[59] = t[88] ^ t[89];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92];
  assign t[62] = t[93] ^ t[94];
  assign t[63] = t[215] ^ t[95];
  assign t[64] = t[96] ^ t[97];
  assign t[65] = ~(t[98] ^ t[99]);
  assign t[66] = t[100] ^ t[101];
  assign t[67] = t[102] ^ t[103];
  assign t[68] = ~(t[74] ^ t[45]);
  assign t[69] = t[104] ^ t[71];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[105] ^ t[106];
  assign t[71] = t[107] ? t[108] : t[220];
  assign t[72] = t[105] ^ t[91];
  assign t[73] = t[109] ^ t[110];
  assign t[74] = t[111] ^ t[112];
  assign t[75] = t[113] ^ t[97];
  assign t[76] = ~(t[79] | t[78]);
  assign t[77] = ~(t[114] | t[52]);
  assign t[78] = ~(t[221]);
  assign t[79] = ~(t[219]);
  assign t[7] = ~(t[15] ^ t[16]);
  assign t[80] = ~(t[20]);
  assign t[81] = ~t[115];
  assign t[82] = ~(t[116]);
  assign t[83] = t[117];
  assign t[84] = t[107] ? t[118] : t[222];
  assign t[85] = t[107] ? t[119] : t[223];
  assign t[86] = ~(t[57] ^ t[120]);
  assign t[87] = t[100] ^ t[121];
  assign t[88] = t[122] ^ t[63];
  assign t[89] = t[96] ^ t[123];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = t[124] ^ t[104];
  assign t[91] = t[125] & t[126];
  assign t[92] = t[9] ? t[127] : t[224];
  assign t[93] = t[128] ^ t[56];
  assign t[94] = t[129] & t[130];
  assign t[95] = t[131] ? t[132] : t[225];
  assign t[96] = t[133] ^ t[134];
  assign t[97] = t[135] & t[136];
  assign t[98] = t[44] ^ t[41];
  assign t[99] = t[137] ^ t[94];
  assign t[9] = ~(t[19] & t[20]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[85] ^ t[111];
  assign t[101] = t[120] ^ t[138];
  assign t[102] = t[139] ^ t[140];
  assign t[103] = t[141] ^ t[134];
  assign t[104] = t[107] ? t[142] : t[226];
  assign t[105] = t[143] ^ t[110];
  assign t[106] = t[144] & t[145];
  assign t[107] = ~(t[146]);
  assign t[108] = t[220] ^ t[147];
  assign t[109] = t[124] ^ t[71];
  assign t[10] = t[210] ^ t[21];
  assign t[110] = t[148] & t[149];
  assign t[111] = t[107] ? t[150] : t[227];
  assign t[112] = t[120] ^ t[58];
  assign t[113] = t[151] ^ t[122];
  assign t[114] = ~(t[214]);
  assign t[115] = t[9] ? t[152] : t[228];
  assign t[116] = t[153];
  assign t[117] = t[9] ? t[154] : t[229];
  assign t[118] = t[222] ^ t[155];
  assign t[119] = t[223] ^ t[156];
  assign t[11] = ~(t[211]);
  assign t[120] = t[157] ^ t[158];
  assign t[121] = t[107] ? t[159] : t[230];
  assign t[122] = t[213] ^ t[160];
  assign t[123] = t[161] & t[162];
  assign t[124] = t[107] ? t[163] : t[231];
  assign t[125] = ~(t[90] ^ t[105]);
  assign t[126] = t[69] ^ t[149];
  assign t[127] = t[224] ^ t[164];
  assign t[128] = t[165] & t[166];
  assign t[129] = ~(t[137] ^ t[93]);
  assign t[12] = ~(t[212]);
  assign t[130] = t[139] ^ t[83];
  assign t[131] = ~(t[146]);
  assign t[132] = t[225] ^ t[167];
  assign t[133] = t[168] & t[169];
  assign t[134] = t[170] & t[171];
  assign t[135] = ~(t[113] ^ t[96]);
  assign t[136] = t[88] ^ t[171];
  assign t[137] = t[81] ^ t[116];
  assign t[138] = t[172] & t[173];
  assign t[139] = t[116] ^ t[61];
  assign t[13] = ~(t[213]);
  assign t[140] = t[93] ^ t[174];
  assign t[141] = t[151] ^ t[63];
  assign t[142] = t[226] ^ t[175];
  assign t[143] = t[176] & t[177];
  assign t[144] = ~(t[143] ^ t[178]);
  assign t[145] = t[109] ^ t[179];
  assign t[146] = ~(t[9]);
  assign t[147] = t[35] ? x[71] : x[70];
  assign t[148] = ~(t[104]);
  assign t[149] = t[107] ? t[180] : t[232];
  assign t[14] = ~(t[22] | t[23]);
  assign t[150] = t[227] ^ t[181];
  assign t[151] = t[9] ? t[182] : t[233];
  assign t[152] = t[228] ^ t[183];
  assign t[153] = t[9] ? t[184] : t[234];
  assign t[154] = t[229] ^ t[185];
  assign t[155] = t[186] ? x[82] : x[81];
  assign t[156] = t[186] ? x[84] : x[83];
  assign t[157] = t[187] & t[188];
  assign t[158] = t[189] & t[121];
  assign t[159] = t[230] ^ t[190];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = t[9] ? t[191] : t[235];
  assign t[161] = ~(t[133] ^ t[192]);
  assign t[162] = t[141] ^ t[193];
  assign t[163] = t[231] ^ t[194];
  assign t[164] = t[80] ? x[89] : x[88];
  assign t[165] = ~(t[195]);
  assign t[166] = ~(t[81]);
  assign t[167] = t[196] ? x[91] : x[90];
  assign t[168] = ~(t[193]);
  assign t[169] = ~(t[151]);
  assign t[16] = ~(t[26] ^ t[27]);
  assign t[170] = ~(t[122]);
  assign t[171] = t[218] ^ t[197];
  assign t[172] = ~(t[157] ^ t[198]);
  assign t[173] = t[199] ^ t[200];
  assign t[174] = t[201] & t[202];
  assign t[175] = t[35] ? x[93] : x[92];
  assign t[176] = ~(t[179]);
  assign t[177] = ~(t[124]);
  assign t[178] = t[69] ^ t[124];
  assign t[179] = t[149] ^ t[104];
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[180] = t[232] ^ t[203];
  assign t[181] = t[186] ? x[95] : x[94];
  assign t[182] = t[233] ^ t[204];
  assign t[183] = t[80] ? x[97] : x[96];
  assign t[184] = t[234] ^ t[205];
  assign t[185] = t[196] ? x[99] : x[98];
  assign t[186] = ~(t[54]);
  assign t[187] = ~(t[200]);
  assign t[188] = ~(t[84]);
  assign t[189] = ~(t[85]);
  assign t[18] = ~(t[30] ^ t[31]);
  assign t[190] = t[186] ? x[101] : x[100];
  assign t[191] = t[235] ^ t[206];
  assign t[192] = t[88] ^ t[151];
  assign t[193] = t[171] ^ t[122];
  assign t[194] = t[35] ? x[103] : x[102];
  assign t[195] = t[83] ^ t[116];
  assign t[196] = ~(t[54]);
  assign t[197] = t[9] ? t[207] : t[236];
  assign t[198] = t[100] ^ t[84];
  assign t[199] = t[84] ^ t[111];
  assign t[19] = ~(t[32] & t[33]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[121] ^ t[85];
  assign t[201] = ~(t[128] ^ t[208]);
  assign t[202] = t[55] ^ t[195];
  assign t[203] = t[35] ? x[108] : x[107];
  assign t[204] = t[186] ? x[110] : x[109];
  assign t[205] = t[196] ? x[112] : x[111];
  assign t[206] = t[186] ? x[114] : x[113];
  assign t[207] = t[236] ^ t[209];
  assign t[208] = t[139] ^ t[81];
  assign t[209] = t[80] ? x[116] : x[115];
  assign t[20] = t[214] | t[34];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[35] ? x[18] : x[17];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[215]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[7];
  assign t[239] = t[266] ^ x[10];
  assign t[23] = ~(t[36] & t[216]);
  assign t[240] = t[267] ^ x[13];
  assign t[241] = t[268] ^ x[16];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = t[37] ^ t[38];
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[51];
  assign t[253] = t[280] ^ x[54];
  assign t[254] = t[281] ^ x[57];
  assign t[255] = t[282] ^ x[60];
  assign t[256] = t[283] ^ x[63];
  assign t[257] = t[284] ^ x[66];
  assign t[258] = t[285] ^ x[69];
  assign t[259] = t[286] ^ x[74];
  assign t[25] = ~(t[39] ^ t[40]);
  assign t[260] = t[287] ^ x[77];
  assign t[261] = t[288] ^ x[80];
  assign t[262] = t[289] ^ x[87];
  assign t[263] = t[290] ^ x[106];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = ~(t[41] ^ t[39]);
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = t[42] ^ t[43];
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = t[27] ^ t[38];
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[7];
  assign t[294] = t[348] ^ x[6];
  assign t[295] = t[349] ^ x[10];
  assign t[296] = t[350] ^ x[9];
  assign t[297] = t[351] ^ x[13];
  assign t[298] = t[352] ^ x[12];
  assign t[299] = t[353] ^ x[16];
  assign t[29] = ~(t[44] ^ t[45]);
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[15];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = ~(t[46] ^ t[47]);
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[48] ^ t[49]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[51];
  assign t[322] = t[376] ^ x[50];
  assign t[323] = t[377] ^ x[54];
  assign t[324] = t[378] ^ x[53];
  assign t[325] = t[379] ^ x[57];
  assign t[326] = t[380] ^ x[56];
  assign t[327] = t[381] ^ x[60];
  assign t[328] = t[382] ^ x[59];
  assign t[329] = t[383] ^ x[63];
  assign t[32] = ~(t[34] & t[50]);
  assign t[330] = t[384] ^ x[62];
  assign t[331] = t[385] ^ x[66];
  assign t[332] = t[386] ^ x[65];
  assign t[333] = t[387] ^ x[69];
  assign t[334] = t[388] ^ x[68];
  assign t[335] = t[389] ^ x[74];
  assign t[336] = t[390] ^ x[73];
  assign t[337] = t[391] ^ x[77];
  assign t[338] = t[392] ^ x[76];
  assign t[339] = t[393] ^ x[80];
  assign t[33] = ~(t[217] ^ t[51]);
  assign t[340] = t[394] ^ x[79];
  assign t[341] = t[395] ^ x[87];
  assign t[342] = t[396] ^ x[86];
  assign t[343] = t[397] ^ x[106];
  assign t[344] = t[398] ^ x[105];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[5]);
  assign t[348] = (x[5]);
  assign t[349] = (x[8]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[8]);
  assign t[351] = (x[11]);
  assign t[352] = (x[11]);
  assign t[353] = (x[14]);
  assign t[354] = (x[14]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = ~(t[54]);
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = ~(t[218]);
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[49]);
  assign t[376] = (x[49]);
  assign t[377] = (x[52]);
  assign t[378] = (x[52]);
  assign t[379] = (x[55]);
  assign t[37] = t[55] ^ t[56];
  assign t[380] = (x[55]);
  assign t[381] = (x[58]);
  assign t[382] = (x[58]);
  assign t[383] = (x[61]);
  assign t[384] = (x[61]);
  assign t[385] = (x[64]);
  assign t[386] = (x[64]);
  assign t[387] = (x[67]);
  assign t[388] = (x[67]);
  assign t[389] = (x[72]);
  assign t[38] = t[57] ^ t[58];
  assign t[390] = (x[72]);
  assign t[391] = (x[75]);
  assign t[392] = (x[75]);
  assign t[393] = (x[78]);
  assign t[394] = (x[78]);
  assign t[395] = (x[85]);
  assign t[396] = (x[85]);
  assign t[397] = (x[104]);
  assign t[398] = (x[104]);
  assign t[39] = t[59] ^ t[60];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = ~(t[65] ^ t[66]);
  assign t[43] = ~(t[67] ^ t[68]);
  assign t[44] = t[69] ^ t[70];
  assign t[45] = t[71] ^ t[72];
  assign t[46] = t[73] ^ t[59];
  assign t[47] = ~(t[42] ^ t[74]);
  assign t[48] = t[15] ^ t[75];
  assign t[49] = ~(t[66] ^ t[45]);
  assign t[4] = t[9] ? t[10] : t[210];
  assign t[50] = ~(t[76] & t[77]);
  assign t[51] = t[78] ^ t[219];
  assign t[52] = ~(t[217]);
  assign t[53] = t[79] & t[78];
  assign t[54] = ~(t[80]);
  assign t[55] = t[81] ^ t[61];
  assign t[56] = t[82] & t[83];
  assign t[57] = t[84] ^ t[85];
  assign t[58] = t[86] & t[87];
  assign t[59] = t[88] ^ t[89];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92];
  assign t[62] = t[93] ^ t[94];
  assign t[63] = t[215] ^ t[95];
  assign t[64] = t[96] ^ t[97];
  assign t[65] = ~(t[98] ^ t[99]);
  assign t[66] = t[100] ^ t[101];
  assign t[67] = t[102] ^ t[103];
  assign t[68] = ~(t[74] ^ t[45]);
  assign t[69] = t[104] ^ t[71];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[105] ^ t[106];
  assign t[71] = t[107] ? t[108] : t[220];
  assign t[72] = t[105] ^ t[91];
  assign t[73] = t[109] ^ t[110];
  assign t[74] = t[111] ^ t[112];
  assign t[75] = t[113] ^ t[97];
  assign t[76] = ~(t[79] | t[78]);
  assign t[77] = ~(t[114] | t[52]);
  assign t[78] = ~(t[221]);
  assign t[79] = ~(t[219]);
  assign t[7] = ~(t[15] ^ t[16]);
  assign t[80] = ~(t[20]);
  assign t[81] = ~t[115];
  assign t[82] = ~(t[116]);
  assign t[83] = t[117];
  assign t[84] = t[107] ? t[118] : t[222];
  assign t[85] = t[107] ? t[119] : t[223];
  assign t[86] = ~(t[57] ^ t[120]);
  assign t[87] = t[100] ^ t[121];
  assign t[88] = t[122] ^ t[63];
  assign t[89] = t[96] ^ t[123];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = t[124] ^ t[104];
  assign t[91] = t[125] & t[126];
  assign t[92] = t[9] ? t[127] : t[224];
  assign t[93] = t[128] ^ t[56];
  assign t[94] = t[129] & t[130];
  assign t[95] = t[131] ? t[132] : t[225];
  assign t[96] = t[133] ^ t[134];
  assign t[97] = t[135] & t[136];
  assign t[98] = t[44] ^ t[41];
  assign t[99] = t[137] ^ t[94];
  assign t[9] = ~(t[19] & t[20]);
  assign y = (t[0]);
endmodule

module R2ind126(x, y);
 input [116:0] x;
 output y;

 wire [396:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ? x[49] : x[48];
  assign t[101] = t[219] ^ t[141];
  assign t[102] = ~(t[142] & t[143]);
  assign t[103] = t[144] ^ t[222];
  assign t[104] = ~(t[220]);
  assign t[105] = t[145] & t[144];
  assign t[106] = t[85] ^ t[125];
  assign t[107] = t[146] & t[147];
  assign t[108] = t[148];
  assign t[109] = t[110] ^ t[61];
  assign t[10] = t[208] ^ t[20];
  assign t[110] = t[149] ^ t[150];
  assign t[111] = t[151] & t[152];
  assign t[112] = t[153] ? t[154] : t[223];
  assign t[113] = t[155] ^ t[58];
  assign t[114] = t[125] ^ t[76];
  assign t[115] = t[113] ^ t[156];
  assign t[116] = t[157] ^ t[127];
  assign t[117] = t[158] & t[159];
  assign t[118] = t[62] ^ t[160];
  assign t[119] = t[138] ^ t[96];
  assign t[11] = ~(t[209]);
  assign t[120] = t[157] ^ t[122];
  assign t[121] = t[161] & t[162];
  assign t[122] = t[9] ? t[163] : t[224];
  assign t[123] = t[128] ^ t[117];
  assign t[124] = t[221] ^ t[164];
  assign t[125] = t[211] ^ t[165];
  assign t[126] = t[31] ? t[166] : t[225];
  assign t[127] = t[9] ? t[167] : t[226];
  assign t[128] = t[168] ^ t[121];
  assign t[129] = t[169] & t[170];
  assign t[12] = ~(t[210]);
  assign t[130] = t[31] ? t[171] : t[227];
  assign t[131] = t[31] ? t[172] : t[228];
  assign t[132] = t[173];
  assign t[133] = t[140] ? x[72] : x[71];
  assign t[134] = ~(t[139]);
  assign t[135] = ~(t[43]);
  assign t[136] = ~(t[44]);
  assign t[137] = t[41] ^ t[43];
  assign t[138] = t[43] ^ t[62];
  assign t[139] = t[67] ^ t[44];
  assign t[13] = ~(t[211]);
  assign t[140] = ~(t[49]);
  assign t[141] = t[140] ? x[74] : x[73];
  assign t[142] = ~(t[145] | t[144]);
  assign t[143] = ~(t[174] | t[104]);
  assign t[144] = ~(t[229]);
  assign t[145] = ~(t[222]);
  assign t[146] = ~(t[106] ^ t[113]);
  assign t[147] = t[114] ^ t[87];
  assign t[148] = t[31] ? t[175] : t[230];
  assign t[149] = t[176] & t[177];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = t[178] & t[132];
  assign t[151] = ~(t[149] ^ t[179]);
  assign t[152] = t[180] ^ t[181];
  assign t[153] = ~(t[19]);
  assign t[154] = t[223] ^ t[182];
  assign t[155] = t[183] & t[184];
  assign t[156] = t[185] & t[186];
  assign t[157] = t[9] ? t[187] : t[231];
  assign t[158] = ~(t[116] ^ t[128]);
  assign t[159] = t[88] ^ t[162];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[63] ^ t[30];
  assign t[161] = ~(t[127]);
  assign t[162] = t[9] ? t[188] : t[232];
  assign t[163] = t[224] ^ t[189];
  assign t[164] = t[140] ? x[88] : x[87];
  assign t[165] = t[31] ? t[190] : t[233];
  assign t[166] = t[225] ^ t[191];
  assign t[167] = t[226] ^ t[192];
  assign t[168] = t[193] & t[194];
  assign t[169] = ~(t[168] ^ t[195]);
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = t[120] ^ t[196];
  assign t[171] = t[227] ^ t[197];
  assign t[172] = t[228] ^ t[198];
  assign t[173] = t[31] ? t[199] : t[234];
  assign t[174] = ~(t[217]);
  assign t[175] = t[230] ^ t[200];
  assign t[176] = ~(t[181]);
  assign t[177] = ~(t[90]);
  assign t[178] = ~(t[91]);
  assign t[179] = t[74] ^ t[90];
  assign t[17] = ~(t[27] ^ t[28]);
  assign t[180] = t[90] ^ t[108];
  assign t[181] = t[132] ^ t[91];
  assign t[182] = t[201] ? x[96] : x[95];
  assign t[183] = ~(t[202]);
  assign t[184] = ~(t[85]);
  assign t[185] = ~(t[155] ^ t[203]);
  assign t[186] = t[57] ^ t[202];
  assign t[187] = t[231] ^ t[204];
  assign t[188] = t[232] ^ t[205];
  assign t[189] = t[32] ? x[98] : x[97];
  assign t[18] = t[29] ^ t[30];
  assign t[190] = t[233] ^ t[206];
  assign t[191] = t[71] ? x[100] : x[99];
  assign t[192] = t[32] ? x[102] : x[101];
  assign t[193] = ~(t[196]);
  assign t[194] = ~(t[157]);
  assign t[195] = t[88] ^ t[157];
  assign t[196] = t[162] ^ t[127];
  assign t[197] = t[71] ? x[104] : x[103];
  assign t[198] = t[201] ? x[106] : x[105];
  assign t[199] = t[234] ^ t[207];
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[71] ? x[108] : x[107];
  assign t[201] = ~(t[49]);
  assign t[202] = t[87] ^ t[125];
  assign t[203] = t[114] ^ t[85];
  assign t[204] = t[32] ? x[110] : x[109];
  assign t[205] = t[32] ? x[112] : x[111];
  assign t[206] = t[140] ? x[114] : x[113];
  assign t[207] = t[201] ? x[116] : x[115];
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[212]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[33] & t[213]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = t[262] ^ x[4];
  assign t[236] = t[263] ^ x[7];
  assign t[237] = t[264] ^ x[10];
  assign t[238] = t[265] ^ x[13];
  assign t[239] = t[266] ^ x[18];
  assign t[23] = ~(t[28] ^ t[34]);
  assign t[240] = t[267] ^ x[21];
  assign t[241] = t[268] ^ x[24];
  assign t[242] = t[269] ^ x[27];
  assign t[243] = t[270] ^ x[30];
  assign t[244] = t[271] ^ x[33];
  assign t[245] = t[272] ^ x[36];
  assign t[246] = t[273] ^ x[39];
  assign t[247] = t[274] ^ x[42];
  assign t[248] = t[275] ^ x[45];
  assign t[249] = t[276] ^ x[52];
  assign t[24] = ~(t[35] ^ t[36]);
  assign t[250] = t[277] ^ x[55];
  assign t[251] = t[278] ^ x[58];
  assign t[252] = t[279] ^ x[61];
  assign t[253] = t[280] ^ x[64];
  assign t[254] = t[281] ^ x[67];
  assign t[255] = t[282] ^ x[70];
  assign t[256] = t[283] ^ x[77];
  assign t[257] = t[284] ^ x[80];
  assign t[258] = t[285] ^ x[83];
  assign t[259] = t[286] ^ x[86];
  assign t[25] = t[37] ^ t[38];
  assign t[260] = t[287] ^ x[91];
  assign t[261] = t[288] ^ x[94];
  assign t[262] = (t[289] & ~t[290]);
  assign t[263] = (t[291] & ~t[292]);
  assign t[264] = (t[293] & ~t[294]);
  assign t[265] = (t[295] & ~t[296]);
  assign t[266] = (t[297] & ~t[298]);
  assign t[267] = (t[299] & ~t[300]);
  assign t[268] = (t[301] & ~t[302]);
  assign t[269] = (t[303] & ~t[304]);
  assign t[26] = ~(t[39] ^ t[18]);
  assign t[270] = (t[305] & ~t[306]);
  assign t[271] = (t[307] & ~t[308]);
  assign t[272] = (t[309] & ~t[310]);
  assign t[273] = (t[311] & ~t[312]);
  assign t[274] = (t[313] & ~t[314]);
  assign t[275] = (t[315] & ~t[316]);
  assign t[276] = (t[317] & ~t[318]);
  assign t[277] = (t[319] & ~t[320]);
  assign t[278] = (t[321] & ~t[322]);
  assign t[279] = (t[323] & ~t[324]);
  assign t[27] = ~(t[39] ^ t[40]);
  assign t[280] = (t[325] & ~t[326]);
  assign t[281] = (t[327] & ~t[328]);
  assign t[282] = (t[329] & ~t[330]);
  assign t[283] = (t[331] & ~t[332]);
  assign t[284] = (t[333] & ~t[334]);
  assign t[285] = (t[335] & ~t[336]);
  assign t[286] = (t[337] & ~t[338]);
  assign t[287] = (t[339] & ~t[340]);
  assign t[288] = (t[341] & ~t[342]);
  assign t[289] = t[343] ^ x[4];
  assign t[28] = t[41] ^ t[42];
  assign t[290] = t[344] ^ x[3];
  assign t[291] = t[345] ^ x[7];
  assign t[292] = t[346] ^ x[6];
  assign t[293] = t[347] ^ x[10];
  assign t[294] = t[348] ^ x[9];
  assign t[295] = t[349] ^ x[13];
  assign t[296] = t[350] ^ x[12];
  assign t[297] = t[351] ^ x[18];
  assign t[298] = t[352] ^ x[17];
  assign t[299] = t[353] ^ x[21];
  assign t[29] = t[43] ^ t[44];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[20];
  assign t[301] = t[355] ^ x[24];
  assign t[302] = t[356] ^ x[23];
  assign t[303] = t[357] ^ x[27];
  assign t[304] = t[358] ^ x[26];
  assign t[305] = t[359] ^ x[30];
  assign t[306] = t[360] ^ x[29];
  assign t[307] = t[361] ^ x[33];
  assign t[308] = t[362] ^ x[32];
  assign t[309] = t[363] ^ x[36];
  assign t[30] = t[45] & t[46];
  assign t[310] = t[364] ^ x[35];
  assign t[311] = t[365] ^ x[39];
  assign t[312] = t[366] ^ x[38];
  assign t[313] = t[367] ^ x[42];
  assign t[314] = t[368] ^ x[41];
  assign t[315] = t[369] ^ x[45];
  assign t[316] = t[370] ^ x[44];
  assign t[317] = t[371] ^ x[52];
  assign t[318] = t[372] ^ x[51];
  assign t[319] = t[373] ^ x[55];
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = t[374] ^ x[54];
  assign t[321] = t[375] ^ x[58];
  assign t[322] = t[376] ^ x[57];
  assign t[323] = t[377] ^ x[61];
  assign t[324] = t[378] ^ x[60];
  assign t[325] = t[379] ^ x[64];
  assign t[326] = t[380] ^ x[63];
  assign t[327] = t[381] ^ x[67];
  assign t[328] = t[382] ^ x[66];
  assign t[329] = t[383] ^ x[70];
  assign t[32] = ~(t[49]);
  assign t[330] = t[384] ^ x[69];
  assign t[331] = t[385] ^ x[77];
  assign t[332] = t[386] ^ x[76];
  assign t[333] = t[387] ^ x[80];
  assign t[334] = t[388] ^ x[79];
  assign t[335] = t[389] ^ x[83];
  assign t[336] = t[390] ^ x[82];
  assign t[337] = t[391] ^ x[86];
  assign t[338] = t[392] ^ x[85];
  assign t[339] = t[393] ^ x[91];
  assign t[33] = ~(t[214]);
  assign t[340] = t[394] ^ x[90];
  assign t[341] = t[395] ^ x[94];
  assign t[342] = t[396] ^ x[93];
  assign t[343] = (x[2]);
  assign t[344] = (x[2]);
  assign t[345] = (x[5]);
  assign t[346] = (x[5]);
  assign t[347] = (x[8]);
  assign t[348] = (x[8]);
  assign t[349] = (x[11]);
  assign t[34] = ~(t[50] ^ t[51]);
  assign t[350] = (x[11]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[52] ^ t[53]);
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = t[17] ^ t[54];
  assign t[370] = (x[43]);
  assign t[371] = (x[50]);
  assign t[372] = (x[50]);
  assign t[373] = (x[53]);
  assign t[374] = (x[53]);
  assign t[375] = (x[56]);
  assign t[376] = (x[56]);
  assign t[377] = (x[59]);
  assign t[378] = (x[59]);
  assign t[379] = (x[62]);
  assign t[37] = ~(t[55] ^ t[56]);
  assign t[380] = (x[62]);
  assign t[381] = (x[65]);
  assign t[382] = (x[65]);
  assign t[383] = (x[68]);
  assign t[384] = (x[68]);
  assign t[385] = (x[75]);
  assign t[386] = (x[75]);
  assign t[387] = (x[78]);
  assign t[388] = (x[78]);
  assign t[389] = (x[81]);
  assign t[38] = t[57] ^ t[58];
  assign t[390] = (x[81]);
  assign t[391] = (x[84]);
  assign t[392] = (x[84]);
  assign t[393] = (x[89]);
  assign t[394] = (x[89]);
  assign t[395] = (x[92]);
  assign t[396] = (x[92]);
  assign t[39] = t[59] ^ t[52];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = t[44] ^ t[62];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[9] ? t[65] : t[215];
  assign t[44] = t[9] ? t[66] : t[216];
  assign t[45] = ~(t[29] ^ t[63]);
  assign t[46] = t[41] ^ t[67];
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = t[217] | t[70];
  assign t[49] = ~(t[71]);
  assign t[4] = t[9] ? t[10] : t[208];
  assign t[50] = ~(t[72] ^ t[73]);
  assign t[51] = t[74] ^ t[75];
  assign t[52] = t[76] ^ t[77];
  assign t[53] = t[78] ^ t[79];
  assign t[54] = ~(t[80] ^ t[81]);
  assign t[55] = t[82] ^ t[34];
  assign t[56] = ~(t[83] ^ t[84]);
  assign t[57] = t[85] ^ t[76];
  assign t[58] = t[86] & t[87];
  assign t[59] = t[88] ^ t[89];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92] & t[93];
  assign t[62] = t[9] ? t[94] : t[218];
  assign t[63] = t[95] ^ t[96];
  assign t[64] = t[97] & t[98];
  assign t[65] = t[215] ^ t[99];
  assign t[66] = t[216] ^ t[100];
  assign t[67] = t[9] ? t[101] : t[219];
  assign t[68] = ~(t[70] & t[102]);
  assign t[69] = ~(t[220] ^ t[103]);
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = ~(t[104] & t[105]);
  assign t[71] = ~(t[48]);
  assign t[72] = t[106] ^ t[107];
  assign t[73] = t[108] ^ t[109];
  assign t[74] = t[91] ^ t[108];
  assign t[75] = t[110] ^ t[111];
  assign t[76] = t[212] ^ t[112];
  assign t[77] = t[113] ^ t[107];
  assign t[78] = t[114] ^ t[115];
  assign t[79] = t[116] ^ t[117];
  assign t[7] = t[15] ^ t[16];
  assign t[80] = t[51] ^ t[38];
  assign t[81] = ~(t[118] ^ t[84]);
  assign t[82] = t[118] ^ t[119];
  assign t[83] = t[120] ^ t[121];
  assign t[84] = t[122] ^ t[123];
  assign t[85] = t[31] ? t[124] : t[221];
  assign t[86] = ~(t[125]);
  assign t[87] = t[214] ^ t[126];
  assign t[88] = t[127] ^ t[122];
  assign t[89] = t[128] ^ t[129];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = ~t[130];
  assign t[91] = t[131];
  assign t[92] = ~(t[60] ^ t[110]);
  assign t[93] = t[74] ^ t[132];
  assign t[94] = t[218] ^ t[133];
  assign t[95] = t[134] & t[135];
  assign t[96] = t[136] & t[67];
  assign t[97] = ~(t[95] ^ t[137]);
  assign t[98] = t[138] ^ t[139];
  assign t[99] = t[140] ? x[47] : x[46];
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [116:0] x;
 output y;

 wire [396:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ? x[49] : x[48];
  assign t[101] = t[219] ^ t[141];
  assign t[102] = ~(t[142] & t[143]);
  assign t[103] = t[144] ^ t[222];
  assign t[104] = ~(t[220]);
  assign t[105] = t[145] & t[144];
  assign t[106] = t[85] ^ t[125];
  assign t[107] = t[146] & t[147];
  assign t[108] = t[148];
  assign t[109] = t[110] ^ t[61];
  assign t[10] = t[208] ^ t[20];
  assign t[110] = t[149] ^ t[150];
  assign t[111] = t[151] & t[152];
  assign t[112] = t[153] ? t[154] : t[223];
  assign t[113] = t[155] ^ t[58];
  assign t[114] = t[125] ^ t[76];
  assign t[115] = t[113] ^ t[156];
  assign t[116] = t[157] ^ t[127];
  assign t[117] = t[158] & t[159];
  assign t[118] = t[62] ^ t[160];
  assign t[119] = t[138] ^ t[96];
  assign t[11] = ~(t[209]);
  assign t[120] = t[157] ^ t[122];
  assign t[121] = t[161] & t[162];
  assign t[122] = t[9] ? t[163] : t[224];
  assign t[123] = t[128] ^ t[117];
  assign t[124] = t[221] ^ t[164];
  assign t[125] = t[211] ^ t[165];
  assign t[126] = t[31] ? t[166] : t[225];
  assign t[127] = t[9] ? t[167] : t[226];
  assign t[128] = t[168] ^ t[121];
  assign t[129] = t[169] & t[170];
  assign t[12] = ~(t[210]);
  assign t[130] = t[31] ? t[171] : t[227];
  assign t[131] = t[31] ? t[172] : t[228];
  assign t[132] = t[173];
  assign t[133] = t[140] ? x[72] : x[71];
  assign t[134] = ~(t[139]);
  assign t[135] = ~(t[43]);
  assign t[136] = ~(t[44]);
  assign t[137] = t[41] ^ t[43];
  assign t[138] = t[43] ^ t[62];
  assign t[139] = t[67] ^ t[44];
  assign t[13] = ~(t[211]);
  assign t[140] = ~(t[49]);
  assign t[141] = t[140] ? x[74] : x[73];
  assign t[142] = ~(t[145] | t[144]);
  assign t[143] = ~(t[174] | t[104]);
  assign t[144] = ~(t[229]);
  assign t[145] = ~(t[222]);
  assign t[146] = ~(t[106] ^ t[113]);
  assign t[147] = t[114] ^ t[87];
  assign t[148] = t[31] ? t[175] : t[230];
  assign t[149] = t[176] & t[177];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = t[178] & t[132];
  assign t[151] = ~(t[149] ^ t[179]);
  assign t[152] = t[180] ^ t[181];
  assign t[153] = ~(t[19]);
  assign t[154] = t[223] ^ t[182];
  assign t[155] = t[183] & t[184];
  assign t[156] = t[185] & t[186];
  assign t[157] = t[9] ? t[187] : t[231];
  assign t[158] = ~(t[116] ^ t[128]);
  assign t[159] = t[88] ^ t[162];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[63] ^ t[30];
  assign t[161] = ~(t[127]);
  assign t[162] = t[9] ? t[188] : t[232];
  assign t[163] = t[224] ^ t[189];
  assign t[164] = t[140] ? x[88] : x[87];
  assign t[165] = t[31] ? t[190] : t[233];
  assign t[166] = t[225] ^ t[191];
  assign t[167] = t[226] ^ t[192];
  assign t[168] = t[193] & t[194];
  assign t[169] = ~(t[168] ^ t[195]);
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = t[120] ^ t[196];
  assign t[171] = t[227] ^ t[197];
  assign t[172] = t[228] ^ t[198];
  assign t[173] = t[31] ? t[199] : t[234];
  assign t[174] = ~(t[217]);
  assign t[175] = t[230] ^ t[200];
  assign t[176] = ~(t[181]);
  assign t[177] = ~(t[90]);
  assign t[178] = ~(t[91]);
  assign t[179] = t[74] ^ t[90];
  assign t[17] = ~(t[27] ^ t[28]);
  assign t[180] = t[90] ^ t[108];
  assign t[181] = t[132] ^ t[91];
  assign t[182] = t[201] ? x[96] : x[95];
  assign t[183] = ~(t[202]);
  assign t[184] = ~(t[85]);
  assign t[185] = ~(t[155] ^ t[203]);
  assign t[186] = t[57] ^ t[202];
  assign t[187] = t[231] ^ t[204];
  assign t[188] = t[232] ^ t[205];
  assign t[189] = t[32] ? x[98] : x[97];
  assign t[18] = t[29] ^ t[30];
  assign t[190] = t[233] ^ t[206];
  assign t[191] = t[71] ? x[100] : x[99];
  assign t[192] = t[32] ? x[102] : x[101];
  assign t[193] = ~(t[196]);
  assign t[194] = ~(t[157]);
  assign t[195] = t[88] ^ t[157];
  assign t[196] = t[162] ^ t[127];
  assign t[197] = t[71] ? x[104] : x[103];
  assign t[198] = t[201] ? x[106] : x[105];
  assign t[199] = t[234] ^ t[207];
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[71] ? x[108] : x[107];
  assign t[201] = ~(t[49]);
  assign t[202] = t[87] ^ t[125];
  assign t[203] = t[114] ^ t[85];
  assign t[204] = t[32] ? x[110] : x[109];
  assign t[205] = t[32] ? x[112] : x[111];
  assign t[206] = t[140] ? x[114] : x[113];
  assign t[207] = t[201] ? x[116] : x[115];
  assign t[208] = (t[235]);
  assign t[209] = (t[236]);
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[212]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[33] & t[213]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = t[262] ^ x[4];
  assign t[236] = t[263] ^ x[7];
  assign t[237] = t[264] ^ x[10];
  assign t[238] = t[265] ^ x[13];
  assign t[239] = t[266] ^ x[18];
  assign t[23] = ~(t[28] ^ t[34]);
  assign t[240] = t[267] ^ x[21];
  assign t[241] = t[268] ^ x[24];
  assign t[242] = t[269] ^ x[27];
  assign t[243] = t[270] ^ x[30];
  assign t[244] = t[271] ^ x[33];
  assign t[245] = t[272] ^ x[36];
  assign t[246] = t[273] ^ x[39];
  assign t[247] = t[274] ^ x[42];
  assign t[248] = t[275] ^ x[45];
  assign t[249] = t[276] ^ x[52];
  assign t[24] = ~(t[35] ^ t[36]);
  assign t[250] = t[277] ^ x[55];
  assign t[251] = t[278] ^ x[58];
  assign t[252] = t[279] ^ x[61];
  assign t[253] = t[280] ^ x[64];
  assign t[254] = t[281] ^ x[67];
  assign t[255] = t[282] ^ x[70];
  assign t[256] = t[283] ^ x[77];
  assign t[257] = t[284] ^ x[80];
  assign t[258] = t[285] ^ x[83];
  assign t[259] = t[286] ^ x[86];
  assign t[25] = t[37] ^ t[38];
  assign t[260] = t[287] ^ x[91];
  assign t[261] = t[288] ^ x[94];
  assign t[262] = (t[289] & ~t[290]);
  assign t[263] = (t[291] & ~t[292]);
  assign t[264] = (t[293] & ~t[294]);
  assign t[265] = (t[295] & ~t[296]);
  assign t[266] = (t[297] & ~t[298]);
  assign t[267] = (t[299] & ~t[300]);
  assign t[268] = (t[301] & ~t[302]);
  assign t[269] = (t[303] & ~t[304]);
  assign t[26] = ~(t[39] ^ t[18]);
  assign t[270] = (t[305] & ~t[306]);
  assign t[271] = (t[307] & ~t[308]);
  assign t[272] = (t[309] & ~t[310]);
  assign t[273] = (t[311] & ~t[312]);
  assign t[274] = (t[313] & ~t[314]);
  assign t[275] = (t[315] & ~t[316]);
  assign t[276] = (t[317] & ~t[318]);
  assign t[277] = (t[319] & ~t[320]);
  assign t[278] = (t[321] & ~t[322]);
  assign t[279] = (t[323] & ~t[324]);
  assign t[27] = ~(t[39] ^ t[40]);
  assign t[280] = (t[325] & ~t[326]);
  assign t[281] = (t[327] & ~t[328]);
  assign t[282] = (t[329] & ~t[330]);
  assign t[283] = (t[331] & ~t[332]);
  assign t[284] = (t[333] & ~t[334]);
  assign t[285] = (t[335] & ~t[336]);
  assign t[286] = (t[337] & ~t[338]);
  assign t[287] = (t[339] & ~t[340]);
  assign t[288] = (t[341] & ~t[342]);
  assign t[289] = t[343] ^ x[4];
  assign t[28] = t[41] ^ t[42];
  assign t[290] = t[344] ^ x[3];
  assign t[291] = t[345] ^ x[7];
  assign t[292] = t[346] ^ x[6];
  assign t[293] = t[347] ^ x[10];
  assign t[294] = t[348] ^ x[9];
  assign t[295] = t[349] ^ x[13];
  assign t[296] = t[350] ^ x[12];
  assign t[297] = t[351] ^ x[18];
  assign t[298] = t[352] ^ x[17];
  assign t[299] = t[353] ^ x[21];
  assign t[29] = t[43] ^ t[44];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[20];
  assign t[301] = t[355] ^ x[24];
  assign t[302] = t[356] ^ x[23];
  assign t[303] = t[357] ^ x[27];
  assign t[304] = t[358] ^ x[26];
  assign t[305] = t[359] ^ x[30];
  assign t[306] = t[360] ^ x[29];
  assign t[307] = t[361] ^ x[33];
  assign t[308] = t[362] ^ x[32];
  assign t[309] = t[363] ^ x[36];
  assign t[30] = t[45] & t[46];
  assign t[310] = t[364] ^ x[35];
  assign t[311] = t[365] ^ x[39];
  assign t[312] = t[366] ^ x[38];
  assign t[313] = t[367] ^ x[42];
  assign t[314] = t[368] ^ x[41];
  assign t[315] = t[369] ^ x[45];
  assign t[316] = t[370] ^ x[44];
  assign t[317] = t[371] ^ x[52];
  assign t[318] = t[372] ^ x[51];
  assign t[319] = t[373] ^ x[55];
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = t[374] ^ x[54];
  assign t[321] = t[375] ^ x[58];
  assign t[322] = t[376] ^ x[57];
  assign t[323] = t[377] ^ x[61];
  assign t[324] = t[378] ^ x[60];
  assign t[325] = t[379] ^ x[64];
  assign t[326] = t[380] ^ x[63];
  assign t[327] = t[381] ^ x[67];
  assign t[328] = t[382] ^ x[66];
  assign t[329] = t[383] ^ x[70];
  assign t[32] = ~(t[49]);
  assign t[330] = t[384] ^ x[69];
  assign t[331] = t[385] ^ x[77];
  assign t[332] = t[386] ^ x[76];
  assign t[333] = t[387] ^ x[80];
  assign t[334] = t[388] ^ x[79];
  assign t[335] = t[389] ^ x[83];
  assign t[336] = t[390] ^ x[82];
  assign t[337] = t[391] ^ x[86];
  assign t[338] = t[392] ^ x[85];
  assign t[339] = t[393] ^ x[91];
  assign t[33] = ~(t[214]);
  assign t[340] = t[394] ^ x[90];
  assign t[341] = t[395] ^ x[94];
  assign t[342] = t[396] ^ x[93];
  assign t[343] = (x[2]);
  assign t[344] = (x[2]);
  assign t[345] = (x[5]);
  assign t[346] = (x[5]);
  assign t[347] = (x[8]);
  assign t[348] = (x[8]);
  assign t[349] = (x[11]);
  assign t[34] = ~(t[50] ^ t[51]);
  assign t[350] = (x[11]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[52] ^ t[53]);
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = t[17] ^ t[54];
  assign t[370] = (x[43]);
  assign t[371] = (x[50]);
  assign t[372] = (x[50]);
  assign t[373] = (x[53]);
  assign t[374] = (x[53]);
  assign t[375] = (x[56]);
  assign t[376] = (x[56]);
  assign t[377] = (x[59]);
  assign t[378] = (x[59]);
  assign t[379] = (x[62]);
  assign t[37] = ~(t[55] ^ t[56]);
  assign t[380] = (x[62]);
  assign t[381] = (x[65]);
  assign t[382] = (x[65]);
  assign t[383] = (x[68]);
  assign t[384] = (x[68]);
  assign t[385] = (x[75]);
  assign t[386] = (x[75]);
  assign t[387] = (x[78]);
  assign t[388] = (x[78]);
  assign t[389] = (x[81]);
  assign t[38] = t[57] ^ t[58];
  assign t[390] = (x[81]);
  assign t[391] = (x[84]);
  assign t[392] = (x[84]);
  assign t[393] = (x[89]);
  assign t[394] = (x[89]);
  assign t[395] = (x[92]);
  assign t[396] = (x[92]);
  assign t[39] = t[59] ^ t[52];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = t[44] ^ t[62];
  assign t[42] = t[63] ^ t[64];
  assign t[43] = t[9] ? t[65] : t[215];
  assign t[44] = t[9] ? t[66] : t[216];
  assign t[45] = ~(t[29] ^ t[63]);
  assign t[46] = t[41] ^ t[67];
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = t[217] | t[70];
  assign t[49] = ~(t[71]);
  assign t[4] = t[9] ? t[10] : t[208];
  assign t[50] = ~(t[72] ^ t[73]);
  assign t[51] = t[74] ^ t[75];
  assign t[52] = t[76] ^ t[77];
  assign t[53] = t[78] ^ t[79];
  assign t[54] = ~(t[80] ^ t[81]);
  assign t[55] = t[82] ^ t[34];
  assign t[56] = ~(t[83] ^ t[84]);
  assign t[57] = t[85] ^ t[76];
  assign t[58] = t[86] & t[87];
  assign t[59] = t[88] ^ t[89];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92] & t[93];
  assign t[62] = t[9] ? t[94] : t[218];
  assign t[63] = t[95] ^ t[96];
  assign t[64] = t[97] & t[98];
  assign t[65] = t[215] ^ t[99];
  assign t[66] = t[216] ^ t[100];
  assign t[67] = t[9] ? t[101] : t[219];
  assign t[68] = ~(t[70] & t[102]);
  assign t[69] = ~(t[220] ^ t[103]);
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = ~(t[104] & t[105]);
  assign t[71] = ~(t[48]);
  assign t[72] = t[106] ^ t[107];
  assign t[73] = t[108] ^ t[109];
  assign t[74] = t[91] ^ t[108];
  assign t[75] = t[110] ^ t[111];
  assign t[76] = t[212] ^ t[112];
  assign t[77] = t[113] ^ t[107];
  assign t[78] = t[114] ^ t[115];
  assign t[79] = t[116] ^ t[117];
  assign t[7] = t[15] ^ t[16];
  assign t[80] = t[51] ^ t[38];
  assign t[81] = ~(t[118] ^ t[84]);
  assign t[82] = t[118] ^ t[119];
  assign t[83] = t[120] ^ t[121];
  assign t[84] = t[122] ^ t[123];
  assign t[85] = t[31] ? t[124] : t[221];
  assign t[86] = ~(t[125]);
  assign t[87] = t[214] ^ t[126];
  assign t[88] = t[127] ^ t[122];
  assign t[89] = t[128] ^ t[129];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = ~t[130];
  assign t[91] = t[131];
  assign t[92] = ~(t[60] ^ t[110]);
  assign t[93] = t[74] ^ t[132];
  assign t[94] = t[218] ^ t[133];
  assign t[95] = t[134] & t[135];
  assign t[96] = t[136] & t[67];
  assign t[97] = ~(t[95] ^ t[137]);
  assign t[98] = t[138] ^ t[139];
  assign t[99] = t[140] ? x[47] : x[46];
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[221] ^ t[143];
  assign t[101] = t[222] ^ t[144];
  assign t[102] = ~(t[114] ^ t[56]);
  assign t[103] = t[36] ^ t[124];
  assign t[104] = t[145] ? x[59] : x[58];
  assign t[105] = t[146] & t[147];
  assign t[106] = t[148] & t[149];
  assign t[107] = ~(t[91] ^ t[71]);
  assign t[108] = t[150] ^ t[149];
  assign t[109] = ~(t[151] & t[152]);
  assign t[10] = t[210] ^ t[20];
  assign t[110] = t[153] ^ t[228];
  assign t[111] = ~(t[223]);
  assign t[112] = t[154] & t[153];
  assign t[113] = t[155] ^ t[61];
  assign t[114] = t[156] ^ t[55];
  assign t[115] = t[119] ^ t[157];
  assign t[116] = t[62] ^ t[158];
  assign t[117] = t[224] ^ t[159];
  assign t[118] = t[160] ^ t[43];
  assign t[119] = t[81] ^ t[65];
  assign t[11] = ~(t[211]);
  assign t[120] = t[225] ^ t[161];
  assign t[121] = ~(t[127]);
  assign t[122] = ~(t[156]);
  assign t[123] = ~(t[55]);
  assign t[124] = t[162];
  assign t[125] = t[36] ^ t[156];
  assign t[126] = t[156] ^ t[44];
  assign t[127] = t[124] ^ t[55];
  assign t[128] = ~(t[163] ^ t[164]);
  assign t[129] = t[165] ^ t[166];
  assign t[12] = ~(t[212]);
  assign t[130] = t[9] ? t[167] : t[229];
  assign t[131] = t[9] ? t[168] : t[230];
  assign t[132] = ~(t[19]);
  assign t[133] = t[226] ^ t[169];
  assign t[134] = t[227] ^ t[170];
  assign t[135] = ~(t[140]);
  assign t[136] = ~(t[155]);
  assign t[137] = ~(t[60]);
  assign t[138] = t[212] ^ t[171];
  assign t[139] = t[40] ^ t[155];
  assign t[13] = ~(t[213]);
  assign t[140] = t[138] ^ t[60];
  assign t[141] = t[32] ? x[70] : x[69];
  assign t[142] = t[76] ? x[72] : x[71];
  assign t[143] = t[76] ? x[74] : x[73];
  assign t[144] = t[145] ? x[76] : x[75];
  assign t[145] = ~(t[50]);
  assign t[146] = ~(t[172]);
  assign t[147] = ~(t[130]);
  assign t[148] = ~(t[131]);
  assign t[149] = t[9] ? t[173] : t[231];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = t[131] ^ t[46];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[174] | t[111]);
  assign t[153] = ~(t[232]);
  assign t[154] = ~(t[228]);
  assign t[155] = t[132] ? t[175] : t[233];
  assign t[156] = t[176];
  assign t[157] = t[118] ^ t[177];
  assign t[158] = t[178] & t[179];
  assign t[159] = t[32] ? x[87] : x[86];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[180] & t[181];
  assign t[161] = t[145] ? x[89] : x[88];
  assign t[162] = t[31] ? t[182] : t[234];
  assign t[163] = t[183] ^ t[184];
  assign t[164] = ~(t[185] ^ t[30]);
  assign t[165] = t[150] ^ t[186];
  assign t[166] = t[65] ^ t[187];
  assign t[167] = t[229] ^ t[188];
  assign t[168] = t[230] ^ t[189];
  assign t[169] = t[190] ? x[94] : x[93];
  assign t[16] = t[25] ^ t[26];
  assign t[170] = t[190] ? x[96] : x[95];
  assign t[171] = t[132] ? t[191] : t[235];
  assign t[172] = t[149] ^ t[131];
  assign t[173] = t[231] ^ t[192];
  assign t[174] = ~(t[218]);
  assign t[175] = t[233] ^ t[193];
  assign t[176] = t[9] ? t[194] : t[236];
  assign t[177] = t[195] & t[196];
  assign t[178] = ~(t[197] ^ t[62]);
  assign t[179] = t[40] ^ t[138];
  assign t[17] = t[27] ^ t[28];
  assign t[180] = ~(t[198]);
  assign t[181] = ~(t[64]);
  assign t[182] = t[234] ^ t[199];
  assign t[183] = t[29] ^ t[200];
  assign t[184] = ~(t[201] ^ t[27]);
  assign t[185] = t[202] ^ t[106];
  assign t[186] = t[71] ^ t[203];
  assign t[187] = t[118] ^ t[54];
  assign t[188] = t[145] ? x[104] : x[103];
  assign t[189] = t[145] ? x[106] : x[105];
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[190] = ~(t[50]);
  assign t[191] = t[235] ^ t[204];
  assign t[192] = t[145] ? x[108] : x[107];
  assign t[193] = t[190] ? x[110] : x[109];
  assign t[194] = t[236] ^ t[205];
  assign t[195] = ~(t[160] ^ t[206]);
  assign t[196] = t[42] ^ t[198];
  assign t[197] = t[155] ^ t[60];
  assign t[198] = t[67] ^ t[81];
  assign t[199] = t[145] ? x[112] : x[111];
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[126] ^ t[86];
  assign t[201] = ~(t[35] ^ t[80]);
  assign t[202] = t[130] ^ t[46];
  assign t[203] = t[207] & t[208];
  assign t[204] = t[190] ? x[114] : x[113];
  assign t[205] = t[145] ? x[116] : x[115];
  assign t[206] = t[119] ^ t[64];
  assign t[207] = ~(t[105] ^ t[209]);
  assign t[208] = t[202] ^ t[172];
  assign t[209] = t[150] ^ t[130];
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[214]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[33] & t[215]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[7];
  assign t[239] = t[266] ^ x[10];
  assign t[23] = t[34] ^ t[35];
  assign t[240] = t[267] ^ x[13];
  assign t[241] = t[268] ^ x[18];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = ~(t[25] ^ t[30]);
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[51];
  assign t[253] = t[280] ^ x[54];
  assign t[254] = t[281] ^ x[57];
  assign t[255] = t[282] ^ x[62];
  assign t[256] = t[283] ^ x[65];
  assign t[257] = t[284] ^ x[68];
  assign t[258] = t[285] ^ x[79];
  assign t[259] = t[286] ^ x[82];
  assign t[25] = t[36] ^ t[37];
  assign t[260] = t[287] ^ x[85];
  assign t[261] = t[288] ^ x[92];
  assign t[262] = t[289] ^ x[99];
  assign t[263] = t[290] ^ x[102];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = t[42] ^ t[43];
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[7];
  assign t[294] = t[348] ^ x[6];
  assign t[295] = t[349] ^ x[10];
  assign t[296] = t[350] ^ x[9];
  assign t[297] = t[351] ^ x[13];
  assign t[298] = t[352] ^ x[12];
  assign t[299] = t[353] ^ x[18];
  assign t[29] = t[44] ^ t[45];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[17];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = t[46] ^ t[47];
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[51];
  assign t[322] = t[376] ^ x[50];
  assign t[323] = t[377] ^ x[54];
  assign t[324] = t[378] ^ x[53];
  assign t[325] = t[379] ^ x[57];
  assign t[326] = t[380] ^ x[56];
  assign t[327] = t[381] ^ x[62];
  assign t[328] = t[382] ^ x[61];
  assign t[329] = t[383] ^ x[65];
  assign t[32] = ~(t[50]);
  assign t[330] = t[384] ^ x[64];
  assign t[331] = t[385] ^ x[68];
  assign t[332] = t[386] ^ x[67];
  assign t[333] = t[387] ^ x[79];
  assign t[334] = t[388] ^ x[78];
  assign t[335] = t[389] ^ x[82];
  assign t[336] = t[390] ^ x[81];
  assign t[337] = t[391] ^ x[85];
  assign t[338] = t[392] ^ x[84];
  assign t[339] = t[393] ^ x[92];
  assign t[33] = ~(t[216]);
  assign t[340] = t[394] ^ x[91];
  assign t[341] = t[395] ^ x[99];
  assign t[342] = t[396] ^ x[98];
  assign t[343] = t[397] ^ x[102];
  assign t[344] = t[398] ^ x[101];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[5]);
  assign t[348] = (x[5]);
  assign t[349] = (x[8]);
  assign t[34] = ~(t[51] ^ t[52]);
  assign t[350] = (x[8]);
  assign t[351] = (x[11]);
  assign t[352] = (x[11]);
  assign t[353] = (x[16]);
  assign t[354] = (x[16]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = t[53] ^ t[54];
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = t[55] ^ t[44];
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[49]);
  assign t[376] = (x[49]);
  assign t[377] = (x[52]);
  assign t[378] = (x[52]);
  assign t[379] = (x[55]);
  assign t[37] = t[56] ^ t[57];
  assign t[380] = (x[55]);
  assign t[381] = (x[60]);
  assign t[382] = (x[60]);
  assign t[383] = (x[63]);
  assign t[384] = (x[63]);
  assign t[385] = (x[66]);
  assign t[386] = (x[66]);
  assign t[387] = (x[77]);
  assign t[388] = (x[77]);
  assign t[389] = (x[80]);
  assign t[38] = t[58] ^ t[34];
  assign t[390] = (x[80]);
  assign t[391] = (x[83]);
  assign t[392] = (x[83]);
  assign t[393] = (x[90]);
  assign t[394] = (x[90]);
  assign t[395] = (x[97]);
  assign t[396] = (x[97]);
  assign t[397] = (x[100]);
  assign t[398] = (x[100]);
  assign t[39] = ~(t[29] ^ t[59]);
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = ~t[68];
  assign t[45] = t[56] ^ t[69];
  assign t[46] = t[9] ? t[70] : t[217];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[218] | t[75];
  assign t[4] = t[9] ? t[10] : t[210];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[64] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = ~t[84];
  assign t[56] = t[85] ^ t[86];
  assign t[57] = t[87] & t[88];
  assign t[58] = ~(t[89] ^ t[90]);
  assign t[59] = t[91] ^ t[72];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[211] ^ t[92];
  assign t[61] = t[215] ^ t[93];
  assign t[62] = t[94] ^ t[95];
  assign t[63] = t[96] & t[97];
  assign t[64] = t[31] ? t[98] : t[219];
  assign t[65] = t[31] ? t[99] : t[220];
  assign t[66] = ~(t[81]);
  assign t[67] = t[31] ? t[100] : t[221];
  assign t[68] = t[9] ? t[101] : t[222];
  assign t[69] = t[102] & t[103];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[217] ^ t[104];
  assign t[71] = t[105] ^ t[106];
  assign t[72] = t[107] & t[108];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[223] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[113] ^ t[95];
  assign t[78] = t[114] ^ t[69];
  assign t[79] = t[115] ^ t[59];
  assign t[7] = ~(t[15] ^ t[16]);
  assign t[80] = t[61] ^ t[116];
  assign t[81] = t[31] ? t[117] : t[224];
  assign t[82] = ~(t[53] ^ t[118]);
  assign t[83] = t[119] ^ t[67];
  assign t[84] = t[9] ? t[120] : t[225];
  assign t[85] = t[121] & t[122];
  assign t[86] = t[123] & t[124];
  assign t[87] = ~(t[85] ^ t[125]);
  assign t[88] = t[126] ^ t[127];
  assign t[89] = t[128] ^ t[28];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = ~(t[129] ^ t[78]);
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[132] ? t[133] : t[226];
  assign t[93] = t[132] ? t[134] : t[227];
  assign t[94] = t[135] & t[136];
  assign t[95] = t[137] & t[138];
  assign t[96] = ~(t[94] ^ t[139]);
  assign t[97] = t[113] ^ t[140];
  assign t[98] = t[219] ^ t[141];
  assign t[99] = t[220] ^ t[142];
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[221] ^ t[143];
  assign t[101] = t[222] ^ t[144];
  assign t[102] = ~(t[114] ^ t[56]);
  assign t[103] = t[36] ^ t[124];
  assign t[104] = t[145] ? x[59] : x[58];
  assign t[105] = t[146] & t[147];
  assign t[106] = t[148] & t[149];
  assign t[107] = ~(t[91] ^ t[71]);
  assign t[108] = t[150] ^ t[149];
  assign t[109] = ~(t[151] & t[152]);
  assign t[10] = t[210] ^ t[20];
  assign t[110] = t[153] ^ t[228];
  assign t[111] = ~(t[223]);
  assign t[112] = t[154] & t[153];
  assign t[113] = t[155] ^ t[61];
  assign t[114] = t[156] ^ t[55];
  assign t[115] = t[119] ^ t[157];
  assign t[116] = t[62] ^ t[158];
  assign t[117] = t[224] ^ t[159];
  assign t[118] = t[160] ^ t[43];
  assign t[119] = t[81] ^ t[65];
  assign t[11] = ~(t[211]);
  assign t[120] = t[225] ^ t[161];
  assign t[121] = ~(t[127]);
  assign t[122] = ~(t[156]);
  assign t[123] = ~(t[55]);
  assign t[124] = t[162];
  assign t[125] = t[36] ^ t[156];
  assign t[126] = t[156] ^ t[44];
  assign t[127] = t[124] ^ t[55];
  assign t[128] = ~(t[163] ^ t[164]);
  assign t[129] = t[165] ^ t[166];
  assign t[12] = ~(t[212]);
  assign t[130] = t[9] ? t[167] : t[229];
  assign t[131] = t[9] ? t[168] : t[230];
  assign t[132] = ~(t[19]);
  assign t[133] = t[226] ^ t[169];
  assign t[134] = t[227] ^ t[170];
  assign t[135] = ~(t[140]);
  assign t[136] = ~(t[155]);
  assign t[137] = ~(t[60]);
  assign t[138] = t[212] ^ t[171];
  assign t[139] = t[40] ^ t[155];
  assign t[13] = ~(t[213]);
  assign t[140] = t[138] ^ t[60];
  assign t[141] = t[32] ? x[70] : x[69];
  assign t[142] = t[76] ? x[72] : x[71];
  assign t[143] = t[76] ? x[74] : x[73];
  assign t[144] = t[145] ? x[76] : x[75];
  assign t[145] = ~(t[50]);
  assign t[146] = ~(t[172]);
  assign t[147] = ~(t[130]);
  assign t[148] = ~(t[131]);
  assign t[149] = t[9] ? t[173] : t[231];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = t[131] ^ t[46];
  assign t[151] = ~(t[154] | t[153]);
  assign t[152] = ~(t[174] | t[111]);
  assign t[153] = ~(t[232]);
  assign t[154] = ~(t[228]);
  assign t[155] = t[132] ? t[175] : t[233];
  assign t[156] = t[176];
  assign t[157] = t[118] ^ t[177];
  assign t[158] = t[178] & t[179];
  assign t[159] = t[32] ? x[87] : x[86];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[180] & t[181];
  assign t[161] = t[145] ? x[89] : x[88];
  assign t[162] = t[31] ? t[182] : t[234];
  assign t[163] = t[183] ^ t[184];
  assign t[164] = ~(t[185] ^ t[30]);
  assign t[165] = t[150] ^ t[186];
  assign t[166] = t[65] ^ t[187];
  assign t[167] = t[229] ^ t[188];
  assign t[168] = t[230] ^ t[189];
  assign t[169] = t[190] ? x[94] : x[93];
  assign t[16] = t[25] ^ t[26];
  assign t[170] = t[190] ? x[96] : x[95];
  assign t[171] = t[132] ? t[191] : t[235];
  assign t[172] = t[149] ^ t[131];
  assign t[173] = t[231] ^ t[192];
  assign t[174] = ~(t[218]);
  assign t[175] = t[233] ^ t[193];
  assign t[176] = t[9] ? t[194] : t[236];
  assign t[177] = t[195] & t[196];
  assign t[178] = ~(t[197] ^ t[62]);
  assign t[179] = t[40] ^ t[138];
  assign t[17] = t[27] ^ t[28];
  assign t[180] = ~(t[198]);
  assign t[181] = ~(t[64]);
  assign t[182] = t[234] ^ t[199];
  assign t[183] = t[29] ^ t[200];
  assign t[184] = ~(t[201] ^ t[27]);
  assign t[185] = t[202] ^ t[106];
  assign t[186] = t[71] ^ t[203];
  assign t[187] = t[118] ^ t[54];
  assign t[188] = t[145] ? x[104] : x[103];
  assign t[189] = t[145] ? x[106] : x[105];
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[190] = ~(t[50]);
  assign t[191] = t[235] ^ t[204];
  assign t[192] = t[145] ? x[108] : x[107];
  assign t[193] = t[190] ? x[110] : x[109];
  assign t[194] = t[236] ^ t[205];
  assign t[195] = ~(t[160] ^ t[206]);
  assign t[196] = t[42] ^ t[198];
  assign t[197] = t[155] ^ t[60];
  assign t[198] = t[67] ^ t[81];
  assign t[199] = t[145] ? x[112] : x[111];
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[126] ^ t[86];
  assign t[201] = ~(t[35] ^ t[80]);
  assign t[202] = t[130] ^ t[46];
  assign t[203] = t[207] & t[208];
  assign t[204] = t[190] ? x[114] : x[113];
  assign t[205] = t[145] ? x[116] : x[115];
  assign t[206] = t[119] ^ t[64];
  assign t[207] = ~(t[105] ^ t[209]);
  assign t[208] = t[202] ^ t[172];
  assign t[209] = t[150] ^ t[130];
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[214]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[33] & t[215]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[7];
  assign t[239] = t[266] ^ x[10];
  assign t[23] = t[34] ^ t[35];
  assign t[240] = t[267] ^ x[13];
  assign t[241] = t[268] ^ x[18];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = ~(t[25] ^ t[30]);
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[51];
  assign t[253] = t[280] ^ x[54];
  assign t[254] = t[281] ^ x[57];
  assign t[255] = t[282] ^ x[62];
  assign t[256] = t[283] ^ x[65];
  assign t[257] = t[284] ^ x[68];
  assign t[258] = t[285] ^ x[79];
  assign t[259] = t[286] ^ x[82];
  assign t[25] = t[36] ^ t[37];
  assign t[260] = t[287] ^ x[85];
  assign t[261] = t[288] ^ x[92];
  assign t[262] = t[289] ^ x[99];
  assign t[263] = t[290] ^ x[102];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = t[42] ^ t[43];
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[7];
  assign t[294] = t[348] ^ x[6];
  assign t[295] = t[349] ^ x[10];
  assign t[296] = t[350] ^ x[9];
  assign t[297] = t[351] ^ x[13];
  assign t[298] = t[352] ^ x[12];
  assign t[299] = t[353] ^ x[18];
  assign t[29] = t[44] ^ t[45];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[17];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = t[46] ^ t[47];
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[51];
  assign t[322] = t[376] ^ x[50];
  assign t[323] = t[377] ^ x[54];
  assign t[324] = t[378] ^ x[53];
  assign t[325] = t[379] ^ x[57];
  assign t[326] = t[380] ^ x[56];
  assign t[327] = t[381] ^ x[62];
  assign t[328] = t[382] ^ x[61];
  assign t[329] = t[383] ^ x[65];
  assign t[32] = ~(t[50]);
  assign t[330] = t[384] ^ x[64];
  assign t[331] = t[385] ^ x[68];
  assign t[332] = t[386] ^ x[67];
  assign t[333] = t[387] ^ x[79];
  assign t[334] = t[388] ^ x[78];
  assign t[335] = t[389] ^ x[82];
  assign t[336] = t[390] ^ x[81];
  assign t[337] = t[391] ^ x[85];
  assign t[338] = t[392] ^ x[84];
  assign t[339] = t[393] ^ x[92];
  assign t[33] = ~(t[216]);
  assign t[340] = t[394] ^ x[91];
  assign t[341] = t[395] ^ x[99];
  assign t[342] = t[396] ^ x[98];
  assign t[343] = t[397] ^ x[102];
  assign t[344] = t[398] ^ x[101];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[5]);
  assign t[348] = (x[5]);
  assign t[349] = (x[8]);
  assign t[34] = ~(t[51] ^ t[52]);
  assign t[350] = (x[8]);
  assign t[351] = (x[11]);
  assign t[352] = (x[11]);
  assign t[353] = (x[16]);
  assign t[354] = (x[16]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = t[53] ^ t[54];
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = t[55] ^ t[44];
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[49]);
  assign t[376] = (x[49]);
  assign t[377] = (x[52]);
  assign t[378] = (x[52]);
  assign t[379] = (x[55]);
  assign t[37] = t[56] ^ t[57];
  assign t[380] = (x[55]);
  assign t[381] = (x[60]);
  assign t[382] = (x[60]);
  assign t[383] = (x[63]);
  assign t[384] = (x[63]);
  assign t[385] = (x[66]);
  assign t[386] = (x[66]);
  assign t[387] = (x[77]);
  assign t[388] = (x[77]);
  assign t[389] = (x[80]);
  assign t[38] = t[58] ^ t[34];
  assign t[390] = (x[80]);
  assign t[391] = (x[83]);
  assign t[392] = (x[83]);
  assign t[393] = (x[90]);
  assign t[394] = (x[90]);
  assign t[395] = (x[97]);
  assign t[396] = (x[97]);
  assign t[397] = (x[100]);
  assign t[398] = (x[100]);
  assign t[39] = ~(t[29] ^ t[59]);
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = t[62] ^ t[63];
  assign t[42] = t[64] ^ t[65];
  assign t[43] = t[66] & t[67];
  assign t[44] = ~t[68];
  assign t[45] = t[56] ^ t[69];
  assign t[46] = t[9] ? t[70] : t[217];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[218] | t[75];
  assign t[4] = t[9] ? t[10] : t[210];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = ~(t[79] ^ t[80]);
  assign t[53] = t[64] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = ~t[84];
  assign t[56] = t[85] ^ t[86];
  assign t[57] = t[87] & t[88];
  assign t[58] = ~(t[89] ^ t[90]);
  assign t[59] = t[91] ^ t[72];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[211] ^ t[92];
  assign t[61] = t[215] ^ t[93];
  assign t[62] = t[94] ^ t[95];
  assign t[63] = t[96] & t[97];
  assign t[64] = t[31] ? t[98] : t[219];
  assign t[65] = t[31] ? t[99] : t[220];
  assign t[66] = ~(t[81]);
  assign t[67] = t[31] ? t[100] : t[221];
  assign t[68] = t[9] ? t[101] : t[222];
  assign t[69] = t[102] & t[103];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[217] ^ t[104];
  assign t[71] = t[105] ^ t[106];
  assign t[72] = t[107] & t[108];
  assign t[73] = ~(t[75] & t[109]);
  assign t[74] = ~(t[223] ^ t[110]);
  assign t[75] = ~(t[111] & t[112]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[113] ^ t[95];
  assign t[78] = t[114] ^ t[69];
  assign t[79] = t[115] ^ t[59];
  assign t[7] = ~(t[15] ^ t[16]);
  assign t[80] = t[61] ^ t[116];
  assign t[81] = t[31] ? t[117] : t[224];
  assign t[82] = ~(t[53] ^ t[118]);
  assign t[83] = t[119] ^ t[67];
  assign t[84] = t[9] ? t[120] : t[225];
  assign t[85] = t[121] & t[122];
  assign t[86] = t[123] & t[124];
  assign t[87] = ~(t[85] ^ t[125]);
  assign t[88] = t[126] ^ t[127];
  assign t[89] = t[128] ^ t[28];
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = ~(t[129] ^ t[78]);
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[132] ? t[133] : t[226];
  assign t[93] = t[132] ? t[134] : t[227];
  assign t[94] = t[135] & t[136];
  assign t[95] = t[137] & t[138];
  assign t[96] = ~(t[94] ^ t[139]);
  assign t[97] = t[113] ^ t[140];
  assign t[98] = t[219] ^ t[141];
  assign t[99] = t[220] ^ t[142];
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [116:0] x;
 output y;

 wire [407:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[142] ^ t[143];
  assign t[101] = t[128] ^ t[59];
  assign t[102] = t[43] ^ t[84];
  assign t[103] = t[144] ^ t[145];
  assign t[104] = t[31] ? t[146] : t[234];
  assign t[105] = ~(t[69] ^ t[96]);
  assign t[106] = t[64] ^ t[147];
  assign t[107] = t[228] ^ t[148];
  assign t[108] = t[149] ^ t[63];
  assign t[109] = t[150] & t[151];
  assign t[10] = t[219] ^ t[20];
  assign t[110] = ~(t[152] & t[153]);
  assign t[111] = t[154] ^ t[235];
  assign t[112] = ~(t[229]);
  assign t[113] = t[155] & t[154];
  assign t[114] = t[156];
  assign t[115] = ~(t[81]);
  assign t[116] = t[157];
  assign t[117] = t[9] ? t[158] : t[236];
  assign t[118] = t[159] & t[160];
  assign t[119] = t[9] ? t[161] : t[237];
  assign t[11] = ~(t[220]);
  assign t[120] = ~(t[86] ^ t[162]);
  assign t[121] = t[77] ^ t[163];
  assign t[122] = t[26] ^ t[164];
  assign t[123] = ~(t[98] ^ t[101]);
  assign t[124] = t[91] ^ t[117];
  assign t[125] = t[165] ? x[62] : x[61];
  assign t[126] = ~(t[163]);
  assign t[127] = ~(t[114]);
  assign t[128] = t[114] ^ t[81];
  assign t[129] = t[166] ^ t[144];
  assign t[12] = ~(t[221]);
  assign t[130] = t[167] ^ t[168];
  assign t[131] = t[230] ^ t[169];
  assign t[132] = t[231] ^ t[170];
  assign t[133] = t[232] ^ t[171];
  assign t[134] = t[233] ^ t[172];
  assign t[135] = t[173] & t[174];
  assign t[136] = t[175] & t[147];
  assign t[137] = ~(t[135] ^ t[176]);
  assign t[138] = t[177] ^ t[178];
  assign t[139] = t[95] ^ t[179];
  assign t[13] = ~(t[222]);
  assign t[140] = t[180] ^ t[166];
  assign t[141] = t[181] & t[182];
  assign t[142] = t[180] ^ t[144];
  assign t[143] = t[183] & t[184];
  assign t[144] = t[224] ^ t[185];
  assign t[145] = t[167] ^ t[141];
  assign t[146] = t[234] ^ t[186];
  assign t[147] = t[31] ? t[187] : t[238];
  assign t[148] = t[165] ? x[67] : x[66];
  assign t[149] = t[188] & t[189];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = ~(t[124] ^ t[108]);
  assign t[151] = t[79] ^ t[93];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[190] | t[112]);
  assign t[154] = ~(t[239]);
  assign t[155] = ~(t[235]);
  assign t[156] = t[9] ? t[191] : t[240];
  assign t[157] = t[31] ? t[192] : t[241];
  assign t[158] = t[236] ^ t[193];
  assign t[159] = ~(t[149] ^ t[194]);
  assign t[15] = t[23] ^ t[24];
  assign t[160] = t[62] ^ t[195];
  assign t[161] = t[237] ^ t[196];
  assign t[162] = t[53] ^ t[114];
  assign t[163] = t[116] ^ t[81];
  assign t[164] = t[177] ^ t[136];
  assign t[165] = ~(t[50]);
  assign t[166] = t[220] ^ t[197];
  assign t[167] = t[198] ^ t[143];
  assign t[168] = t[199] & t[200];
  assign t[169] = t[165] ? x[78] : x[77];
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = t[165] ? x[80] : x[79];
  assign t[171] = t[32] ? x[82] : x[81];
  assign t[172] = t[76] ? x[84] : x[83];
  assign t[173] = ~(t[178]);
  assign t[174] = ~(t[104]);
  assign t[175] = ~(t[94]);
  assign t[176] = t[64] ^ t[104];
  assign t[177] = t[104] ^ t[95];
  assign t[178] = t[147] ^ t[94];
  assign t[179] = t[96] ^ t[70];
  assign t[17] = ~(t[27] ^ t[28]);
  assign t[180] = t[201] ? t[202] : t[242];
  assign t[181] = ~(t[140] ^ t[167]);
  assign t[182] = t[129] ^ t[184];
  assign t[183] = ~(t[166]);
  assign t[184] = t[221] ^ t[203];
  assign t[185] = t[201] ? t[204] : t[243];
  assign t[186] = t[32] ? x[92] : x[91];
  assign t[187] = t[238] ^ t[205];
  assign t[188] = ~(t[195]);
  assign t[189] = ~(t[91]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[190] = ~(t[226]);
  assign t[191] = t[240] ^ t[206];
  assign t[192] = t[241] ^ t[207];
  assign t[193] = t[165] ? x[94] : x[93];
  assign t[194] = t[79] ^ t[91];
  assign t[195] = t[93] ^ t[117];
  assign t[196] = t[165] ? x[96] : x[95];
  assign t[197] = t[201] ? t[208] : t[244];
  assign t[198] = t[209] & t[210];
  assign t[199] = ~(t[198] ^ t[211]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[142] ^ t[212];
  assign t[201] = ~(t[19]);
  assign t[202] = t[242] ^ t[213];
  assign t[203] = t[201] ? t[214] : t[245];
  assign t[204] = t[243] ^ t[215];
  assign t[205] = t[76] ? x[104] : x[103];
  assign t[206] = t[165] ? x[106] : x[105];
  assign t[207] = t[165] ? x[108] : x[107];
  assign t[208] = t[244] ^ t[216];
  assign t[209] = ~(t[212]);
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = ~(t[180]);
  assign t[211] = t[129] ^ t[180];
  assign t[212] = t[184] ^ t[166];
  assign t[213] = t[217] ? x[110] : x[109];
  assign t[214] = t[245] ^ t[218];
  assign t[215] = t[217] ? x[112] : x[111];
  assign t[216] = t[217] ? x[114] : x[113];
  assign t[217] = ~(t[50]);
  assign t[218] = t[217] ? x[116] : x[115];
  assign t[219] = (t[246]);
  assign t[21] = ~(t[223]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[33] & t[224]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = (t[266]);
  assign t[23] = ~(t[34] ^ t[35]);
  assign t[240] = (t[267]);
  assign t[241] = (t[268]);
  assign t[242] = (t[269]);
  assign t[243] = (t[270]);
  assign t[244] = (t[271]);
  assign t[245] = (t[272]);
  assign t[246] = t[273] ^ x[4];
  assign t[247] = t[274] ^ x[7];
  assign t[248] = t[275] ^ x[10];
  assign t[249] = t[276] ^ x[13];
  assign t[24] = t[36] ^ t[37];
  assign t[250] = t[277] ^ x[18];
  assign t[251] = t[278] ^ x[21];
  assign t[252] = t[279] ^ x[24];
  assign t[253] = t[280] ^ x[27];
  assign t[254] = t[281] ^ x[30];
  assign t[255] = t[282] ^ x[33];
  assign t[256] = t[283] ^ x[36];
  assign t[257] = t[284] ^ x[39];
  assign t[258] = t[285] ^ x[42];
  assign t[259] = t[286] ^ x[45];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[287] ^ x[48];
  assign t[261] = t[288] ^ x[51];
  assign t[262] = t[289] ^ x[54];
  assign t[263] = t[290] ^ x[57];
  assign t[264] = t[291] ^ x[60];
  assign t[265] = t[292] ^ x[65];
  assign t[266] = t[293] ^ x[70];
  assign t[267] = t[294] ^ x[73];
  assign t[268] = t[295] ^ x[76];
  assign t[269] = t[296] ^ x[87];
  assign t[26] = ~(t[40] ^ t[41]);
  assign t[270] = t[297] ^ x[90];
  assign t[271] = t[298] ^ x[99];
  assign t[272] = t[299] ^ x[102];
  assign t[273] = (t[300] & ~t[301]);
  assign t[274] = (t[302] & ~t[303]);
  assign t[275] = (t[304] & ~t[305]);
  assign t[276] = (t[306] & ~t[307]);
  assign t[277] = (t[308] & ~t[309]);
  assign t[278] = (t[310] & ~t[311]);
  assign t[279] = (t[312] & ~t[313]);
  assign t[27] = t[42] ^ t[43];
  assign t[280] = (t[314] & ~t[315]);
  assign t[281] = (t[316] & ~t[317]);
  assign t[282] = (t[318] & ~t[319]);
  assign t[283] = (t[320] & ~t[321]);
  assign t[284] = (t[322] & ~t[323]);
  assign t[285] = (t[324] & ~t[325]);
  assign t[286] = (t[326] & ~t[327]);
  assign t[287] = (t[328] & ~t[329]);
  assign t[288] = (t[330] & ~t[331]);
  assign t[289] = (t[332] & ~t[333]);
  assign t[28] = ~(t[44] ^ t[25]);
  assign t[290] = (t[334] & ~t[335]);
  assign t[291] = (t[336] & ~t[337]);
  assign t[292] = (t[338] & ~t[339]);
  assign t[293] = (t[340] & ~t[341]);
  assign t[294] = (t[342] & ~t[343]);
  assign t[295] = (t[344] & ~t[345]);
  assign t[296] = (t[346] & ~t[347]);
  assign t[297] = (t[348] & ~t[349]);
  assign t[298] = (t[350] & ~t[351]);
  assign t[299] = (t[352] & ~t[353]);
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[4];
  assign t[301] = t[355] ^ x[3];
  assign t[302] = t[356] ^ x[7];
  assign t[303] = t[357] ^ x[6];
  assign t[304] = t[358] ^ x[10];
  assign t[305] = t[359] ^ x[9];
  assign t[306] = t[360] ^ x[13];
  assign t[307] = t[361] ^ x[12];
  assign t[308] = t[362] ^ x[18];
  assign t[309] = t[363] ^ x[17];
  assign t[30] = ~(t[36] ^ t[47]);
  assign t[310] = t[364] ^ x[21];
  assign t[311] = t[365] ^ x[20];
  assign t[312] = t[366] ^ x[24];
  assign t[313] = t[367] ^ x[23];
  assign t[314] = t[368] ^ x[27];
  assign t[315] = t[369] ^ x[26];
  assign t[316] = t[370] ^ x[30];
  assign t[317] = t[371] ^ x[29];
  assign t[318] = t[372] ^ x[33];
  assign t[319] = t[373] ^ x[32];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[36];
  assign t[321] = t[375] ^ x[35];
  assign t[322] = t[376] ^ x[39];
  assign t[323] = t[377] ^ x[38];
  assign t[324] = t[378] ^ x[42];
  assign t[325] = t[379] ^ x[41];
  assign t[326] = t[380] ^ x[45];
  assign t[327] = t[381] ^ x[44];
  assign t[328] = t[382] ^ x[48];
  assign t[329] = t[383] ^ x[47];
  assign t[32] = ~(t[50]);
  assign t[330] = t[384] ^ x[51];
  assign t[331] = t[385] ^ x[50];
  assign t[332] = t[386] ^ x[54];
  assign t[333] = t[387] ^ x[53];
  assign t[334] = t[388] ^ x[57];
  assign t[335] = t[389] ^ x[56];
  assign t[336] = t[390] ^ x[60];
  assign t[337] = t[391] ^ x[59];
  assign t[338] = t[392] ^ x[65];
  assign t[339] = t[393] ^ x[64];
  assign t[33] = ~(t[225]);
  assign t[340] = t[394] ^ x[70];
  assign t[341] = t[395] ^ x[69];
  assign t[342] = t[396] ^ x[73];
  assign t[343] = t[397] ^ x[72];
  assign t[344] = t[398] ^ x[76];
  assign t[345] = t[399] ^ x[75];
  assign t[346] = t[400] ^ x[87];
  assign t[347] = t[401] ^ x[86];
  assign t[348] = t[402] ^ x[90];
  assign t[349] = t[403] ^ x[89];
  assign t[34] = t[51] ^ t[18];
  assign t[350] = t[404] ^ x[99];
  assign t[351] = t[405] ^ x[98];
  assign t[352] = t[406] ^ x[102];
  assign t[353] = t[407] ^ x[101];
  assign t[354] = (x[2]);
  assign t[355] = (x[2]);
  assign t[356] = (x[5]);
  assign t[357] = (x[5]);
  assign t[358] = (x[8]);
  assign t[359] = (x[8]);
  assign t[35] = ~(t[52] ^ t[44]);
  assign t[360] = (x[11]);
  assign t[361] = (x[11]);
  assign t[362] = (x[16]);
  assign t[363] = (x[16]);
  assign t[364] = (x[19]);
  assign t[365] = (x[19]);
  assign t[366] = (x[22]);
  assign t[367] = (x[22]);
  assign t[368] = (x[25]);
  assign t[369] = (x[25]);
  assign t[36] = t[53] ^ t[54];
  assign t[370] = (x[28]);
  assign t[371] = (x[28]);
  assign t[372] = (x[31]);
  assign t[373] = (x[31]);
  assign t[374] = (x[34]);
  assign t[375] = (x[34]);
  assign t[376] = (x[37]);
  assign t[377] = (x[37]);
  assign t[378] = (x[40]);
  assign t[379] = (x[40]);
  assign t[37] = ~(t[55] ^ t[56]);
  assign t[380] = (x[43]);
  assign t[381] = (x[43]);
  assign t[382] = (x[46]);
  assign t[383] = (x[46]);
  assign t[384] = (x[49]);
  assign t[385] = (x[49]);
  assign t[386] = (x[52]);
  assign t[387] = (x[52]);
  assign t[388] = (x[55]);
  assign t[389] = (x[55]);
  assign t[38] = ~t[57];
  assign t[390] = (x[58]);
  assign t[391] = (x[58]);
  assign t[392] = (x[63]);
  assign t[393] = (x[63]);
  assign t[394] = (x[68]);
  assign t[395] = (x[68]);
  assign t[396] = (x[71]);
  assign t[397] = (x[71]);
  assign t[398] = (x[74]);
  assign t[399] = (x[74]);
  assign t[39] = t[58] ^ t[59];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[400] = (x[85]);
  assign t[401] = (x[85]);
  assign t[402] = (x[88]);
  assign t[403] = (x[88]);
  assign t[404] = (x[97]);
  assign t[405] = (x[97]);
  assign t[406] = (x[100]);
  assign t[407] = (x[100]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[42] ^ t[47]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] ^ t[36]);
  assign t[45] = ~(t[67] ^ t[68]);
  assign t[46] = t[69] ^ t[70];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[226] | t[75];
  assign t[4] = t[9] ? t[10] : t[219];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] ^ t[38];
  assign t[54] = t[58] ^ t[82];
  assign t[55] = t[83] ^ t[45];
  assign t[56] = ~(t[25] ^ t[84]);
  assign t[57] = t[9] ? t[85] : t[227];
  assign t[58] = t[86] ^ t[78];
  assign t[59] = t[87] & t[88];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[25] ^ t[51];
  assign t[61] = ~(t[89] ^ t[90]);
  assign t[62] = t[91] ^ t[71];
  assign t[63] = t[92] & t[93];
  assign t[64] = t[94] ^ t[95];
  assign t[65] = t[96] ^ t[97];
  assign t[66] = ~(t[98] ^ t[99]);
  assign t[67] = t[100] ^ t[101];
  assign t[68] = ~(t[102] ^ t[103]);
  assign t[69] = t[104] ^ t[94];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[105] & t[106];
  assign t[71] = t[9] ? t[107] : t[228];
  assign t[72] = t[108] ^ t[109];
  assign t[73] = ~(t[75] & t[110]);
  assign t[74] = ~(t[229] ^ t[111]);
  assign t[75] = ~(t[112] & t[113]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[114] ^ t[38];
  assign t[78] = t[115] & t[116];
  assign t[79] = t[117] ^ t[71];
  assign t[7] = ~(t[15] ^ t[16]);
  assign t[80] = t[108] ^ t[118];
  assign t[81] = ~t[119];
  assign t[82] = t[120] & t[121];
  assign t[83] = ~(t[122] ^ t[123]);
  assign t[84] = t[124] ^ t[109];
  assign t[85] = t[227] ^ t[125];
  assign t[86] = t[126] & t[127];
  assign t[87] = ~(t[128] ^ t[58]);
  assign t[88] = t[53] ^ t[116];
  assign t[89] = ~(t[46] ^ t[103]);
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[9] ? t[131] : t[230];
  assign t[92] = ~(t[117]);
  assign t[93] = t[9] ? t[132] : t[231];
  assign t[94] = t[31] ? t[133] : t[232];
  assign t[95] = t[31] ? t[134] : t[233];
  assign t[96] = t[135] ^ t[136];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[52] ^ t[139];
  assign t[99] = t[140] ^ t[141];
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind131(x, y);
 input [116:0] x;
 output y;

 wire [407:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[142] ^ t[143];
  assign t[101] = t[128] ^ t[59];
  assign t[102] = t[43] ^ t[84];
  assign t[103] = t[144] ^ t[145];
  assign t[104] = t[31] ? t[146] : t[234];
  assign t[105] = ~(t[69] ^ t[96]);
  assign t[106] = t[64] ^ t[147];
  assign t[107] = t[228] ^ t[148];
  assign t[108] = t[149] ^ t[63];
  assign t[109] = t[150] & t[151];
  assign t[10] = t[219] ^ t[20];
  assign t[110] = ~(t[152] & t[153]);
  assign t[111] = t[154] ^ t[235];
  assign t[112] = ~(t[229]);
  assign t[113] = t[155] & t[154];
  assign t[114] = t[156];
  assign t[115] = ~(t[81]);
  assign t[116] = t[157];
  assign t[117] = t[9] ? t[158] : t[236];
  assign t[118] = t[159] & t[160];
  assign t[119] = t[9] ? t[161] : t[237];
  assign t[11] = ~(t[220]);
  assign t[120] = ~(t[86] ^ t[162]);
  assign t[121] = t[77] ^ t[163];
  assign t[122] = t[26] ^ t[164];
  assign t[123] = ~(t[98] ^ t[101]);
  assign t[124] = t[91] ^ t[117];
  assign t[125] = t[165] ? x[62] : x[61];
  assign t[126] = ~(t[163]);
  assign t[127] = ~(t[114]);
  assign t[128] = t[114] ^ t[81];
  assign t[129] = t[166] ^ t[144];
  assign t[12] = ~(t[221]);
  assign t[130] = t[167] ^ t[168];
  assign t[131] = t[230] ^ t[169];
  assign t[132] = t[231] ^ t[170];
  assign t[133] = t[232] ^ t[171];
  assign t[134] = t[233] ^ t[172];
  assign t[135] = t[173] & t[174];
  assign t[136] = t[175] & t[147];
  assign t[137] = ~(t[135] ^ t[176]);
  assign t[138] = t[177] ^ t[178];
  assign t[139] = t[95] ^ t[179];
  assign t[13] = ~(t[222]);
  assign t[140] = t[180] ^ t[166];
  assign t[141] = t[181] & t[182];
  assign t[142] = t[180] ^ t[144];
  assign t[143] = t[183] & t[184];
  assign t[144] = t[224] ^ t[185];
  assign t[145] = t[167] ^ t[141];
  assign t[146] = t[234] ^ t[186];
  assign t[147] = t[31] ? t[187] : t[238];
  assign t[148] = t[165] ? x[67] : x[66];
  assign t[149] = t[188] & t[189];
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = ~(t[124] ^ t[108]);
  assign t[151] = t[79] ^ t[93];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[190] | t[112]);
  assign t[154] = ~(t[239]);
  assign t[155] = ~(t[235]);
  assign t[156] = t[9] ? t[191] : t[240];
  assign t[157] = t[31] ? t[192] : t[241];
  assign t[158] = t[236] ^ t[193];
  assign t[159] = ~(t[149] ^ t[194]);
  assign t[15] = t[23] ^ t[24];
  assign t[160] = t[62] ^ t[195];
  assign t[161] = t[237] ^ t[196];
  assign t[162] = t[53] ^ t[114];
  assign t[163] = t[116] ^ t[81];
  assign t[164] = t[177] ^ t[136];
  assign t[165] = ~(t[50]);
  assign t[166] = t[220] ^ t[197];
  assign t[167] = t[198] ^ t[143];
  assign t[168] = t[199] & t[200];
  assign t[169] = t[165] ? x[78] : x[77];
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = t[165] ? x[80] : x[79];
  assign t[171] = t[32] ? x[82] : x[81];
  assign t[172] = t[76] ? x[84] : x[83];
  assign t[173] = ~(t[178]);
  assign t[174] = ~(t[104]);
  assign t[175] = ~(t[94]);
  assign t[176] = t[64] ^ t[104];
  assign t[177] = t[104] ^ t[95];
  assign t[178] = t[147] ^ t[94];
  assign t[179] = t[96] ^ t[70];
  assign t[17] = ~(t[27] ^ t[28]);
  assign t[180] = t[201] ? t[202] : t[242];
  assign t[181] = ~(t[140] ^ t[167]);
  assign t[182] = t[129] ^ t[184];
  assign t[183] = ~(t[166]);
  assign t[184] = t[221] ^ t[203];
  assign t[185] = t[201] ? t[204] : t[243];
  assign t[186] = t[32] ? x[92] : x[91];
  assign t[187] = t[238] ^ t[205];
  assign t[188] = ~(t[195]);
  assign t[189] = ~(t[91]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[190] = ~(t[226]);
  assign t[191] = t[240] ^ t[206];
  assign t[192] = t[241] ^ t[207];
  assign t[193] = t[165] ? x[94] : x[93];
  assign t[194] = t[79] ^ t[91];
  assign t[195] = t[93] ^ t[117];
  assign t[196] = t[165] ? x[96] : x[95];
  assign t[197] = t[201] ? t[208] : t[244];
  assign t[198] = t[209] & t[210];
  assign t[199] = ~(t[198] ^ t[211]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[142] ^ t[212];
  assign t[201] = ~(t[19]);
  assign t[202] = t[242] ^ t[213];
  assign t[203] = t[201] ? t[214] : t[245];
  assign t[204] = t[243] ^ t[215];
  assign t[205] = t[76] ? x[104] : x[103];
  assign t[206] = t[165] ? x[106] : x[105];
  assign t[207] = t[165] ? x[108] : x[107];
  assign t[208] = t[244] ^ t[216];
  assign t[209] = ~(t[212]);
  assign t[20] = t[32] ? x[15] : x[14];
  assign t[210] = ~(t[180]);
  assign t[211] = t[129] ^ t[180];
  assign t[212] = t[184] ^ t[166];
  assign t[213] = t[217] ? x[110] : x[109];
  assign t[214] = t[245] ^ t[218];
  assign t[215] = t[217] ? x[112] : x[111];
  assign t[216] = t[217] ? x[114] : x[113];
  assign t[217] = ~(t[50]);
  assign t[218] = t[217] ? x[116] : x[115];
  assign t[219] = (t[246]);
  assign t[21] = ~(t[223]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[33] & t[224]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = (t[266]);
  assign t[23] = ~(t[34] ^ t[35]);
  assign t[240] = (t[267]);
  assign t[241] = (t[268]);
  assign t[242] = (t[269]);
  assign t[243] = (t[270]);
  assign t[244] = (t[271]);
  assign t[245] = (t[272]);
  assign t[246] = t[273] ^ x[4];
  assign t[247] = t[274] ^ x[7];
  assign t[248] = t[275] ^ x[10];
  assign t[249] = t[276] ^ x[13];
  assign t[24] = t[36] ^ t[37];
  assign t[250] = t[277] ^ x[18];
  assign t[251] = t[278] ^ x[21];
  assign t[252] = t[279] ^ x[24];
  assign t[253] = t[280] ^ x[27];
  assign t[254] = t[281] ^ x[30];
  assign t[255] = t[282] ^ x[33];
  assign t[256] = t[283] ^ x[36];
  assign t[257] = t[284] ^ x[39];
  assign t[258] = t[285] ^ x[42];
  assign t[259] = t[286] ^ x[45];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[287] ^ x[48];
  assign t[261] = t[288] ^ x[51];
  assign t[262] = t[289] ^ x[54];
  assign t[263] = t[290] ^ x[57];
  assign t[264] = t[291] ^ x[60];
  assign t[265] = t[292] ^ x[65];
  assign t[266] = t[293] ^ x[70];
  assign t[267] = t[294] ^ x[73];
  assign t[268] = t[295] ^ x[76];
  assign t[269] = t[296] ^ x[87];
  assign t[26] = ~(t[40] ^ t[41]);
  assign t[270] = t[297] ^ x[90];
  assign t[271] = t[298] ^ x[99];
  assign t[272] = t[299] ^ x[102];
  assign t[273] = (t[300] & ~t[301]);
  assign t[274] = (t[302] & ~t[303]);
  assign t[275] = (t[304] & ~t[305]);
  assign t[276] = (t[306] & ~t[307]);
  assign t[277] = (t[308] & ~t[309]);
  assign t[278] = (t[310] & ~t[311]);
  assign t[279] = (t[312] & ~t[313]);
  assign t[27] = t[42] ^ t[43];
  assign t[280] = (t[314] & ~t[315]);
  assign t[281] = (t[316] & ~t[317]);
  assign t[282] = (t[318] & ~t[319]);
  assign t[283] = (t[320] & ~t[321]);
  assign t[284] = (t[322] & ~t[323]);
  assign t[285] = (t[324] & ~t[325]);
  assign t[286] = (t[326] & ~t[327]);
  assign t[287] = (t[328] & ~t[329]);
  assign t[288] = (t[330] & ~t[331]);
  assign t[289] = (t[332] & ~t[333]);
  assign t[28] = ~(t[44] ^ t[25]);
  assign t[290] = (t[334] & ~t[335]);
  assign t[291] = (t[336] & ~t[337]);
  assign t[292] = (t[338] & ~t[339]);
  assign t[293] = (t[340] & ~t[341]);
  assign t[294] = (t[342] & ~t[343]);
  assign t[295] = (t[344] & ~t[345]);
  assign t[296] = (t[346] & ~t[347]);
  assign t[297] = (t[348] & ~t[349]);
  assign t[298] = (t[350] & ~t[351]);
  assign t[299] = (t[352] & ~t[353]);
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[5] | t[6]);
  assign t[300] = t[354] ^ x[4];
  assign t[301] = t[355] ^ x[3];
  assign t[302] = t[356] ^ x[7];
  assign t[303] = t[357] ^ x[6];
  assign t[304] = t[358] ^ x[10];
  assign t[305] = t[359] ^ x[9];
  assign t[306] = t[360] ^ x[13];
  assign t[307] = t[361] ^ x[12];
  assign t[308] = t[362] ^ x[18];
  assign t[309] = t[363] ^ x[17];
  assign t[30] = ~(t[36] ^ t[47]);
  assign t[310] = t[364] ^ x[21];
  assign t[311] = t[365] ^ x[20];
  assign t[312] = t[366] ^ x[24];
  assign t[313] = t[367] ^ x[23];
  assign t[314] = t[368] ^ x[27];
  assign t[315] = t[369] ^ x[26];
  assign t[316] = t[370] ^ x[30];
  assign t[317] = t[371] ^ x[29];
  assign t[318] = t[372] ^ x[33];
  assign t[319] = t[373] ^ x[32];
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = t[374] ^ x[36];
  assign t[321] = t[375] ^ x[35];
  assign t[322] = t[376] ^ x[39];
  assign t[323] = t[377] ^ x[38];
  assign t[324] = t[378] ^ x[42];
  assign t[325] = t[379] ^ x[41];
  assign t[326] = t[380] ^ x[45];
  assign t[327] = t[381] ^ x[44];
  assign t[328] = t[382] ^ x[48];
  assign t[329] = t[383] ^ x[47];
  assign t[32] = ~(t[50]);
  assign t[330] = t[384] ^ x[51];
  assign t[331] = t[385] ^ x[50];
  assign t[332] = t[386] ^ x[54];
  assign t[333] = t[387] ^ x[53];
  assign t[334] = t[388] ^ x[57];
  assign t[335] = t[389] ^ x[56];
  assign t[336] = t[390] ^ x[60];
  assign t[337] = t[391] ^ x[59];
  assign t[338] = t[392] ^ x[65];
  assign t[339] = t[393] ^ x[64];
  assign t[33] = ~(t[225]);
  assign t[340] = t[394] ^ x[70];
  assign t[341] = t[395] ^ x[69];
  assign t[342] = t[396] ^ x[73];
  assign t[343] = t[397] ^ x[72];
  assign t[344] = t[398] ^ x[76];
  assign t[345] = t[399] ^ x[75];
  assign t[346] = t[400] ^ x[87];
  assign t[347] = t[401] ^ x[86];
  assign t[348] = t[402] ^ x[90];
  assign t[349] = t[403] ^ x[89];
  assign t[34] = t[51] ^ t[18];
  assign t[350] = t[404] ^ x[99];
  assign t[351] = t[405] ^ x[98];
  assign t[352] = t[406] ^ x[102];
  assign t[353] = t[407] ^ x[101];
  assign t[354] = (x[2]);
  assign t[355] = (x[2]);
  assign t[356] = (x[5]);
  assign t[357] = (x[5]);
  assign t[358] = (x[8]);
  assign t[359] = (x[8]);
  assign t[35] = ~(t[52] ^ t[44]);
  assign t[360] = (x[11]);
  assign t[361] = (x[11]);
  assign t[362] = (x[16]);
  assign t[363] = (x[16]);
  assign t[364] = (x[19]);
  assign t[365] = (x[19]);
  assign t[366] = (x[22]);
  assign t[367] = (x[22]);
  assign t[368] = (x[25]);
  assign t[369] = (x[25]);
  assign t[36] = t[53] ^ t[54];
  assign t[370] = (x[28]);
  assign t[371] = (x[28]);
  assign t[372] = (x[31]);
  assign t[373] = (x[31]);
  assign t[374] = (x[34]);
  assign t[375] = (x[34]);
  assign t[376] = (x[37]);
  assign t[377] = (x[37]);
  assign t[378] = (x[40]);
  assign t[379] = (x[40]);
  assign t[37] = ~(t[55] ^ t[56]);
  assign t[380] = (x[43]);
  assign t[381] = (x[43]);
  assign t[382] = (x[46]);
  assign t[383] = (x[46]);
  assign t[384] = (x[49]);
  assign t[385] = (x[49]);
  assign t[386] = (x[52]);
  assign t[387] = (x[52]);
  assign t[388] = (x[55]);
  assign t[389] = (x[55]);
  assign t[38] = ~t[57];
  assign t[390] = (x[58]);
  assign t[391] = (x[58]);
  assign t[392] = (x[63]);
  assign t[393] = (x[63]);
  assign t[394] = (x[68]);
  assign t[395] = (x[68]);
  assign t[396] = (x[71]);
  assign t[397] = (x[71]);
  assign t[398] = (x[74]);
  assign t[399] = (x[74]);
  assign t[39] = t[58] ^ t[59];
  assign t[3] = ~(t[7] ^ t[8]);
  assign t[400] = (x[85]);
  assign t[401] = (x[85]);
  assign t[402] = (x[88]);
  assign t[403] = (x[88]);
  assign t[404] = (x[97]);
  assign t[405] = (x[97]);
  assign t[406] = (x[100]);
  assign t[407] = (x[100]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[42] ^ t[47]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] ^ t[36]);
  assign t[45] = ~(t[67] ^ t[68]);
  assign t[46] = t[69] ^ t[70];
  assign t[47] = t[71] ^ t[72];
  assign t[48] = ~(t[73] & t[74]);
  assign t[49] = t[226] | t[75];
  assign t[4] = t[9] ? t[10] : t[219];
  assign t[50] = ~(t[76]);
  assign t[51] = t[77] ^ t[78];
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] ^ t[38];
  assign t[54] = t[58] ^ t[82];
  assign t[55] = t[83] ^ t[45];
  assign t[56] = ~(t[25] ^ t[84]);
  assign t[57] = t[9] ? t[85] : t[227];
  assign t[58] = t[86] ^ t[78];
  assign t[59] = t[87] & t[88];
  assign t[5] = ~(t[11] & t[12]);
  assign t[60] = t[25] ^ t[51];
  assign t[61] = ~(t[89] ^ t[90]);
  assign t[62] = t[91] ^ t[71];
  assign t[63] = t[92] & t[93];
  assign t[64] = t[94] ^ t[95];
  assign t[65] = t[96] ^ t[97];
  assign t[66] = ~(t[98] ^ t[99]);
  assign t[67] = t[100] ^ t[101];
  assign t[68] = ~(t[102] ^ t[103]);
  assign t[69] = t[104] ^ t[94];
  assign t[6] = ~(t[13] & t[14]);
  assign t[70] = t[105] & t[106];
  assign t[71] = t[9] ? t[107] : t[228];
  assign t[72] = t[108] ^ t[109];
  assign t[73] = ~(t[75] & t[110]);
  assign t[74] = ~(t[229] ^ t[111]);
  assign t[75] = ~(t[112] & t[113]);
  assign t[76] = ~(t[49]);
  assign t[77] = t[114] ^ t[38];
  assign t[78] = t[115] & t[116];
  assign t[79] = t[117] ^ t[71];
  assign t[7] = ~(t[15] ^ t[16]);
  assign t[80] = t[108] ^ t[118];
  assign t[81] = ~t[119];
  assign t[82] = t[120] & t[121];
  assign t[83] = ~(t[122] ^ t[123]);
  assign t[84] = t[124] ^ t[109];
  assign t[85] = t[227] ^ t[125];
  assign t[86] = t[126] & t[127];
  assign t[87] = ~(t[128] ^ t[58]);
  assign t[88] = t[53] ^ t[116];
  assign t[89] = ~(t[46] ^ t[103]);
  assign t[8] = ~(t[17] ^ t[18]);
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[9] ? t[131] : t[230];
  assign t[92] = ~(t[117]);
  assign t[93] = t[9] ? t[132] : t[231];
  assign t[94] = t[31] ? t[133] : t[232];
  assign t[95] = t[31] ? t[134] : t[233];
  assign t[96] = t[135] ^ t[136];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[52] ^ t[139];
  assign t[99] = t[140] ^ t[141];
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [116:0] x;
 output y;

 wire [400:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[8] ? t[140] : t[225];
  assign t[101] = t[141] ^ t[105];
  assign t[102] = t[142] & t[143];
  assign t[103] = t[220] ^ t[144];
  assign t[104] = t[123] ^ t[67];
  assign t[105] = t[145] & t[146];
  assign t[106] = ~t[147];
  assign t[107] = t[119] ^ t[54];
  assign t[108] = t[148] ^ t[121];
  assign t[109] = ~(t[149] & t[150]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[151] ^ t[226];
  assign t[111] = ~(t[221]);
  assign t[112] = t[152] & t[151];
  assign t[113] = ~(t[15]);
  assign t[114] = t[223] ^ t[153];
  assign t[115] = t[213] ^ t[154];
  assign t[116] = t[113] ? t[155] : t[227];
  assign t[117] = t[8] ? t[156] : t[228];
  assign t[118] = t[8] ? t[157] : t[229];
  assign t[119] = t[158] ^ t[159];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[160];
  assign t[121] = t[27] ? t[161] : t[230];
  assign t[122] = t[162] & t[163];
  assign t[123] = t[8] ? t[164] : t[231];
  assign t[124] = ~(t[86] ^ t[101]);
  assign t[125] = t[65] ^ t[146];
  assign t[126] = t[224] ^ t[165];
  assign t[127] = t[166] & t[167];
  assign t[128] = ~(t[135] ^ t[89]);
  assign t[129] = t[137] ^ t[79];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[75] ? x[65] : x[64];
  assign t[131] = t[168] & t[169];
  assign t[132] = t[170] & t[171];
  assign t[133] = ~(t[108] ^ t[92]);
  assign t[134] = t[84] ^ t[171];
  assign t[135] = t[77] ^ t[115];
  assign t[136] = t[172] & t[173];
  assign t[137] = t[115] ^ t[57];
  assign t[138] = t[89] ^ t[174];
  assign t[139] = t[148] ^ t[59];
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[225] ^ t[175];
  assign t[141] = t[176] & t[177];
  assign t[142] = ~(t[141] ^ t[178]);
  assign t[143] = t[104] ^ t[179];
  assign t[144] = t[180] ? x[67] : x[66];
  assign t[145] = ~(t[100]);
  assign t[146] = t[8] ? t[181] : t[232];
  assign t[147] = t[8] ? t[182] : t[233];
  assign t[148] = t[27] ? t[183] : t[234];
  assign t[149] = ~(t[152] | t[151]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[184] | t[111]);
  assign t[151] = ~(t[235]);
  assign t[152] = ~(t[226]);
  assign t[153] = t[185] ? x[81] : x[80];
  assign t[154] = t[113] ? t[186] : t[236];
  assign t[155] = t[227] ^ t[187];
  assign t[156] = t[228] ^ t[188];
  assign t[157] = t[229] ^ t[189];
  assign t[158] = t[190] & t[191];
  assign t[159] = t[192] & t[120];
  assign t[15] = ~(t[27]);
  assign t[160] = t[27] ? t[193] : t[237];
  assign t[161] = t[230] ^ t[194];
  assign t[162] = ~(t[131] ^ t[195]);
  assign t[163] = t[139] ^ t[196];
  assign t[164] = t[231] ^ t[197];
  assign t[165] = t[185] ? x[89] : x[88];
  assign t[166] = ~(t[198]);
  assign t[167] = ~(t[77]);
  assign t[168] = ~(t[196]);
  assign t[169] = ~(t[148]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[121]);
  assign t[171] = t[27] ? t[199] : t[238];
  assign t[172] = ~(t[158] ^ t[200]);
  assign t[173] = t[201] ^ t[202];
  assign t[174] = t[203] & t[204];
  assign t[175] = t[180] ? x[94] : x[93];
  assign t[176] = ~(t[179]);
  assign t[177] = ~(t[123]);
  assign t[178] = t[65] ^ t[123];
  assign t[179] = t[146] ^ t[100];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[48]);
  assign t[181] = t[232] ^ t[205];
  assign t[182] = t[233] ^ t[206];
  assign t[183] = t[234] ^ t[207];
  assign t[184] = ~(t[216]);
  assign t[185] = ~(t[48]);
  assign t[186] = t[236] ^ t[208];
  assign t[187] = t[185] ? x[96] : x[95];
  assign t[188] = t[180] ? x[98] : x[97];
  assign t[189] = t[180] ? x[100] : x[99];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = ~(t[202]);
  assign t[191] = ~(t[80]);
  assign t[192] = ~(t[81]);
  assign t[193] = t[237] ^ t[209];
  assign t[194] = t[28] ? x[102] : x[101];
  assign t[195] = t[84] ^ t[148];
  assign t[196] = t[171] ^ t[121];
  assign t[197] = t[180] ? x[104] : x[103];
  assign t[198] = t[79] ^ t[115];
  assign t[199] = t[238] ^ t[210];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[96] ^ t[80];
  assign t[201] = t[80] ^ t[106];
  assign t[202] = t[120] ^ t[81];
  assign t[203] = ~(t[127] ^ t[211]);
  assign t[204] = t[51] ^ t[198];
  assign t[205] = t[180] ? x[106] : x[105];
  assign t[206] = t[180] ? x[108] : x[107];
  assign t[207] = t[28] ? x[110] : x[109];
  assign t[208] = t[185] ? x[112] : x[111];
  assign t[209] = t[180] ? x[114] : x[113];
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = t[75] ? x[116] : x[115];
  assign t[211] = t[137] ^ t[77];
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[35]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[38] ^ t[39];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = t[266] ^ x[4];
  assign t[23] = t[22] ^ t[34];
  assign t[240] = t[267] ^ x[9];
  assign t[241] = t[268] ^ x[12];
  assign t[242] = t[269] ^ x[15];
  assign t[243] = t[270] ^ x[18];
  assign t[244] = t[271] ^ x[21];
  assign t[245] = t[272] ^ x[24];
  assign t[246] = t[273] ^ x[27];
  assign t[247] = t[274] ^ x[30];
  assign t[248] = t[275] ^ x[33];
  assign t[249] = t[276] ^ x[36];
  assign t[24] = ~(t[40] ^ t[41]);
  assign t[250] = t[277] ^ x[39];
  assign t[251] = t[278] ^ x[42];
  assign t[252] = t[279] ^ x[45];
  assign t[253] = t[280] ^ x[48];
  assign t[254] = t[281] ^ x[51];
  assign t[255] = t[282] ^ x[54];
  assign t[256] = t[283] ^ x[57];
  assign t[257] = t[284] ^ x[60];
  assign t[258] = t[285] ^ x[63];
  assign t[259] = t[286] ^ x[70];
  assign t[25] = ~(t[42] ^ t[43]);
  assign t[260] = t[287] ^ x[73];
  assign t[261] = t[288] ^ x[76];
  assign t[262] = t[289] ^ x[79];
  assign t[263] = t[290] ^ x[84];
  assign t[264] = t[291] ^ x[87];
  assign t[265] = t[292] ^ x[92];
  assign t[266] = (t[293] & ~t[294]);
  assign t[267] = (t[295] & ~t[296]);
  assign t[268] = (t[297] & ~t[298]);
  assign t[269] = (t[299] & ~t[300]);
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[270] = (t[301] & ~t[302]);
  assign t[271] = (t[303] & ~t[304]);
  assign t[272] = (t[305] & ~t[306]);
  assign t[273] = (t[307] & ~t[308]);
  assign t[274] = (t[309] & ~t[310]);
  assign t[275] = (t[311] & ~t[312]);
  assign t[276] = (t[313] & ~t[314]);
  assign t[277] = (t[315] & ~t[316]);
  assign t[278] = (t[317] & ~t[318]);
  assign t[279] = (t[319] & ~t[320]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = t[347] ^ x[4];
  assign t[294] = t[348] ^ x[3];
  assign t[295] = t[349] ^ x[9];
  assign t[296] = t[350] ^ x[8];
  assign t[297] = t[351] ^ x[12];
  assign t[298] = t[352] ^ x[11];
  assign t[299] = t[353] ^ x[15];
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[14];
  assign t[301] = t[355] ^ x[18];
  assign t[302] = t[356] ^ x[17];
  assign t[303] = t[357] ^ x[21];
  assign t[304] = t[358] ^ x[20];
  assign t[305] = t[359] ^ x[24];
  assign t[306] = t[360] ^ x[23];
  assign t[307] = t[361] ^ x[27];
  assign t[308] = t[362] ^ x[26];
  assign t[309] = t[363] ^ x[30];
  assign t[30] = ~(t[214]);
  assign t[310] = t[364] ^ x[29];
  assign t[311] = t[365] ^ x[33];
  assign t[312] = t[366] ^ x[32];
  assign t[313] = t[367] ^ x[36];
  assign t[314] = t[368] ^ x[35];
  assign t[315] = t[369] ^ x[39];
  assign t[316] = t[370] ^ x[38];
  assign t[317] = t[371] ^ x[42];
  assign t[318] = t[372] ^ x[41];
  assign t[319] = t[373] ^ x[45];
  assign t[31] = ~(t[215]);
  assign t[320] = t[374] ^ x[44];
  assign t[321] = t[375] ^ x[48];
  assign t[322] = t[376] ^ x[47];
  assign t[323] = t[377] ^ x[51];
  assign t[324] = t[378] ^ x[50];
  assign t[325] = t[379] ^ x[54];
  assign t[326] = t[380] ^ x[53];
  assign t[327] = t[381] ^ x[57];
  assign t[328] = t[382] ^ x[56];
  assign t[329] = t[383] ^ x[60];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[59];
  assign t[331] = t[385] ^ x[63];
  assign t[332] = t[386] ^ x[62];
  assign t[333] = t[387] ^ x[70];
  assign t[334] = t[388] ^ x[69];
  assign t[335] = t[389] ^ x[73];
  assign t[336] = t[390] ^ x[72];
  assign t[337] = t[391] ^ x[76];
  assign t[338] = t[392] ^ x[75];
  assign t[339] = t[393] ^ x[79];
  assign t[33] = t[51] ^ t[52];
  assign t[340] = t[394] ^ x[78];
  assign t[341] = t[395] ^ x[84];
  assign t[342] = t[396] ^ x[83];
  assign t[343] = t[397] ^ x[87];
  assign t[344] = t[398] ^ x[86];
  assign t[345] = t[399] ^ x[92];
  assign t[346] = t[400] ^ x[91];
  assign t[347] = (x[2]);
  assign t[348] = (x[2]);
  assign t[349] = (x[7]);
  assign t[34] = t[53] ^ t[54];
  assign t[350] = (x[7]);
  assign t[351] = (x[10]);
  assign t[352] = (x[10]);
  assign t[353] = (x[13]);
  assign t[354] = (x[13]);
  assign t[355] = (x[16]);
  assign t[356] = (x[16]);
  assign t[357] = (x[19]);
  assign t[358] = (x[19]);
  assign t[359] = (x[22]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[22]);
  assign t[361] = (x[25]);
  assign t[362] = (x[25]);
  assign t[363] = (x[28]);
  assign t[364] = (x[28]);
  assign t[365] = (x[31]);
  assign t[366] = (x[31]);
  assign t[367] = (x[34]);
  assign t[368] = (x[34]);
  assign t[369] = (x[37]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[37]);
  assign t[371] = (x[40]);
  assign t[372] = (x[40]);
  assign t[373] = (x[43]);
  assign t[374] = (x[43]);
  assign t[375] = (x[46]);
  assign t[376] = (x[46]);
  assign t[377] = (x[49]);
  assign t[378] = (x[49]);
  assign t[379] = (x[52]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[52]);
  assign t[381] = (x[55]);
  assign t[382] = (x[55]);
  assign t[383] = (x[58]);
  assign t[384] = (x[58]);
  assign t[385] = (x[61]);
  assign t[386] = (x[61]);
  assign t[387] = (x[68]);
  assign t[388] = (x[68]);
  assign t[389] = (x[71]);
  assign t[38] = ~(t[61] ^ t[62]);
  assign t[390] = (x[71]);
  assign t[391] = (x[74]);
  assign t[392] = (x[74]);
  assign t[393] = (x[77]);
  assign t[394] = (x[77]);
  assign t[395] = (x[82]);
  assign t[396] = (x[82]);
  assign t[397] = (x[85]);
  assign t[398] = (x[85]);
  assign t[399] = (x[90]);
  assign t[39] = ~(t[63] ^ t[64]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[90]);
  assign t[40] = t[65] ^ t[66];
  assign t[41] = t[67] ^ t[68];
  assign t[42] = t[69] ^ t[55];
  assign t[43] = ~(t[38] ^ t[70]);
  assign t[44] = t[11] ^ t[71];
  assign t[45] = ~(t[62] ^ t[41]);
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[216] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[217]);
  assign t[4] = t[8] ? t[9] : t[212];
  assign t[50] = ~(t[76] & t[218]);
  assign t[51] = t[77] ^ t[57];
  assign t[52] = t[78] & t[79];
  assign t[53] = t[80] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = t[84] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[218] ^ t[88];
  assign t[58] = t[89] ^ t[90];
  assign t[59] = t[27] ? t[91] : t[219];
  assign t[5] = ~(t[10]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = ~(t[94] ^ t[95]);
  assign t[62] = t[96] ^ t[97];
  assign t[63] = t[98] ^ t[99];
  assign t[64] = ~(t[70] ^ t[41]);
  assign t[65] = t[100] ^ t[67];
  assign t[66] = t[101] ^ t[102];
  assign t[67] = t[8] ? t[103] : t[220];
  assign t[68] = t[101] ^ t[87];
  assign t[69] = t[104] ^ t[105];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[106] ^ t[107];
  assign t[71] = t[108] ^ t[93];
  assign t[72] = ~(t[74] & t[109]);
  assign t[73] = ~(t[221] ^ t[110]);
  assign t[74] = ~(t[111] & t[112]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[222]);
  assign t[77] = t[113] ? t[114] : t[223];
  assign t[78] = ~(t[115]);
  assign t[79] = t[214] ^ t[116];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117];
  assign t[81] = ~t[118];
  assign t[82] = ~(t[53] ^ t[119]);
  assign t[83] = t[96] ^ t[120];
  assign t[84] = t[121] ^ t[59];
  assign t[85] = t[92] ^ t[122];
  assign t[86] = t[123] ^ t[100];
  assign t[87] = t[124] & t[125];
  assign t[88] = t[113] ? t[126] : t[224];
  assign t[89] = t[127] ^ t[52];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] & t[129];
  assign t[91] = t[219] ^ t[130];
  assign t[92] = t[131] ^ t[132];
  assign t[93] = t[133] & t[134];
  assign t[94] = t[40] ^ t[37];
  assign t[95] = t[135] ^ t[90];
  assign t[96] = t[81] ^ t[106];
  assign t[97] = t[119] ^ t[136];
  assign t[98] = t[137] ^ t[138];
  assign t[99] = t[139] ^ t[132];
  assign t[9] = t[212] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [116:0] x;
 output y;

 wire [400:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[8] ? t[140] : t[225];
  assign t[101] = t[141] ^ t[105];
  assign t[102] = t[142] & t[143];
  assign t[103] = t[220] ^ t[144];
  assign t[104] = t[123] ^ t[67];
  assign t[105] = t[145] & t[146];
  assign t[106] = ~t[147];
  assign t[107] = t[119] ^ t[54];
  assign t[108] = t[148] ^ t[121];
  assign t[109] = ~(t[149] & t[150]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[151] ^ t[226];
  assign t[111] = ~(t[221]);
  assign t[112] = t[152] & t[151];
  assign t[113] = ~(t[15]);
  assign t[114] = t[223] ^ t[153];
  assign t[115] = t[213] ^ t[154];
  assign t[116] = t[113] ? t[155] : t[227];
  assign t[117] = t[8] ? t[156] : t[228];
  assign t[118] = t[8] ? t[157] : t[229];
  assign t[119] = t[158] ^ t[159];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[160];
  assign t[121] = t[27] ? t[161] : t[230];
  assign t[122] = t[162] & t[163];
  assign t[123] = t[8] ? t[164] : t[231];
  assign t[124] = ~(t[86] ^ t[101]);
  assign t[125] = t[65] ^ t[146];
  assign t[126] = t[224] ^ t[165];
  assign t[127] = t[166] & t[167];
  assign t[128] = ~(t[135] ^ t[89]);
  assign t[129] = t[137] ^ t[79];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[75] ? x[65] : x[64];
  assign t[131] = t[168] & t[169];
  assign t[132] = t[170] & t[171];
  assign t[133] = ~(t[108] ^ t[92]);
  assign t[134] = t[84] ^ t[171];
  assign t[135] = t[77] ^ t[115];
  assign t[136] = t[172] & t[173];
  assign t[137] = t[115] ^ t[57];
  assign t[138] = t[89] ^ t[174];
  assign t[139] = t[148] ^ t[59];
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[225] ^ t[175];
  assign t[141] = t[176] & t[177];
  assign t[142] = ~(t[141] ^ t[178]);
  assign t[143] = t[104] ^ t[179];
  assign t[144] = t[180] ? x[67] : x[66];
  assign t[145] = ~(t[100]);
  assign t[146] = t[8] ? t[181] : t[232];
  assign t[147] = t[8] ? t[182] : t[233];
  assign t[148] = t[27] ? t[183] : t[234];
  assign t[149] = ~(t[152] | t[151]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[184] | t[111]);
  assign t[151] = ~(t[235]);
  assign t[152] = ~(t[226]);
  assign t[153] = t[185] ? x[81] : x[80];
  assign t[154] = t[113] ? t[186] : t[236];
  assign t[155] = t[227] ^ t[187];
  assign t[156] = t[228] ^ t[188];
  assign t[157] = t[229] ^ t[189];
  assign t[158] = t[190] & t[191];
  assign t[159] = t[192] & t[120];
  assign t[15] = ~(t[27]);
  assign t[160] = t[27] ? t[193] : t[237];
  assign t[161] = t[230] ^ t[194];
  assign t[162] = ~(t[131] ^ t[195]);
  assign t[163] = t[139] ^ t[196];
  assign t[164] = t[231] ^ t[197];
  assign t[165] = t[185] ? x[89] : x[88];
  assign t[166] = ~(t[198]);
  assign t[167] = ~(t[77]);
  assign t[168] = ~(t[196]);
  assign t[169] = ~(t[148]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[121]);
  assign t[171] = t[27] ? t[199] : t[238];
  assign t[172] = ~(t[158] ^ t[200]);
  assign t[173] = t[201] ^ t[202];
  assign t[174] = t[203] & t[204];
  assign t[175] = t[180] ? x[94] : x[93];
  assign t[176] = ~(t[179]);
  assign t[177] = ~(t[123]);
  assign t[178] = t[65] ^ t[123];
  assign t[179] = t[146] ^ t[100];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[48]);
  assign t[181] = t[232] ^ t[205];
  assign t[182] = t[233] ^ t[206];
  assign t[183] = t[234] ^ t[207];
  assign t[184] = ~(t[216]);
  assign t[185] = ~(t[48]);
  assign t[186] = t[236] ^ t[208];
  assign t[187] = t[185] ? x[96] : x[95];
  assign t[188] = t[180] ? x[98] : x[97];
  assign t[189] = t[180] ? x[100] : x[99];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = ~(t[202]);
  assign t[191] = ~(t[80]);
  assign t[192] = ~(t[81]);
  assign t[193] = t[237] ^ t[209];
  assign t[194] = t[28] ? x[102] : x[101];
  assign t[195] = t[84] ^ t[148];
  assign t[196] = t[171] ^ t[121];
  assign t[197] = t[180] ? x[104] : x[103];
  assign t[198] = t[79] ^ t[115];
  assign t[199] = t[238] ^ t[210];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[96] ^ t[80];
  assign t[201] = t[80] ^ t[106];
  assign t[202] = t[120] ^ t[81];
  assign t[203] = ~(t[127] ^ t[211]);
  assign t[204] = t[51] ^ t[198];
  assign t[205] = t[180] ? x[106] : x[105];
  assign t[206] = t[180] ? x[108] : x[107];
  assign t[207] = t[28] ? x[110] : x[109];
  assign t[208] = t[185] ? x[112] : x[111];
  assign t[209] = t[180] ? x[114] : x[113];
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = t[75] ? x[116] : x[115];
  assign t[211] = t[137] ^ t[77];
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[35]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[38] ^ t[39];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = t[266] ^ x[4];
  assign t[23] = t[22] ^ t[34];
  assign t[240] = t[267] ^ x[9];
  assign t[241] = t[268] ^ x[12];
  assign t[242] = t[269] ^ x[15];
  assign t[243] = t[270] ^ x[18];
  assign t[244] = t[271] ^ x[21];
  assign t[245] = t[272] ^ x[24];
  assign t[246] = t[273] ^ x[27];
  assign t[247] = t[274] ^ x[30];
  assign t[248] = t[275] ^ x[33];
  assign t[249] = t[276] ^ x[36];
  assign t[24] = ~(t[40] ^ t[41]);
  assign t[250] = t[277] ^ x[39];
  assign t[251] = t[278] ^ x[42];
  assign t[252] = t[279] ^ x[45];
  assign t[253] = t[280] ^ x[48];
  assign t[254] = t[281] ^ x[51];
  assign t[255] = t[282] ^ x[54];
  assign t[256] = t[283] ^ x[57];
  assign t[257] = t[284] ^ x[60];
  assign t[258] = t[285] ^ x[63];
  assign t[259] = t[286] ^ x[70];
  assign t[25] = ~(t[42] ^ t[43]);
  assign t[260] = t[287] ^ x[73];
  assign t[261] = t[288] ^ x[76];
  assign t[262] = t[289] ^ x[79];
  assign t[263] = t[290] ^ x[84];
  assign t[264] = t[291] ^ x[87];
  assign t[265] = t[292] ^ x[92];
  assign t[266] = (t[293] & ~t[294]);
  assign t[267] = (t[295] & ~t[296]);
  assign t[268] = (t[297] & ~t[298]);
  assign t[269] = (t[299] & ~t[300]);
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[270] = (t[301] & ~t[302]);
  assign t[271] = (t[303] & ~t[304]);
  assign t[272] = (t[305] & ~t[306]);
  assign t[273] = (t[307] & ~t[308]);
  assign t[274] = (t[309] & ~t[310]);
  assign t[275] = (t[311] & ~t[312]);
  assign t[276] = (t[313] & ~t[314]);
  assign t[277] = (t[315] & ~t[316]);
  assign t[278] = (t[317] & ~t[318]);
  assign t[279] = (t[319] & ~t[320]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = t[347] ^ x[4];
  assign t[294] = t[348] ^ x[3];
  assign t[295] = t[349] ^ x[9];
  assign t[296] = t[350] ^ x[8];
  assign t[297] = t[351] ^ x[12];
  assign t[298] = t[352] ^ x[11];
  assign t[299] = t[353] ^ x[15];
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[14];
  assign t[301] = t[355] ^ x[18];
  assign t[302] = t[356] ^ x[17];
  assign t[303] = t[357] ^ x[21];
  assign t[304] = t[358] ^ x[20];
  assign t[305] = t[359] ^ x[24];
  assign t[306] = t[360] ^ x[23];
  assign t[307] = t[361] ^ x[27];
  assign t[308] = t[362] ^ x[26];
  assign t[309] = t[363] ^ x[30];
  assign t[30] = ~(t[214]);
  assign t[310] = t[364] ^ x[29];
  assign t[311] = t[365] ^ x[33];
  assign t[312] = t[366] ^ x[32];
  assign t[313] = t[367] ^ x[36];
  assign t[314] = t[368] ^ x[35];
  assign t[315] = t[369] ^ x[39];
  assign t[316] = t[370] ^ x[38];
  assign t[317] = t[371] ^ x[42];
  assign t[318] = t[372] ^ x[41];
  assign t[319] = t[373] ^ x[45];
  assign t[31] = ~(t[215]);
  assign t[320] = t[374] ^ x[44];
  assign t[321] = t[375] ^ x[48];
  assign t[322] = t[376] ^ x[47];
  assign t[323] = t[377] ^ x[51];
  assign t[324] = t[378] ^ x[50];
  assign t[325] = t[379] ^ x[54];
  assign t[326] = t[380] ^ x[53];
  assign t[327] = t[381] ^ x[57];
  assign t[328] = t[382] ^ x[56];
  assign t[329] = t[383] ^ x[60];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[59];
  assign t[331] = t[385] ^ x[63];
  assign t[332] = t[386] ^ x[62];
  assign t[333] = t[387] ^ x[70];
  assign t[334] = t[388] ^ x[69];
  assign t[335] = t[389] ^ x[73];
  assign t[336] = t[390] ^ x[72];
  assign t[337] = t[391] ^ x[76];
  assign t[338] = t[392] ^ x[75];
  assign t[339] = t[393] ^ x[79];
  assign t[33] = t[51] ^ t[52];
  assign t[340] = t[394] ^ x[78];
  assign t[341] = t[395] ^ x[84];
  assign t[342] = t[396] ^ x[83];
  assign t[343] = t[397] ^ x[87];
  assign t[344] = t[398] ^ x[86];
  assign t[345] = t[399] ^ x[92];
  assign t[346] = t[400] ^ x[91];
  assign t[347] = (x[2]);
  assign t[348] = (x[2]);
  assign t[349] = (x[7]);
  assign t[34] = t[53] ^ t[54];
  assign t[350] = (x[7]);
  assign t[351] = (x[10]);
  assign t[352] = (x[10]);
  assign t[353] = (x[13]);
  assign t[354] = (x[13]);
  assign t[355] = (x[16]);
  assign t[356] = (x[16]);
  assign t[357] = (x[19]);
  assign t[358] = (x[19]);
  assign t[359] = (x[22]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[22]);
  assign t[361] = (x[25]);
  assign t[362] = (x[25]);
  assign t[363] = (x[28]);
  assign t[364] = (x[28]);
  assign t[365] = (x[31]);
  assign t[366] = (x[31]);
  assign t[367] = (x[34]);
  assign t[368] = (x[34]);
  assign t[369] = (x[37]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[37]);
  assign t[371] = (x[40]);
  assign t[372] = (x[40]);
  assign t[373] = (x[43]);
  assign t[374] = (x[43]);
  assign t[375] = (x[46]);
  assign t[376] = (x[46]);
  assign t[377] = (x[49]);
  assign t[378] = (x[49]);
  assign t[379] = (x[52]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[52]);
  assign t[381] = (x[55]);
  assign t[382] = (x[55]);
  assign t[383] = (x[58]);
  assign t[384] = (x[58]);
  assign t[385] = (x[61]);
  assign t[386] = (x[61]);
  assign t[387] = (x[68]);
  assign t[388] = (x[68]);
  assign t[389] = (x[71]);
  assign t[38] = ~(t[61] ^ t[62]);
  assign t[390] = (x[71]);
  assign t[391] = (x[74]);
  assign t[392] = (x[74]);
  assign t[393] = (x[77]);
  assign t[394] = (x[77]);
  assign t[395] = (x[82]);
  assign t[396] = (x[82]);
  assign t[397] = (x[85]);
  assign t[398] = (x[85]);
  assign t[399] = (x[90]);
  assign t[39] = ~(t[63] ^ t[64]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[90]);
  assign t[40] = t[65] ^ t[66];
  assign t[41] = t[67] ^ t[68];
  assign t[42] = t[69] ^ t[55];
  assign t[43] = ~(t[38] ^ t[70]);
  assign t[44] = t[11] ^ t[71];
  assign t[45] = ~(t[62] ^ t[41]);
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[216] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[217]);
  assign t[4] = t[8] ? t[9] : t[212];
  assign t[50] = ~(t[76] & t[218]);
  assign t[51] = t[77] ^ t[57];
  assign t[52] = t[78] & t[79];
  assign t[53] = t[80] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = t[84] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[218] ^ t[88];
  assign t[58] = t[89] ^ t[90];
  assign t[59] = t[27] ? t[91] : t[219];
  assign t[5] = ~(t[10]);
  assign t[60] = t[92] ^ t[93];
  assign t[61] = ~(t[94] ^ t[95]);
  assign t[62] = t[96] ^ t[97];
  assign t[63] = t[98] ^ t[99];
  assign t[64] = ~(t[70] ^ t[41]);
  assign t[65] = t[100] ^ t[67];
  assign t[66] = t[101] ^ t[102];
  assign t[67] = t[8] ? t[103] : t[220];
  assign t[68] = t[101] ^ t[87];
  assign t[69] = t[104] ^ t[105];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[106] ^ t[107];
  assign t[71] = t[108] ^ t[93];
  assign t[72] = ~(t[74] & t[109]);
  assign t[73] = ~(t[221] ^ t[110]);
  assign t[74] = ~(t[111] & t[112]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[222]);
  assign t[77] = t[113] ? t[114] : t[223];
  assign t[78] = ~(t[115]);
  assign t[79] = t[214] ^ t[116];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117];
  assign t[81] = ~t[118];
  assign t[82] = ~(t[53] ^ t[119]);
  assign t[83] = t[96] ^ t[120];
  assign t[84] = t[121] ^ t[59];
  assign t[85] = t[92] ^ t[122];
  assign t[86] = t[123] ^ t[100];
  assign t[87] = t[124] & t[125];
  assign t[88] = t[113] ? t[126] : t[224];
  assign t[89] = t[127] ^ t[52];
  assign t[8] = ~(t[15]);
  assign t[90] = t[128] & t[129];
  assign t[91] = t[219] ^ t[130];
  assign t[92] = t[131] ^ t[132];
  assign t[93] = t[133] & t[134];
  assign t[94] = t[40] ^ t[37];
  assign t[95] = t[135] ^ t[90];
  assign t[96] = t[81] ^ t[106];
  assign t[97] = t[119] ^ t[136];
  assign t[98] = t[137] ^ t[138];
  assign t[99] = t[139] ^ t[132];
  assign t[9] = t[212] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[141] ^ t[142];
  assign t[101] = t[217] ^ t[143];
  assign t[102] = t[218] ^ t[144];
  assign t[103] = t[27] ? t[145] : t[226];
  assign t[104] = ~(t[146] & t[147]);
  assign t[105] = t[148] ^ t[227];
  assign t[106] = ~(t[219]);
  assign t[107] = t[149] & t[148];
  assign t[108] = t[87] ^ t[127];
  assign t[109] = t[150] & t[151];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[216] ^ t[152];
  assign t[111] = t[112] ^ t[62];
  assign t[112] = t[153] ^ t[154];
  assign t[113] = t[155] & t[156];
  assign t[114] = t[221] ^ t[157];
  assign t[115] = t[158] ^ t[59];
  assign t[116] = t[127] ^ t[78];
  assign t[117] = t[115] ^ t[159];
  assign t[118] = t[160] ^ t[129];
  assign t[119] = t[161] & t[162];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[63] ^ t[163];
  assign t[121] = t[141] ^ t[98];
  assign t[122] = t[160] ^ t[124];
  assign t[123] = t[164] & t[165];
  assign t[124] = t[8] ? t[166] : t[228];
  assign t[125] = t[130] ^ t[119];
  assign t[126] = t[222] ^ t[167];
  assign t[127] = t[27] ? t[168] : t[229];
  assign t[128] = t[223] ^ t[169];
  assign t[129] = t[8] ? t[170] : t[230];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[171] ^ t[123];
  assign t[131] = t[172] & t[173];
  assign t[132] = ~(t[15]);
  assign t[133] = t[224] ^ t[174];
  assign t[134] = t[132] ? t[175] : t[231];
  assign t[135] = t[212] ^ t[176];
  assign t[136] = t[225] ^ t[177];
  assign t[137] = ~(t[142]);
  assign t[138] = ~(t[42]);
  assign t[139] = ~(t[43]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[40] ^ t[42];
  assign t[141] = t[42] ^ t[63];
  assign t[142] = t[68] ^ t[43];
  assign t[143] = t[178] ? x[71] : x[70];
  assign t[144] = t[178] ? x[73] : x[72];
  assign t[145] = t[226] ^ t[179];
  assign t[146] = ~(t[149] | t[148]);
  assign t[147] = ~(t[180] | t[106]);
  assign t[148] = ~(t[232]);
  assign t[149] = ~(t[227]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = ~(t[108] ^ t[115]);
  assign t[151] = t[116] ^ t[89];
  assign t[152] = t[132] ? t[181] : t[233];
  assign t[153] = t[182] & t[183];
  assign t[154] = t[184] & t[135];
  assign t[155] = ~(t[153] ^ t[185]);
  assign t[156] = t[186] ^ t[187];
  assign t[157] = t[72] ? x[81] : x[80];
  assign t[158] = t[188] & t[189];
  assign t[159] = t[190] & t[191];
  assign t[15] = ~(t[27]);
  assign t[160] = t[8] ? t[192] : t[234];
  assign t[161] = ~(t[118] ^ t[130]);
  assign t[162] = t[90] ^ t[165];
  assign t[163] = t[64] ^ t[26];
  assign t[164] = ~(t[129]);
  assign t[165] = t[8] ? t[193] : t[235];
  assign t[166] = t[228] ^ t[194];
  assign t[167] = t[28] ? x[89] : x[88];
  assign t[168] = t[229] ^ t[195];
  assign t[169] = t[72] ? x[91] : x[90];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[230] ^ t[196];
  assign t[171] = t[197] & t[198];
  assign t[172] = ~(t[171] ^ t[199]);
  assign t[173] = t[122] ^ t[200];
  assign t[174] = t[201] ? x[93] : x[92];
  assign t[175] = t[231] ^ t[202];
  assign t[176] = t[132] ? t[203] : t[236];
  assign t[177] = t[178] ? x[98] : x[97];
  assign t[178] = ~(t[48]);
  assign t[179] = t[178] ? x[100] : x[99];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[214]);
  assign t[181] = t[233] ^ t[204];
  assign t[182] = ~(t[187]);
  assign t[183] = ~(t[92]);
  assign t[184] = ~(t[93]);
  assign t[185] = t[76] ^ t[92];
  assign t[186] = t[92] ^ t[110];
  assign t[187] = t[135] ^ t[93];
  assign t[188] = ~(t[205]);
  assign t[189] = ~(t[87]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = ~(t[158] ^ t[206]);
  assign t[191] = t[58] ^ t[205];
  assign t[192] = t[234] ^ t[207];
  assign t[193] = t[235] ^ t[208];
  assign t[194] = t[178] ? x[102] : x[101];
  assign t[195] = t[28] ? x[104] : x[103];
  assign t[196] = t[178] ? x[106] : x[105];
  assign t[197] = ~(t[200]);
  assign t[198] = ~(t[160]);
  assign t[199] = t[90] ^ t[160];
  assign t[19] = ~(t[24] ^ t[33]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[165] ^ t[129];
  assign t[201] = ~(t[48]);
  assign t[202] = t[201] ? x[108] : x[107];
  assign t[203] = t[236] ^ t[209];
  assign t[204] = t[201] ? x[110] : x[109];
  assign t[205] = t[89] ^ t[127];
  assign t[206] = t[116] ^ t[87];
  assign t[207] = t[178] ? x[112] : x[111];
  assign t[208] = t[178] ? x[114] : x[113];
  assign t[209] = t[201] ? x[116] : x[115];
  assign t[20] = ~(t[34] ^ t[35]);
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[38] ^ t[14]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[9];
  assign t[239] = t[266] ^ x[12];
  assign t[23] = ~(t[38] ^ t[39]);
  assign t[240] = t[267] ^ x[15];
  assign t[241] = t[268] ^ x[18];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = t[40] ^ t[41];
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[51];
  assign t[253] = t[280] ^ x[54];
  assign t[254] = t[281] ^ x[57];
  assign t[255] = t[282] ^ x[60];
  assign t[256] = t[283] ^ x[63];
  assign t[257] = t[284] ^ x[66];
  assign t[258] = t[285] ^ x[69];
  assign t[259] = t[286] ^ x[76];
  assign t[25] = t[42] ^ t[43];
  assign t[260] = t[287] ^ x[79];
  assign t[261] = t[288] ^ x[84];
  assign t[262] = t[289] ^ x[87];
  assign t[263] = t[290] ^ x[96];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = t[44] & t[45];
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[9];
  assign t[294] = t[348] ^ x[8];
  assign t[295] = t[349] ^ x[12];
  assign t[296] = t[350] ^ x[11];
  assign t[297] = t[351] ^ x[15];
  assign t[298] = t[352] ^ x[14];
  assign t[299] = t[353] ^ x[18];
  assign t[29] = ~(t[211]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[17];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = ~(t[212]);
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[213]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[51];
  assign t[322] = t[376] ^ x[50];
  assign t[323] = t[377] ^ x[54];
  assign t[324] = t[378] ^ x[53];
  assign t[325] = t[379] ^ x[57];
  assign t[326] = t[380] ^ x[56];
  assign t[327] = t[381] ^ x[60];
  assign t[328] = t[382] ^ x[59];
  assign t[329] = t[383] ^ x[63];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[62];
  assign t[331] = t[385] ^ x[66];
  assign t[332] = t[386] ^ x[65];
  assign t[333] = t[387] ^ x[69];
  assign t[334] = t[388] ^ x[68];
  assign t[335] = t[389] ^ x[76];
  assign t[336] = t[390] ^ x[75];
  assign t[337] = t[391] ^ x[79];
  assign t[338] = t[392] ^ x[78];
  assign t[339] = t[393] ^ x[84];
  assign t[33] = ~(t[51] ^ t[52]);
  assign t[340] = t[394] ^ x[83];
  assign t[341] = t[395] ^ x[87];
  assign t[342] = t[396] ^ x[86];
  assign t[343] = t[397] ^ x[96];
  assign t[344] = t[398] ^ x[95];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[7]);
  assign t[348] = (x[7]);
  assign t[349] = (x[10]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[10]);
  assign t[351] = (x[13]);
  assign t[352] = (x[13]);
  assign t[353] = (x[16]);
  assign t[354] = (x[16]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = t[13] ^ t[55];
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[49]);
  assign t[376] = (x[49]);
  assign t[377] = (x[52]);
  assign t[378] = (x[52]);
  assign t[379] = (x[55]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[55]);
  assign t[381] = (x[58]);
  assign t[382] = (x[58]);
  assign t[383] = (x[61]);
  assign t[384] = (x[61]);
  assign t[385] = (x[64]);
  assign t[386] = (x[64]);
  assign t[387] = (x[67]);
  assign t[388] = (x[67]);
  assign t[389] = (x[74]);
  assign t[38] = t[60] ^ t[53];
  assign t[390] = (x[74]);
  assign t[391] = (x[77]);
  assign t[392] = (x[77]);
  assign t[393] = (x[82]);
  assign t[394] = (x[82]);
  assign t[395] = (x[85]);
  assign t[396] = (x[85]);
  assign t[397] = (x[94]);
  assign t[398] = (x[94]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[43] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66];
  assign t[43] = ~t[67];
  assign t[44] = ~(t[25] ^ t[64]);
  assign t[45] = t[40] ^ t[68];
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = t[214] | t[71];
  assign t[48] = ~(t[72]);
  assign t[49] = ~(t[215]);
  assign t[4] = t[8] ? t[9] : t[210];
  assign t[50] = ~(t[73] & t[216]);
  assign t[51] = ~(t[74] ^ t[75]);
  assign t[52] = t[76] ^ t[77];
  assign t[53] = t[78] ^ t[79];
  assign t[54] = t[80] ^ t[81];
  assign t[55] = ~(t[82] ^ t[83]);
  assign t[56] = t[84] ^ t[33];
  assign t[57] = ~(t[85] ^ t[86]);
  assign t[58] = t[87] ^ t[78];
  assign t[59] = t[88] & t[89];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92] ^ t[93];
  assign t[62] = t[94] & t[95];
  assign t[63] = ~t[96];
  assign t[64] = t[97] ^ t[98];
  assign t[65] = t[99] & t[100];
  assign t[66] = t[8] ? t[101] : t[217];
  assign t[67] = t[8] ? t[102] : t[218];
  assign t[68] = t[103];
  assign t[69] = ~(t[71] & t[104]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[219] ^ t[105]);
  assign t[71] = ~(t[106] & t[107]);
  assign t[72] = ~(t[47]);
  assign t[73] = ~(t[220]);
  assign t[74] = t[108] ^ t[109];
  assign t[75] = t[110] ^ t[111];
  assign t[76] = t[93] ^ t[110];
  assign t[77] = t[112] ^ t[113];
  assign t[78] = t[27] ? t[114] : t[221];
  assign t[79] = t[115] ^ t[109];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[116] ^ t[117];
  assign t[81] = t[118] ^ t[119];
  assign t[82] = t[52] ^ t[37];
  assign t[83] = ~(t[120] ^ t[86]);
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[122] ^ t[123];
  assign t[86] = t[124] ^ t[125];
  assign t[87] = t[27] ? t[126] : t[222];
  assign t[88] = ~(t[127]);
  assign t[89] = t[27] ? t[128] : t[223];
  assign t[8] = ~(t[15]);
  assign t[90] = t[129] ^ t[124];
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[132] ? t[133] : t[224];
  assign t[93] = t[211] ^ t[134];
  assign t[94] = ~(t[61] ^ t[112]);
  assign t[95] = t[76] ^ t[135];
  assign t[96] = t[8] ? t[136] : t[225];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[139] & t[68];
  assign t[99] = ~(t[97] ^ t[140]);
  assign t[9] = t[210] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[141] ^ t[142];
  assign t[101] = t[217] ^ t[143];
  assign t[102] = t[218] ^ t[144];
  assign t[103] = t[27] ? t[145] : t[226];
  assign t[104] = ~(t[146] & t[147]);
  assign t[105] = t[148] ^ t[227];
  assign t[106] = ~(t[219]);
  assign t[107] = t[149] & t[148];
  assign t[108] = t[87] ^ t[127];
  assign t[109] = t[150] & t[151];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[216] ^ t[152];
  assign t[111] = t[112] ^ t[62];
  assign t[112] = t[153] ^ t[154];
  assign t[113] = t[155] & t[156];
  assign t[114] = t[221] ^ t[157];
  assign t[115] = t[158] ^ t[59];
  assign t[116] = t[127] ^ t[78];
  assign t[117] = t[115] ^ t[159];
  assign t[118] = t[160] ^ t[129];
  assign t[119] = t[161] & t[162];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[63] ^ t[163];
  assign t[121] = t[141] ^ t[98];
  assign t[122] = t[160] ^ t[124];
  assign t[123] = t[164] & t[165];
  assign t[124] = t[8] ? t[166] : t[228];
  assign t[125] = t[130] ^ t[119];
  assign t[126] = t[222] ^ t[167];
  assign t[127] = t[27] ? t[168] : t[229];
  assign t[128] = t[223] ^ t[169];
  assign t[129] = t[8] ? t[170] : t[230];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[171] ^ t[123];
  assign t[131] = t[172] & t[173];
  assign t[132] = ~(t[15]);
  assign t[133] = t[224] ^ t[174];
  assign t[134] = t[132] ? t[175] : t[231];
  assign t[135] = t[212] ^ t[176];
  assign t[136] = t[225] ^ t[177];
  assign t[137] = ~(t[142]);
  assign t[138] = ~(t[42]);
  assign t[139] = ~(t[43]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[40] ^ t[42];
  assign t[141] = t[42] ^ t[63];
  assign t[142] = t[68] ^ t[43];
  assign t[143] = t[178] ? x[71] : x[70];
  assign t[144] = t[178] ? x[73] : x[72];
  assign t[145] = t[226] ^ t[179];
  assign t[146] = ~(t[149] | t[148]);
  assign t[147] = ~(t[180] | t[106]);
  assign t[148] = ~(t[232]);
  assign t[149] = ~(t[227]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = ~(t[108] ^ t[115]);
  assign t[151] = t[116] ^ t[89];
  assign t[152] = t[132] ? t[181] : t[233];
  assign t[153] = t[182] & t[183];
  assign t[154] = t[184] & t[135];
  assign t[155] = ~(t[153] ^ t[185]);
  assign t[156] = t[186] ^ t[187];
  assign t[157] = t[72] ? x[81] : x[80];
  assign t[158] = t[188] & t[189];
  assign t[159] = t[190] & t[191];
  assign t[15] = ~(t[27]);
  assign t[160] = t[8] ? t[192] : t[234];
  assign t[161] = ~(t[118] ^ t[130]);
  assign t[162] = t[90] ^ t[165];
  assign t[163] = t[64] ^ t[26];
  assign t[164] = ~(t[129]);
  assign t[165] = t[8] ? t[193] : t[235];
  assign t[166] = t[228] ^ t[194];
  assign t[167] = t[28] ? x[89] : x[88];
  assign t[168] = t[229] ^ t[195];
  assign t[169] = t[72] ? x[91] : x[90];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[230] ^ t[196];
  assign t[171] = t[197] & t[198];
  assign t[172] = ~(t[171] ^ t[199]);
  assign t[173] = t[122] ^ t[200];
  assign t[174] = t[201] ? x[93] : x[92];
  assign t[175] = t[231] ^ t[202];
  assign t[176] = t[132] ? t[203] : t[236];
  assign t[177] = t[178] ? x[98] : x[97];
  assign t[178] = ~(t[48]);
  assign t[179] = t[178] ? x[100] : x[99];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[214]);
  assign t[181] = t[233] ^ t[204];
  assign t[182] = ~(t[187]);
  assign t[183] = ~(t[92]);
  assign t[184] = ~(t[93]);
  assign t[185] = t[76] ^ t[92];
  assign t[186] = t[92] ^ t[110];
  assign t[187] = t[135] ^ t[93];
  assign t[188] = ~(t[205]);
  assign t[189] = ~(t[87]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = ~(t[158] ^ t[206]);
  assign t[191] = t[58] ^ t[205];
  assign t[192] = t[234] ^ t[207];
  assign t[193] = t[235] ^ t[208];
  assign t[194] = t[178] ? x[102] : x[101];
  assign t[195] = t[28] ? x[104] : x[103];
  assign t[196] = t[178] ? x[106] : x[105];
  assign t[197] = ~(t[200]);
  assign t[198] = ~(t[160]);
  assign t[199] = t[90] ^ t[160];
  assign t[19] = ~(t[24] ^ t[33]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[165] ^ t[129];
  assign t[201] = ~(t[48]);
  assign t[202] = t[201] ? x[108] : x[107];
  assign t[203] = t[236] ^ t[209];
  assign t[204] = t[201] ? x[110] : x[109];
  assign t[205] = t[89] ^ t[127];
  assign t[206] = t[116] ^ t[87];
  assign t[207] = t[178] ? x[112] : x[111];
  assign t[208] = t[178] ? x[114] : x[113];
  assign t[209] = t[201] ? x[116] : x[115];
  assign t[20] = ~(t[34] ^ t[35]);
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[38] ^ t[14]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[9];
  assign t[239] = t[266] ^ x[12];
  assign t[23] = ~(t[38] ^ t[39]);
  assign t[240] = t[267] ^ x[15];
  assign t[241] = t[268] ^ x[18];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = t[40] ^ t[41];
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[51];
  assign t[253] = t[280] ^ x[54];
  assign t[254] = t[281] ^ x[57];
  assign t[255] = t[282] ^ x[60];
  assign t[256] = t[283] ^ x[63];
  assign t[257] = t[284] ^ x[66];
  assign t[258] = t[285] ^ x[69];
  assign t[259] = t[286] ^ x[76];
  assign t[25] = t[42] ^ t[43];
  assign t[260] = t[287] ^ x[79];
  assign t[261] = t[288] ^ x[84];
  assign t[262] = t[289] ^ x[87];
  assign t[263] = t[290] ^ x[96];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = t[44] & t[45];
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[9];
  assign t[294] = t[348] ^ x[8];
  assign t[295] = t[349] ^ x[12];
  assign t[296] = t[350] ^ x[11];
  assign t[297] = t[351] ^ x[15];
  assign t[298] = t[352] ^ x[14];
  assign t[299] = t[353] ^ x[18];
  assign t[29] = ~(t[211]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[17];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = ~(t[212]);
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[213]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[51];
  assign t[322] = t[376] ^ x[50];
  assign t[323] = t[377] ^ x[54];
  assign t[324] = t[378] ^ x[53];
  assign t[325] = t[379] ^ x[57];
  assign t[326] = t[380] ^ x[56];
  assign t[327] = t[381] ^ x[60];
  assign t[328] = t[382] ^ x[59];
  assign t[329] = t[383] ^ x[63];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[62];
  assign t[331] = t[385] ^ x[66];
  assign t[332] = t[386] ^ x[65];
  assign t[333] = t[387] ^ x[69];
  assign t[334] = t[388] ^ x[68];
  assign t[335] = t[389] ^ x[76];
  assign t[336] = t[390] ^ x[75];
  assign t[337] = t[391] ^ x[79];
  assign t[338] = t[392] ^ x[78];
  assign t[339] = t[393] ^ x[84];
  assign t[33] = ~(t[51] ^ t[52]);
  assign t[340] = t[394] ^ x[83];
  assign t[341] = t[395] ^ x[87];
  assign t[342] = t[396] ^ x[86];
  assign t[343] = t[397] ^ x[96];
  assign t[344] = t[398] ^ x[95];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[7]);
  assign t[348] = (x[7]);
  assign t[349] = (x[10]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[10]);
  assign t[351] = (x[13]);
  assign t[352] = (x[13]);
  assign t[353] = (x[16]);
  assign t[354] = (x[16]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = t[13] ^ t[55];
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[49]);
  assign t[376] = (x[49]);
  assign t[377] = (x[52]);
  assign t[378] = (x[52]);
  assign t[379] = (x[55]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[55]);
  assign t[381] = (x[58]);
  assign t[382] = (x[58]);
  assign t[383] = (x[61]);
  assign t[384] = (x[61]);
  assign t[385] = (x[64]);
  assign t[386] = (x[64]);
  assign t[387] = (x[67]);
  assign t[388] = (x[67]);
  assign t[389] = (x[74]);
  assign t[38] = t[60] ^ t[53];
  assign t[390] = (x[74]);
  assign t[391] = (x[77]);
  assign t[392] = (x[77]);
  assign t[393] = (x[82]);
  assign t[394] = (x[82]);
  assign t[395] = (x[85]);
  assign t[396] = (x[85]);
  assign t[397] = (x[94]);
  assign t[398] = (x[94]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[43] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[66];
  assign t[43] = ~t[67];
  assign t[44] = ~(t[25] ^ t[64]);
  assign t[45] = t[40] ^ t[68];
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = t[214] | t[71];
  assign t[48] = ~(t[72]);
  assign t[49] = ~(t[215]);
  assign t[4] = t[8] ? t[9] : t[210];
  assign t[50] = ~(t[73] & t[216]);
  assign t[51] = ~(t[74] ^ t[75]);
  assign t[52] = t[76] ^ t[77];
  assign t[53] = t[78] ^ t[79];
  assign t[54] = t[80] ^ t[81];
  assign t[55] = ~(t[82] ^ t[83]);
  assign t[56] = t[84] ^ t[33];
  assign t[57] = ~(t[85] ^ t[86]);
  assign t[58] = t[87] ^ t[78];
  assign t[59] = t[88] & t[89];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92] ^ t[93];
  assign t[62] = t[94] & t[95];
  assign t[63] = ~t[96];
  assign t[64] = t[97] ^ t[98];
  assign t[65] = t[99] & t[100];
  assign t[66] = t[8] ? t[101] : t[217];
  assign t[67] = t[8] ? t[102] : t[218];
  assign t[68] = t[103];
  assign t[69] = ~(t[71] & t[104]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[219] ^ t[105]);
  assign t[71] = ~(t[106] & t[107]);
  assign t[72] = ~(t[47]);
  assign t[73] = ~(t[220]);
  assign t[74] = t[108] ^ t[109];
  assign t[75] = t[110] ^ t[111];
  assign t[76] = t[93] ^ t[110];
  assign t[77] = t[112] ^ t[113];
  assign t[78] = t[27] ? t[114] : t[221];
  assign t[79] = t[115] ^ t[109];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[116] ^ t[117];
  assign t[81] = t[118] ^ t[119];
  assign t[82] = t[52] ^ t[37];
  assign t[83] = ~(t[120] ^ t[86]);
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[122] ^ t[123];
  assign t[86] = t[124] ^ t[125];
  assign t[87] = t[27] ? t[126] : t[222];
  assign t[88] = ~(t[127]);
  assign t[89] = t[27] ? t[128] : t[223];
  assign t[8] = ~(t[15]);
  assign t[90] = t[129] ^ t[124];
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[132] ? t[133] : t[224];
  assign t[93] = t[211] ^ t[134];
  assign t[94] = ~(t[61] ^ t[112]);
  assign t[95] = t[76] ^ t[135];
  assign t[96] = t[8] ? t[136] : t[225];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[139] & t[68];
  assign t[99] = ~(t[97] ^ t[140]);
  assign t[9] = t[210] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind136(x, y);
 input [116:0] x;
 output y;

 wire [400:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[116] ^ t[142];
  assign t[101] = t[221] ^ t[143];
  assign t[102] = t[222] ^ t[144];
  assign t[103] = t[223] ^ t[145];
  assign t[104] = t[224] ^ t[146];
  assign t[105] = ~(t[117] ^ t[57]);
  assign t[106] = t[35] ^ t[127];
  assign t[107] = t[225] ^ t[147];
  assign t[108] = t[148] & t[149];
  assign t[109] = t[150] & t[151];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[93] ^ t[72]);
  assign t[111] = t[152] ^ t[151];
  assign t[112] = ~(t[153] & t[154]);
  assign t[113] = t[155] ^ t[230];
  assign t[114] = ~(t[226]);
  assign t[115] = t[156] & t[155];
  assign t[116] = t[157] ^ t[62];
  assign t[117] = t[158] ^ t[56];
  assign t[118] = t[122] ^ t[159];
  assign t[119] = t[63] ^ t[160];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[228] ^ t[161];
  assign t[121] = t[162] ^ t[42];
  assign t[122] = t[83] ^ t[66];
  assign t[123] = t[229] ^ t[163];
  assign t[124] = ~(t[130]);
  assign t[125] = ~(t[158]);
  assign t[126] = ~(t[56]);
  assign t[127] = t[227] ^ t[164];
  assign t[128] = t[35] ^ t[158];
  assign t[129] = t[158] ^ t[43];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[127] ^ t[56];
  assign t[131] = ~(t[165] ^ t[166]);
  assign t[132] = t[167] ^ t[168];
  assign t[133] = t[169];
  assign t[134] = ~t[170];
  assign t[135] = t[171] ? x[62] : x[61];
  assign t[136] = t[171] ? x[64] : x[63];
  assign t[137] = ~(t[142]);
  assign t[138] = ~(t[157]);
  assign t[139] = ~(t[61]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[94] ? t[172] : t[231];
  assign t[141] = t[39] ^ t[157];
  assign t[142] = t[140] ^ t[61];
  assign t[143] = t[173] ? x[69] : x[68];
  assign t[144] = t[77] ? x[71] : x[70];
  assign t[145] = t[173] ? x[73] : x[72];
  assign t[146] = t[28] ? x[75] : x[74];
  assign t[147] = t[77] ? x[77] : x[76];
  assign t[148] = ~(t[174]);
  assign t[149] = ~(t[133]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[134]);
  assign t[151] = t[175];
  assign t[152] = t[134] ^ t[45];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[176] | t[114]);
  assign t[155] = ~(t[232]);
  assign t[156] = ~(t[230]);
  assign t[157] = t[94] ? t[177] : t[233];
  assign t[158] = t[8] ? t[178] : t[234];
  assign t[159] = t[121] ^ t[179];
  assign t[15] = ~(t[27]);
  assign t[160] = t[180] & t[181];
  assign t[161] = t[173] ? x[88] : x[87];
  assign t[162] = t[182] & t[183];
  assign t[163] = t[28] ? x[90] : x[89];
  assign t[164] = t[8] ? t[184] : t[235];
  assign t[165] = t[185] ^ t[186];
  assign t[166] = ~(t[187] ^ t[26]);
  assign t[167] = t[152] ^ t[188];
  assign t[168] = t[66] ^ t[189];
  assign t[169] = t[8] ? t[190] : t[236];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[8] ? t[191] : t[237];
  assign t[171] = ~(t[49]);
  assign t[172] = t[231] ^ t[192];
  assign t[173] = ~(t[49]);
  assign t[174] = t[151] ^ t[134];
  assign t[175] = t[8] ? t[193] : t[238];
  assign t[176] = ~(t[217]);
  assign t[177] = t[233] ^ t[194];
  assign t[178] = t[234] ^ t[195];
  assign t[179] = t[196] & t[197];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[198] ^ t[63]);
  assign t[181] = t[39] ^ t[140];
  assign t[182] = ~(t[199]);
  assign t[183] = ~(t[65]);
  assign t[184] = t[235] ^ t[200];
  assign t[185] = t[25] ^ t[201];
  assign t[186] = ~(t[202] ^ t[23]);
  assign t[187] = t[203] ^ t[109];
  assign t[188] = t[72] ^ t[204];
  assign t[189] = t[121] ^ t[55];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[236] ^ t[205];
  assign t[191] = t[237] ^ t[206];
  assign t[192] = t[171] ? x[104] : x[103];
  assign t[193] = t[238] ^ t[207];
  assign t[194] = t[171] ? x[106] : x[105];
  assign t[195] = t[28] ? x[108] : x[107];
  assign t[196] = ~(t[162] ^ t[208]);
  assign t[197] = t[41] ^ t[199];
  assign t[198] = t[157] ^ t[61];
  assign t[199] = t[68] ^ t[83];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[28] ? x[110] : x[109];
  assign t[201] = t[129] ^ t[88];
  assign t[202] = ~(t[34] ^ t[82]);
  assign t[203] = t[133] ^ t[45];
  assign t[204] = t[209] & t[210];
  assign t[205] = t[77] ? x[112] : x[111];
  assign t[206] = t[28] ? x[114] : x[113];
  assign t[207] = t[77] ? x[116] : x[115];
  assign t[208] = t[122] ^ t[65];
  assign t[209] = ~(t[108] ^ t[211]);
  assign t[20] = ~(t[21] ^ t[26]);
  assign t[210] = t[203] ^ t[174];
  assign t[211] = t[152] ^ t[133];
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[35] ^ t[36];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[37] ^ t[38]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = t[266] ^ x[4];
  assign t[23] = t[39] ^ t[40];
  assign t[240] = t[267] ^ x[9];
  assign t[241] = t[268] ^ x[12];
  assign t[242] = t[269] ^ x[15];
  assign t[243] = t[270] ^ x[18];
  assign t[244] = t[271] ^ x[21];
  assign t[245] = t[272] ^ x[24];
  assign t[246] = t[273] ^ x[27];
  assign t[247] = t[274] ^ x[30];
  assign t[248] = t[275] ^ x[33];
  assign t[249] = t[276] ^ x[36];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[277] ^ x[39];
  assign t[251] = t[278] ^ x[42];
  assign t[252] = t[279] ^ x[45];
  assign t[253] = t[280] ^ x[48];
  assign t[254] = t[281] ^ x[51];
  assign t[255] = t[282] ^ x[54];
  assign t[256] = t[283] ^ x[57];
  assign t[257] = t[284] ^ x[60];
  assign t[258] = t[285] ^ x[67];
  assign t[259] = t[286] ^ x[80];
  assign t[25] = t[43] ^ t[44];
  assign t[260] = t[287] ^ x[83];
  assign t[261] = t[288] ^ x[86];
  assign t[262] = t[289] ^ x[93];
  assign t[263] = t[290] ^ x[96];
  assign t[264] = t[291] ^ x[99];
  assign t[265] = t[292] ^ x[102];
  assign t[266] = (t[293] & ~t[294]);
  assign t[267] = (t[295] & ~t[296]);
  assign t[268] = (t[297] & ~t[298]);
  assign t[269] = (t[299] & ~t[300]);
  assign t[26] = t[45] ^ t[46];
  assign t[270] = (t[301] & ~t[302]);
  assign t[271] = (t[303] & ~t[304]);
  assign t[272] = (t[305] & ~t[306]);
  assign t[273] = (t[307] & ~t[308]);
  assign t[274] = (t[309] & ~t[310]);
  assign t[275] = (t[311] & ~t[312]);
  assign t[276] = (t[313] & ~t[314]);
  assign t[277] = (t[315] & ~t[316]);
  assign t[278] = (t[317] & ~t[318]);
  assign t[279] = (t[319] & ~t[320]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = ~(t[49]);
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = t[347] ^ x[4];
  assign t[294] = t[348] ^ x[3];
  assign t[295] = t[349] ^ x[9];
  assign t[296] = t[350] ^ x[8];
  assign t[297] = t[351] ^ x[12];
  assign t[298] = t[352] ^ x[11];
  assign t[299] = t[353] ^ x[15];
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[14];
  assign t[301] = t[355] ^ x[18];
  assign t[302] = t[356] ^ x[17];
  assign t[303] = t[357] ^ x[21];
  assign t[304] = t[358] ^ x[20];
  assign t[305] = t[359] ^ x[24];
  assign t[306] = t[360] ^ x[23];
  assign t[307] = t[361] ^ x[27];
  assign t[308] = t[362] ^ x[26];
  assign t[309] = t[363] ^ x[30];
  assign t[30] = ~(t[214]);
  assign t[310] = t[364] ^ x[29];
  assign t[311] = t[365] ^ x[33];
  assign t[312] = t[366] ^ x[32];
  assign t[313] = t[367] ^ x[36];
  assign t[314] = t[368] ^ x[35];
  assign t[315] = t[369] ^ x[39];
  assign t[316] = t[370] ^ x[38];
  assign t[317] = t[371] ^ x[42];
  assign t[318] = t[372] ^ x[41];
  assign t[319] = t[373] ^ x[45];
  assign t[31] = ~(t[215]);
  assign t[320] = t[374] ^ x[44];
  assign t[321] = t[375] ^ x[48];
  assign t[322] = t[376] ^ x[47];
  assign t[323] = t[377] ^ x[51];
  assign t[324] = t[378] ^ x[50];
  assign t[325] = t[379] ^ x[54];
  assign t[326] = t[380] ^ x[53];
  assign t[327] = t[381] ^ x[57];
  assign t[328] = t[382] ^ x[56];
  assign t[329] = t[383] ^ x[60];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[59];
  assign t[331] = t[385] ^ x[67];
  assign t[332] = t[386] ^ x[66];
  assign t[333] = t[387] ^ x[80];
  assign t[334] = t[388] ^ x[79];
  assign t[335] = t[389] ^ x[83];
  assign t[336] = t[390] ^ x[82];
  assign t[337] = t[391] ^ x[86];
  assign t[338] = t[392] ^ x[85];
  assign t[339] = t[393] ^ x[93];
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[340] = t[394] ^ x[92];
  assign t[341] = t[395] ^ x[96];
  assign t[342] = t[396] ^ x[95];
  assign t[343] = t[397] ^ x[99];
  assign t[344] = t[398] ^ x[98];
  assign t[345] = t[399] ^ x[102];
  assign t[346] = t[400] ^ x[101];
  assign t[347] = (x[2]);
  assign t[348] = (x[2]);
  assign t[349] = (x[7]);
  assign t[34] = t[54] ^ t[55];
  assign t[350] = (x[7]);
  assign t[351] = (x[10]);
  assign t[352] = (x[10]);
  assign t[353] = (x[13]);
  assign t[354] = (x[13]);
  assign t[355] = (x[16]);
  assign t[356] = (x[16]);
  assign t[357] = (x[19]);
  assign t[358] = (x[19]);
  assign t[359] = (x[22]);
  assign t[35] = t[56] ^ t[43];
  assign t[360] = (x[22]);
  assign t[361] = (x[25]);
  assign t[362] = (x[25]);
  assign t[363] = (x[28]);
  assign t[364] = (x[28]);
  assign t[365] = (x[31]);
  assign t[366] = (x[31]);
  assign t[367] = (x[34]);
  assign t[368] = (x[34]);
  assign t[369] = (x[37]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[37]);
  assign t[371] = (x[40]);
  assign t[372] = (x[40]);
  assign t[373] = (x[43]);
  assign t[374] = (x[43]);
  assign t[375] = (x[46]);
  assign t[376] = (x[46]);
  assign t[377] = (x[49]);
  assign t[378] = (x[49]);
  assign t[379] = (x[52]);
  assign t[37] = t[59] ^ t[33];
  assign t[380] = (x[52]);
  assign t[381] = (x[55]);
  assign t[382] = (x[55]);
  assign t[383] = (x[58]);
  assign t[384] = (x[58]);
  assign t[385] = (x[65]);
  assign t[386] = (x[65]);
  assign t[387] = (x[78]);
  assign t[388] = (x[78]);
  assign t[389] = (x[81]);
  assign t[38] = ~(t[25] ^ t[60]);
  assign t[390] = (x[81]);
  assign t[391] = (x[84]);
  assign t[392] = (x[84]);
  assign t[393] = (x[91]);
  assign t[394] = (x[91]);
  assign t[395] = (x[94]);
  assign t[396] = (x[94]);
  assign t[397] = (x[97]);
  assign t[398] = (x[97]);
  assign t[399] = (x[100]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[100]);
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] & t[68];
  assign t[43] = t[216] ^ t[69];
  assign t[44] = t[57] ^ t[70];
  assign t[45] = t[71];
  assign t[46] = t[72] ^ t[73];
  assign t[47] = ~(t[74] & t[75]);
  assign t[48] = t[217] | t[76];
  assign t[49] = ~(t[77]);
  assign t[4] = t[8] ? t[9] : t[212];
  assign t[50] = ~(t[216]);
  assign t[51] = ~(t[78] & t[218]);
  assign t[52] = t[79] ^ t[80];
  assign t[53] = ~(t[81] ^ t[82]);
  assign t[54] = t[65] ^ t[83];
  assign t[55] = t[84] & t[85];
  assign t[56] = t[215] ^ t[86];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] & t[90];
  assign t[59] = ~(t[91] ^ t[92]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] ^ t[73];
  assign t[61] = t[94] ? t[95] : t[219];
  assign t[62] = t[94] ? t[96] : t[220];
  assign t[63] = t[97] ^ t[98];
  assign t[64] = t[99] & t[100];
  assign t[65] = t[8] ? t[101] : t[221];
  assign t[66] = t[8] ? t[102] : t[222];
  assign t[67] = ~(t[83]);
  assign t[68] = t[8] ? t[103] : t[223];
  assign t[69] = t[8] ? t[104] : t[224];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[105] & t[106];
  assign t[71] = t[8] ? t[107] : t[225];
  assign t[72] = t[108] ^ t[109];
  assign t[73] = t[110] & t[111];
  assign t[74] = ~(t[76] & t[112]);
  assign t[75] = ~(t[226] ^ t[113]);
  assign t[76] = ~(t[114] & t[115]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[227]);
  assign t[79] = t[116] ^ t[98];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] ^ t[70];
  assign t[81] = t[118] ^ t[60];
  assign t[82] = t[62] ^ t[119];
  assign t[83] = t[8] ? t[120] : t[228];
  assign t[84] = ~(t[54] ^ t[121]);
  assign t[85] = t[122] ^ t[68];
  assign t[86] = t[8] ? t[123] : t[229];
  assign t[87] = t[124] & t[125];
  assign t[88] = t[126] & t[127];
  assign t[89] = ~(t[87] ^ t[128]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[131] ^ t[24];
  assign t[92] = ~(t[132] ^ t[80]);
  assign t[93] = t[133] ^ t[134];
  assign t[94] = ~(t[15]);
  assign t[95] = t[219] ^ t[135];
  assign t[96] = t[220] ^ t[136];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[139] & t[140];
  assign t[99] = ~(t[97] ^ t[141]);
  assign t[9] = t[212] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [116:0] x;
 output y;

 wire [400:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[116] ^ t[142];
  assign t[101] = t[221] ^ t[143];
  assign t[102] = t[222] ^ t[144];
  assign t[103] = t[223] ^ t[145];
  assign t[104] = t[224] ^ t[146];
  assign t[105] = ~(t[117] ^ t[57]);
  assign t[106] = t[35] ^ t[127];
  assign t[107] = t[225] ^ t[147];
  assign t[108] = t[148] & t[149];
  assign t[109] = t[150] & t[151];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[93] ^ t[72]);
  assign t[111] = t[152] ^ t[151];
  assign t[112] = ~(t[153] & t[154]);
  assign t[113] = t[155] ^ t[230];
  assign t[114] = ~(t[226]);
  assign t[115] = t[156] & t[155];
  assign t[116] = t[157] ^ t[62];
  assign t[117] = t[158] ^ t[56];
  assign t[118] = t[122] ^ t[159];
  assign t[119] = t[63] ^ t[160];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[228] ^ t[161];
  assign t[121] = t[162] ^ t[42];
  assign t[122] = t[83] ^ t[66];
  assign t[123] = t[229] ^ t[163];
  assign t[124] = ~(t[130]);
  assign t[125] = ~(t[158]);
  assign t[126] = ~(t[56]);
  assign t[127] = t[227] ^ t[164];
  assign t[128] = t[35] ^ t[158];
  assign t[129] = t[158] ^ t[43];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[127] ^ t[56];
  assign t[131] = ~(t[165] ^ t[166]);
  assign t[132] = t[167] ^ t[168];
  assign t[133] = t[169];
  assign t[134] = ~t[170];
  assign t[135] = t[171] ? x[62] : x[61];
  assign t[136] = t[171] ? x[64] : x[63];
  assign t[137] = ~(t[142]);
  assign t[138] = ~(t[157]);
  assign t[139] = ~(t[61]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[94] ? t[172] : t[231];
  assign t[141] = t[39] ^ t[157];
  assign t[142] = t[140] ^ t[61];
  assign t[143] = t[173] ? x[69] : x[68];
  assign t[144] = t[77] ? x[71] : x[70];
  assign t[145] = t[173] ? x[73] : x[72];
  assign t[146] = t[28] ? x[75] : x[74];
  assign t[147] = t[77] ? x[77] : x[76];
  assign t[148] = ~(t[174]);
  assign t[149] = ~(t[133]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[134]);
  assign t[151] = t[175];
  assign t[152] = t[134] ^ t[45];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[176] | t[114]);
  assign t[155] = ~(t[232]);
  assign t[156] = ~(t[230]);
  assign t[157] = t[94] ? t[177] : t[233];
  assign t[158] = t[8] ? t[178] : t[234];
  assign t[159] = t[121] ^ t[179];
  assign t[15] = ~(t[27]);
  assign t[160] = t[180] & t[181];
  assign t[161] = t[173] ? x[88] : x[87];
  assign t[162] = t[182] & t[183];
  assign t[163] = t[28] ? x[90] : x[89];
  assign t[164] = t[8] ? t[184] : t[235];
  assign t[165] = t[185] ^ t[186];
  assign t[166] = ~(t[187] ^ t[26]);
  assign t[167] = t[152] ^ t[188];
  assign t[168] = t[66] ^ t[189];
  assign t[169] = t[8] ? t[190] : t[236];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[8] ? t[191] : t[237];
  assign t[171] = ~(t[49]);
  assign t[172] = t[231] ^ t[192];
  assign t[173] = ~(t[49]);
  assign t[174] = t[151] ^ t[134];
  assign t[175] = t[8] ? t[193] : t[238];
  assign t[176] = ~(t[217]);
  assign t[177] = t[233] ^ t[194];
  assign t[178] = t[234] ^ t[195];
  assign t[179] = t[196] & t[197];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[198] ^ t[63]);
  assign t[181] = t[39] ^ t[140];
  assign t[182] = ~(t[199]);
  assign t[183] = ~(t[65]);
  assign t[184] = t[235] ^ t[200];
  assign t[185] = t[25] ^ t[201];
  assign t[186] = ~(t[202] ^ t[23]);
  assign t[187] = t[203] ^ t[109];
  assign t[188] = t[72] ^ t[204];
  assign t[189] = t[121] ^ t[55];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[236] ^ t[205];
  assign t[191] = t[237] ^ t[206];
  assign t[192] = t[171] ? x[104] : x[103];
  assign t[193] = t[238] ^ t[207];
  assign t[194] = t[171] ? x[106] : x[105];
  assign t[195] = t[28] ? x[108] : x[107];
  assign t[196] = ~(t[162] ^ t[208]);
  assign t[197] = t[41] ^ t[199];
  assign t[198] = t[157] ^ t[61];
  assign t[199] = t[68] ^ t[83];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[28] ? x[110] : x[109];
  assign t[201] = t[129] ^ t[88];
  assign t[202] = ~(t[34] ^ t[82]);
  assign t[203] = t[133] ^ t[45];
  assign t[204] = t[209] & t[210];
  assign t[205] = t[77] ? x[112] : x[111];
  assign t[206] = t[28] ? x[114] : x[113];
  assign t[207] = t[77] ? x[116] : x[115];
  assign t[208] = t[122] ^ t[65];
  assign t[209] = ~(t[108] ^ t[211]);
  assign t[20] = ~(t[21] ^ t[26]);
  assign t[210] = t[203] ^ t[174];
  assign t[211] = t[152] ^ t[133];
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[35] ^ t[36];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[37] ^ t[38]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = t[266] ^ x[4];
  assign t[23] = t[39] ^ t[40];
  assign t[240] = t[267] ^ x[9];
  assign t[241] = t[268] ^ x[12];
  assign t[242] = t[269] ^ x[15];
  assign t[243] = t[270] ^ x[18];
  assign t[244] = t[271] ^ x[21];
  assign t[245] = t[272] ^ x[24];
  assign t[246] = t[273] ^ x[27];
  assign t[247] = t[274] ^ x[30];
  assign t[248] = t[275] ^ x[33];
  assign t[249] = t[276] ^ x[36];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[277] ^ x[39];
  assign t[251] = t[278] ^ x[42];
  assign t[252] = t[279] ^ x[45];
  assign t[253] = t[280] ^ x[48];
  assign t[254] = t[281] ^ x[51];
  assign t[255] = t[282] ^ x[54];
  assign t[256] = t[283] ^ x[57];
  assign t[257] = t[284] ^ x[60];
  assign t[258] = t[285] ^ x[67];
  assign t[259] = t[286] ^ x[80];
  assign t[25] = t[43] ^ t[44];
  assign t[260] = t[287] ^ x[83];
  assign t[261] = t[288] ^ x[86];
  assign t[262] = t[289] ^ x[93];
  assign t[263] = t[290] ^ x[96];
  assign t[264] = t[291] ^ x[99];
  assign t[265] = t[292] ^ x[102];
  assign t[266] = (t[293] & ~t[294]);
  assign t[267] = (t[295] & ~t[296]);
  assign t[268] = (t[297] & ~t[298]);
  assign t[269] = (t[299] & ~t[300]);
  assign t[26] = t[45] ^ t[46];
  assign t[270] = (t[301] & ~t[302]);
  assign t[271] = (t[303] & ~t[304]);
  assign t[272] = (t[305] & ~t[306]);
  assign t[273] = (t[307] & ~t[308]);
  assign t[274] = (t[309] & ~t[310]);
  assign t[275] = (t[311] & ~t[312]);
  assign t[276] = (t[313] & ~t[314]);
  assign t[277] = (t[315] & ~t[316]);
  assign t[278] = (t[317] & ~t[318]);
  assign t[279] = (t[319] & ~t[320]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = ~(t[49]);
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = t[347] ^ x[4];
  assign t[294] = t[348] ^ x[3];
  assign t[295] = t[349] ^ x[9];
  assign t[296] = t[350] ^ x[8];
  assign t[297] = t[351] ^ x[12];
  assign t[298] = t[352] ^ x[11];
  assign t[299] = t[353] ^ x[15];
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[14];
  assign t[301] = t[355] ^ x[18];
  assign t[302] = t[356] ^ x[17];
  assign t[303] = t[357] ^ x[21];
  assign t[304] = t[358] ^ x[20];
  assign t[305] = t[359] ^ x[24];
  assign t[306] = t[360] ^ x[23];
  assign t[307] = t[361] ^ x[27];
  assign t[308] = t[362] ^ x[26];
  assign t[309] = t[363] ^ x[30];
  assign t[30] = ~(t[214]);
  assign t[310] = t[364] ^ x[29];
  assign t[311] = t[365] ^ x[33];
  assign t[312] = t[366] ^ x[32];
  assign t[313] = t[367] ^ x[36];
  assign t[314] = t[368] ^ x[35];
  assign t[315] = t[369] ^ x[39];
  assign t[316] = t[370] ^ x[38];
  assign t[317] = t[371] ^ x[42];
  assign t[318] = t[372] ^ x[41];
  assign t[319] = t[373] ^ x[45];
  assign t[31] = ~(t[215]);
  assign t[320] = t[374] ^ x[44];
  assign t[321] = t[375] ^ x[48];
  assign t[322] = t[376] ^ x[47];
  assign t[323] = t[377] ^ x[51];
  assign t[324] = t[378] ^ x[50];
  assign t[325] = t[379] ^ x[54];
  assign t[326] = t[380] ^ x[53];
  assign t[327] = t[381] ^ x[57];
  assign t[328] = t[382] ^ x[56];
  assign t[329] = t[383] ^ x[60];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[59];
  assign t[331] = t[385] ^ x[67];
  assign t[332] = t[386] ^ x[66];
  assign t[333] = t[387] ^ x[80];
  assign t[334] = t[388] ^ x[79];
  assign t[335] = t[389] ^ x[83];
  assign t[336] = t[390] ^ x[82];
  assign t[337] = t[391] ^ x[86];
  assign t[338] = t[392] ^ x[85];
  assign t[339] = t[393] ^ x[93];
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[340] = t[394] ^ x[92];
  assign t[341] = t[395] ^ x[96];
  assign t[342] = t[396] ^ x[95];
  assign t[343] = t[397] ^ x[99];
  assign t[344] = t[398] ^ x[98];
  assign t[345] = t[399] ^ x[102];
  assign t[346] = t[400] ^ x[101];
  assign t[347] = (x[2]);
  assign t[348] = (x[2]);
  assign t[349] = (x[7]);
  assign t[34] = t[54] ^ t[55];
  assign t[350] = (x[7]);
  assign t[351] = (x[10]);
  assign t[352] = (x[10]);
  assign t[353] = (x[13]);
  assign t[354] = (x[13]);
  assign t[355] = (x[16]);
  assign t[356] = (x[16]);
  assign t[357] = (x[19]);
  assign t[358] = (x[19]);
  assign t[359] = (x[22]);
  assign t[35] = t[56] ^ t[43];
  assign t[360] = (x[22]);
  assign t[361] = (x[25]);
  assign t[362] = (x[25]);
  assign t[363] = (x[28]);
  assign t[364] = (x[28]);
  assign t[365] = (x[31]);
  assign t[366] = (x[31]);
  assign t[367] = (x[34]);
  assign t[368] = (x[34]);
  assign t[369] = (x[37]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[37]);
  assign t[371] = (x[40]);
  assign t[372] = (x[40]);
  assign t[373] = (x[43]);
  assign t[374] = (x[43]);
  assign t[375] = (x[46]);
  assign t[376] = (x[46]);
  assign t[377] = (x[49]);
  assign t[378] = (x[49]);
  assign t[379] = (x[52]);
  assign t[37] = t[59] ^ t[33];
  assign t[380] = (x[52]);
  assign t[381] = (x[55]);
  assign t[382] = (x[55]);
  assign t[383] = (x[58]);
  assign t[384] = (x[58]);
  assign t[385] = (x[65]);
  assign t[386] = (x[65]);
  assign t[387] = (x[78]);
  assign t[388] = (x[78]);
  assign t[389] = (x[81]);
  assign t[38] = ~(t[25] ^ t[60]);
  assign t[390] = (x[81]);
  assign t[391] = (x[84]);
  assign t[392] = (x[84]);
  assign t[393] = (x[91]);
  assign t[394] = (x[91]);
  assign t[395] = (x[94]);
  assign t[396] = (x[94]);
  assign t[397] = (x[97]);
  assign t[398] = (x[97]);
  assign t[399] = (x[100]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[100]);
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] & t[68];
  assign t[43] = t[216] ^ t[69];
  assign t[44] = t[57] ^ t[70];
  assign t[45] = t[71];
  assign t[46] = t[72] ^ t[73];
  assign t[47] = ~(t[74] & t[75]);
  assign t[48] = t[217] | t[76];
  assign t[49] = ~(t[77]);
  assign t[4] = t[8] ? t[9] : t[212];
  assign t[50] = ~(t[216]);
  assign t[51] = ~(t[78] & t[218]);
  assign t[52] = t[79] ^ t[80];
  assign t[53] = ~(t[81] ^ t[82]);
  assign t[54] = t[65] ^ t[83];
  assign t[55] = t[84] & t[85];
  assign t[56] = t[215] ^ t[86];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] & t[90];
  assign t[59] = ~(t[91] ^ t[92]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] ^ t[73];
  assign t[61] = t[94] ? t[95] : t[219];
  assign t[62] = t[94] ? t[96] : t[220];
  assign t[63] = t[97] ^ t[98];
  assign t[64] = t[99] & t[100];
  assign t[65] = t[8] ? t[101] : t[221];
  assign t[66] = t[8] ? t[102] : t[222];
  assign t[67] = ~(t[83]);
  assign t[68] = t[8] ? t[103] : t[223];
  assign t[69] = t[8] ? t[104] : t[224];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[105] & t[106];
  assign t[71] = t[8] ? t[107] : t[225];
  assign t[72] = t[108] ^ t[109];
  assign t[73] = t[110] & t[111];
  assign t[74] = ~(t[76] & t[112]);
  assign t[75] = ~(t[226] ^ t[113]);
  assign t[76] = ~(t[114] & t[115]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[227]);
  assign t[79] = t[116] ^ t[98];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] ^ t[70];
  assign t[81] = t[118] ^ t[60];
  assign t[82] = t[62] ^ t[119];
  assign t[83] = t[8] ? t[120] : t[228];
  assign t[84] = ~(t[54] ^ t[121]);
  assign t[85] = t[122] ^ t[68];
  assign t[86] = t[8] ? t[123] : t[229];
  assign t[87] = t[124] & t[125];
  assign t[88] = t[126] & t[127];
  assign t[89] = ~(t[87] ^ t[128]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[131] ^ t[24];
  assign t[92] = ~(t[132] ^ t[80]);
  assign t[93] = t[133] ^ t[134];
  assign t[94] = ~(t[15]);
  assign t[95] = t[219] ^ t[135];
  assign t[96] = t[220] ^ t[136];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[139] & t[140];
  assign t[99] = ~(t[97] ^ t[141]);
  assign t[9] = t[212] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [116:0] x;
 output y;

 wire [409:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[53] ^ t[141];
  assign t[101] = t[142] ^ t[143];
  assign t[102] = t[144] ^ t[145];
  assign t[103] = t[130] ^ t[60];
  assign t[104] = t[42] ^ t[86];
  assign t[105] = t[146] ^ t[147];
  assign t[106] = t[8] ? t[148] : t[233];
  assign t[107] = ~(t[70] ^ t[98]);
  assign t[108] = t[65] ^ t[149];
  assign t[109] = t[8] ? t[150] : t[234];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[151] ^ t[64];
  assign t[111] = t[152] & t[153];
  assign t[112] = ~(t[154] & t[155]);
  assign t[113] = t[156] ^ t[235];
  assign t[114] = ~(t[229]);
  assign t[115] = t[157] & t[156];
  assign t[116] = t[8] ? t[158] : t[236];
  assign t[117] = ~(t[83]);
  assign t[118] = t[230] ^ t[159];
  assign t[119] = ~t[160];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[161] & t[162];
  assign t[121] = t[8] ? t[163] : t[237];
  assign t[122] = ~(t[88] ^ t[164]);
  assign t[123] = t[79] ^ t[165];
  assign t[124] = t[22] ^ t[166];
  assign t[125] = ~(t[100] ^ t[103]);
  assign t[126] = t[93] ^ t[119];
  assign t[127] = t[28] ? x[56] : x[55];
  assign t[128] = ~(t[165]);
  assign t[129] = ~(t[116]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[116] ^ t[83];
  assign t[131] = t[167] ^ t[146];
  assign t[132] = t[168] ^ t[169];
  assign t[133] = t[8] ? t[170] : t[238];
  assign t[134] = t[8] ? t[171] : t[239];
  assign t[135] = t[231] ^ t[172];
  assign t[136] = t[232] ^ t[173];
  assign t[137] = t[174] & t[175];
  assign t[138] = t[176] & t[149];
  assign t[139] = ~(t[137] ^ t[177]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[178] ^ t[179];
  assign t[141] = t[97] ^ t[180];
  assign t[142] = t[181] ^ t[167];
  assign t[143] = t[182] & t[183];
  assign t[144] = t[181] ^ t[146];
  assign t[145] = t[184] & t[185];
  assign t[146] = t[186] ? t[187] : t[240];
  assign t[147] = t[168] ^ t[143];
  assign t[148] = t[233] ^ t[188];
  assign t[149] = t[8] ? t[189] : t[241];
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[234] ^ t[190];
  assign t[151] = t[191] & t[192];
  assign t[152] = ~(t[126] ^ t[110]);
  assign t[153] = t[81] ^ t[95];
  assign t[154] = ~(t[157] | t[156]);
  assign t[155] = ~(t[193] | t[114]);
  assign t[156] = ~(t[242]);
  assign t[157] = ~(t[235]);
  assign t[158] = t[236] ^ t[194];
  assign t[159] = t[8] ? t[195] : t[243];
  assign t[15] = ~(t[27]);
  assign t[160] = t[8] ? t[196] : t[244];
  assign t[161] = ~(t[151] ^ t[197]);
  assign t[162] = t[63] ^ t[198];
  assign t[163] = t[237] ^ t[199];
  assign t[164] = t[54] ^ t[116];
  assign t[165] = t[118] ^ t[83];
  assign t[166] = t[178] ^ t[138];
  assign t[167] = t[186] ? t[200] : t[245];
  assign t[168] = t[201] ^ t[145];
  assign t[169] = t[202] & t[203];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[238] ^ t[204];
  assign t[171] = t[239] ^ t[205];
  assign t[172] = t[206] ? x[82] : x[81];
  assign t[173] = t[77] ? x[84] : x[83];
  assign t[174] = ~(t[179]);
  assign t[175] = ~(t[106]);
  assign t[176] = ~(t[96]);
  assign t[177] = t[65] ^ t[106];
  assign t[178] = t[106] ^ t[97];
  assign t[179] = t[149] ^ t[96];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[98] ^ t[71];
  assign t[181] = t[186] ? t[207] : t[246];
  assign t[182] = ~(t[142] ^ t[168]);
  assign t[183] = t[131] ^ t[185];
  assign t[184] = ~(t[167]);
  assign t[185] = t[186] ? t[208] : t[247];
  assign t[186] = ~(t[15]);
  assign t[187] = t[240] ^ t[209];
  assign t[188] = t[206] ? x[92] : x[91];
  assign t[189] = t[241] ^ t[210];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[77] ? x[94] : x[93];
  assign t[191] = ~(t[198]);
  assign t[192] = ~(t[93]);
  assign t[193] = ~(t[226]);
  assign t[194] = t[28] ? x[96] : x[95];
  assign t[195] = t[243] ^ t[211];
  assign t[196] = t[244] ^ t[212];
  assign t[197] = t[81] ^ t[93];
  assign t[198] = t[95] ^ t[119];
  assign t[199] = t[28] ? x[98] : x[97];
  assign t[19] = ~(t[33] ^ t[34]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[245] ^ t[213];
  assign t[201] = t[214] & t[215];
  assign t[202] = ~(t[201] ^ t[216]);
  assign t[203] = t[144] ^ t[217];
  assign t[204] = t[77] ? x[100] : x[99];
  assign t[205] = t[77] ? x[102] : x[101];
  assign t[206] = ~(t[49]);
  assign t[207] = t[246] ^ t[218];
  assign t[208] = t[247] ^ t[219];
  assign t[209] = t[220] ? x[104] : x[103];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[206] ? x[106] : x[105];
  assign t[211] = t[28] ? x[108] : x[107];
  assign t[212] = t[28] ? x[110] : x[109];
  assign t[213] = t[220] ? x[112] : x[111];
  assign t[214] = ~(t[217]);
  assign t[215] = ~(t[181]);
  assign t[216] = t[131] ^ t[181];
  assign t[217] = t[185] ^ t[167];
  assign t[218] = t[220] ? x[114] : x[113];
  assign t[219] = t[220] ? x[116] : x[115];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = ~(t[49]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[39] ^ t[40]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = (t[266]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (t[267]);
  assign t[241] = (t[268]);
  assign t[242] = (t[269]);
  assign t[243] = (t[270]);
  assign t[244] = (t[271]);
  assign t[245] = (t[272]);
  assign t[246] = (t[273]);
  assign t[247] = (t[274]);
  assign t[248] = t[275] ^ x[4];
  assign t[249] = t[276] ^ x[9];
  assign t[24] = ~(t[43] ^ t[21]);
  assign t[250] = t[277] ^ x[12];
  assign t[251] = t[278] ^ x[15];
  assign t[252] = t[279] ^ x[18];
  assign t[253] = t[280] ^ x[21];
  assign t[254] = t[281] ^ x[24];
  assign t[255] = t[282] ^ x[27];
  assign t[256] = t[283] ^ x[30];
  assign t[257] = t[284] ^ x[33];
  assign t[258] = t[285] ^ x[36];
  assign t[259] = t[286] ^ x[39];
  assign t[25] = t[44] ^ t[45];
  assign t[260] = t[287] ^ x[42];
  assign t[261] = t[288] ^ x[45];
  assign t[262] = t[289] ^ x[48];
  assign t[263] = t[290] ^ x[51];
  assign t[264] = t[291] ^ x[54];
  assign t[265] = t[292] ^ x[59];
  assign t[266] = t[293] ^ x[62];
  assign t[267] = t[294] ^ x[65];
  assign t[268] = t[295] ^ x[68];
  assign t[269] = t[296] ^ x[71];
  assign t[26] = ~(t[35] ^ t[46]);
  assign t[270] = t[297] ^ x[74];
  assign t[271] = t[298] ^ x[77];
  assign t[272] = t[299] ^ x[80];
  assign t[273] = t[300] ^ x[87];
  assign t[274] = t[301] ^ x[90];
  assign t[275] = (t[302] & ~t[303]);
  assign t[276] = (t[304] & ~t[305]);
  assign t[277] = (t[306] & ~t[307]);
  assign t[278] = (t[308] & ~t[309]);
  assign t[279] = (t[310] & ~t[311]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[312] & ~t[313]);
  assign t[281] = (t[314] & ~t[315]);
  assign t[282] = (t[316] & ~t[317]);
  assign t[283] = (t[318] & ~t[319]);
  assign t[284] = (t[320] & ~t[321]);
  assign t[285] = (t[322] & ~t[323]);
  assign t[286] = (t[324] & ~t[325]);
  assign t[287] = (t[326] & ~t[327]);
  assign t[288] = (t[328] & ~t[329]);
  assign t[289] = (t[330] & ~t[331]);
  assign t[28] = ~(t[49]);
  assign t[290] = (t[332] & ~t[333]);
  assign t[291] = (t[334] & ~t[335]);
  assign t[292] = (t[336] & ~t[337]);
  assign t[293] = (t[338] & ~t[339]);
  assign t[294] = (t[340] & ~t[341]);
  assign t[295] = (t[342] & ~t[343]);
  assign t[296] = (t[344] & ~t[345]);
  assign t[297] = (t[346] & ~t[347]);
  assign t[298] = (t[348] & ~t[349]);
  assign t[299] = (t[350] & ~t[351]);
  assign t[29] = ~(t[222]);
  assign t[2] = ~(t[5]);
  assign t[300] = (t[352] & ~t[353]);
  assign t[301] = (t[354] & ~t[355]);
  assign t[302] = t[356] ^ x[4];
  assign t[303] = t[357] ^ x[3];
  assign t[304] = t[358] ^ x[9];
  assign t[305] = t[359] ^ x[8];
  assign t[306] = t[360] ^ x[12];
  assign t[307] = t[361] ^ x[11];
  assign t[308] = t[362] ^ x[15];
  assign t[309] = t[363] ^ x[14];
  assign t[30] = ~(t[223]);
  assign t[310] = t[364] ^ x[18];
  assign t[311] = t[365] ^ x[17];
  assign t[312] = t[366] ^ x[21];
  assign t[313] = t[367] ^ x[20];
  assign t[314] = t[368] ^ x[24];
  assign t[315] = t[369] ^ x[23];
  assign t[316] = t[370] ^ x[27];
  assign t[317] = t[371] ^ x[26];
  assign t[318] = t[372] ^ x[30];
  assign t[319] = t[373] ^ x[29];
  assign t[31] = ~(t[224]);
  assign t[320] = t[374] ^ x[33];
  assign t[321] = t[375] ^ x[32];
  assign t[322] = t[376] ^ x[36];
  assign t[323] = t[377] ^ x[35];
  assign t[324] = t[378] ^ x[39];
  assign t[325] = t[379] ^ x[38];
  assign t[326] = t[380] ^ x[42];
  assign t[327] = t[381] ^ x[41];
  assign t[328] = t[382] ^ x[45];
  assign t[329] = t[383] ^ x[44];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[48];
  assign t[331] = t[385] ^ x[47];
  assign t[332] = t[386] ^ x[51];
  assign t[333] = t[387] ^ x[50];
  assign t[334] = t[388] ^ x[54];
  assign t[335] = t[389] ^ x[53];
  assign t[336] = t[390] ^ x[59];
  assign t[337] = t[391] ^ x[58];
  assign t[338] = t[392] ^ x[62];
  assign t[339] = t[393] ^ x[61];
  assign t[33] = t[52] ^ t[14];
  assign t[340] = t[394] ^ x[65];
  assign t[341] = t[395] ^ x[64];
  assign t[342] = t[396] ^ x[68];
  assign t[343] = t[397] ^ x[67];
  assign t[344] = t[398] ^ x[71];
  assign t[345] = t[399] ^ x[70];
  assign t[346] = t[400] ^ x[74];
  assign t[347] = t[401] ^ x[73];
  assign t[348] = t[402] ^ x[77];
  assign t[349] = t[403] ^ x[76];
  assign t[34] = ~(t[53] ^ t[43]);
  assign t[350] = t[404] ^ x[80];
  assign t[351] = t[405] ^ x[79];
  assign t[352] = t[406] ^ x[87];
  assign t[353] = t[407] ^ x[86];
  assign t[354] = t[408] ^ x[90];
  assign t[355] = t[409] ^ x[89];
  assign t[356] = (x[2]);
  assign t[357] = (x[2]);
  assign t[358] = (x[7]);
  assign t[359] = (x[7]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[10]);
  assign t[361] = (x[10]);
  assign t[362] = (x[13]);
  assign t[363] = (x[13]);
  assign t[364] = (x[16]);
  assign t[365] = (x[16]);
  assign t[366] = (x[19]);
  assign t[367] = (x[19]);
  assign t[368] = (x[22]);
  assign t[369] = (x[22]);
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[370] = (x[25]);
  assign t[371] = (x[25]);
  assign t[372] = (x[28]);
  assign t[373] = (x[28]);
  assign t[374] = (x[31]);
  assign t[375] = (x[31]);
  assign t[376] = (x[34]);
  assign t[377] = (x[34]);
  assign t[378] = (x[37]);
  assign t[379] = (x[37]);
  assign t[37] = t[225] ^ t[58];
  assign t[380] = (x[40]);
  assign t[381] = (x[40]);
  assign t[382] = (x[43]);
  assign t[383] = (x[43]);
  assign t[384] = (x[46]);
  assign t[385] = (x[46]);
  assign t[386] = (x[49]);
  assign t[387] = (x[49]);
  assign t[388] = (x[52]);
  assign t[389] = (x[52]);
  assign t[38] = t[59] ^ t[60];
  assign t[390] = (x[57]);
  assign t[391] = (x[57]);
  assign t[392] = (x[60]);
  assign t[393] = (x[60]);
  assign t[394] = (x[63]);
  assign t[395] = (x[63]);
  assign t[396] = (x[66]);
  assign t[397] = (x[66]);
  assign t[398] = (x[69]);
  assign t[399] = (x[69]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[72]);
  assign t[401] = (x[72]);
  assign t[402] = (x[75]);
  assign t[403] = (x[75]);
  assign t[404] = (x[78]);
  assign t[405] = (x[78]);
  assign t[406] = (x[85]);
  assign t[407] = (x[85]);
  assign t[408] = (x[88]);
  assign t[409] = (x[88]);
  assign t[40] = ~(t[41] ^ t[46]);
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[67] ^ t[35]);
  assign t[44] = ~(t[68] ^ t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] ^ t[73];
  assign t[47] = ~(t[74] & t[75]);
  assign t[48] = t[226] | t[76];
  assign t[49] = ~(t[77]);
  assign t[4] = t[8] ? t[9] : t[221];
  assign t[50] = ~(t[225]);
  assign t[51] = ~(t[78] & t[227]);
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] ^ t[37];
  assign t[55] = t[59] ^ t[84];
  assign t[56] = t[85] ^ t[44];
  assign t[57] = ~(t[21] ^ t[86]);
  assign t[58] = t[8] ? t[87] : t[228];
  assign t[59] = t[88] ^ t[80];
  assign t[5] = ~(t[10]);
  assign t[60] = t[89] & t[90];
  assign t[61] = t[21] ^ t[52];
  assign t[62] = ~(t[91] ^ t[92]);
  assign t[63] = t[93] ^ t[72];
  assign t[64] = t[94] & t[95];
  assign t[65] = t[96] ^ t[97];
  assign t[66] = t[98] ^ t[99];
  assign t[67] = ~(t[100] ^ t[101]);
  assign t[68] = t[102] ^ t[103];
  assign t[69] = ~(t[104] ^ t[105]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[106] ^ t[96];
  assign t[71] = t[107] & t[108];
  assign t[72] = t[109];
  assign t[73] = t[110] ^ t[111];
  assign t[74] = ~(t[76] & t[112]);
  assign t[75] = ~(t[229] ^ t[113]);
  assign t[76] = ~(t[114] & t[115]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[230]);
  assign t[79] = t[116] ^ t[37];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] & t[118];
  assign t[81] = t[119] ^ t[72];
  assign t[82] = t[110] ^ t[120];
  assign t[83] = t[224] ^ t[121];
  assign t[84] = t[122] & t[123];
  assign t[85] = ~(t[124] ^ t[125]);
  assign t[86] = t[126] ^ t[111];
  assign t[87] = t[228] ^ t[127];
  assign t[88] = t[128] & t[129];
  assign t[89] = ~(t[130] ^ t[59]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[54] ^ t[118];
  assign t[91] = ~(t[45] ^ t[105]);
  assign t[92] = t[131] ^ t[132];
  assign t[93] = t[133];
  assign t[94] = ~(t[119]);
  assign t[95] = t[134];
  assign t[96] = t[8] ? t[135] : t[231];
  assign t[97] = t[8] ? t[136] : t[232];
  assign t[98] = t[137] ^ t[138];
  assign t[99] = t[139] & t[140];
  assign t[9] = t[221] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [116:0] x;
 output y;

 wire [409:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[53] ^ t[141];
  assign t[101] = t[142] ^ t[143];
  assign t[102] = t[144] ^ t[145];
  assign t[103] = t[130] ^ t[60];
  assign t[104] = t[42] ^ t[86];
  assign t[105] = t[146] ^ t[147];
  assign t[106] = t[8] ? t[148] : t[233];
  assign t[107] = ~(t[70] ^ t[98]);
  assign t[108] = t[65] ^ t[149];
  assign t[109] = t[8] ? t[150] : t[234];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[151] ^ t[64];
  assign t[111] = t[152] & t[153];
  assign t[112] = ~(t[154] & t[155]);
  assign t[113] = t[156] ^ t[235];
  assign t[114] = ~(t[229]);
  assign t[115] = t[157] & t[156];
  assign t[116] = t[8] ? t[158] : t[236];
  assign t[117] = ~(t[83]);
  assign t[118] = t[230] ^ t[159];
  assign t[119] = ~t[160];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[161] & t[162];
  assign t[121] = t[8] ? t[163] : t[237];
  assign t[122] = ~(t[88] ^ t[164]);
  assign t[123] = t[79] ^ t[165];
  assign t[124] = t[22] ^ t[166];
  assign t[125] = ~(t[100] ^ t[103]);
  assign t[126] = t[93] ^ t[119];
  assign t[127] = t[28] ? x[56] : x[55];
  assign t[128] = ~(t[165]);
  assign t[129] = ~(t[116]);
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[116] ^ t[83];
  assign t[131] = t[167] ^ t[146];
  assign t[132] = t[168] ^ t[169];
  assign t[133] = t[8] ? t[170] : t[238];
  assign t[134] = t[8] ? t[171] : t[239];
  assign t[135] = t[231] ^ t[172];
  assign t[136] = t[232] ^ t[173];
  assign t[137] = t[174] & t[175];
  assign t[138] = t[176] & t[149];
  assign t[139] = ~(t[137] ^ t[177]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[178] ^ t[179];
  assign t[141] = t[97] ^ t[180];
  assign t[142] = t[181] ^ t[167];
  assign t[143] = t[182] & t[183];
  assign t[144] = t[181] ^ t[146];
  assign t[145] = t[184] & t[185];
  assign t[146] = t[186] ? t[187] : t[240];
  assign t[147] = t[168] ^ t[143];
  assign t[148] = t[233] ^ t[188];
  assign t[149] = t[8] ? t[189] : t[241];
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[234] ^ t[190];
  assign t[151] = t[191] & t[192];
  assign t[152] = ~(t[126] ^ t[110]);
  assign t[153] = t[81] ^ t[95];
  assign t[154] = ~(t[157] | t[156]);
  assign t[155] = ~(t[193] | t[114]);
  assign t[156] = ~(t[242]);
  assign t[157] = ~(t[235]);
  assign t[158] = t[236] ^ t[194];
  assign t[159] = t[8] ? t[195] : t[243];
  assign t[15] = ~(t[27]);
  assign t[160] = t[8] ? t[196] : t[244];
  assign t[161] = ~(t[151] ^ t[197]);
  assign t[162] = t[63] ^ t[198];
  assign t[163] = t[237] ^ t[199];
  assign t[164] = t[54] ^ t[116];
  assign t[165] = t[118] ^ t[83];
  assign t[166] = t[178] ^ t[138];
  assign t[167] = t[186] ? t[200] : t[245];
  assign t[168] = t[201] ^ t[145];
  assign t[169] = t[202] & t[203];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[238] ^ t[204];
  assign t[171] = t[239] ^ t[205];
  assign t[172] = t[206] ? x[82] : x[81];
  assign t[173] = t[77] ? x[84] : x[83];
  assign t[174] = ~(t[179]);
  assign t[175] = ~(t[106]);
  assign t[176] = ~(t[96]);
  assign t[177] = t[65] ^ t[106];
  assign t[178] = t[106] ^ t[97];
  assign t[179] = t[149] ^ t[96];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[98] ^ t[71];
  assign t[181] = t[186] ? t[207] : t[246];
  assign t[182] = ~(t[142] ^ t[168]);
  assign t[183] = t[131] ^ t[185];
  assign t[184] = ~(t[167]);
  assign t[185] = t[186] ? t[208] : t[247];
  assign t[186] = ~(t[15]);
  assign t[187] = t[240] ^ t[209];
  assign t[188] = t[206] ? x[92] : x[91];
  assign t[189] = t[241] ^ t[210];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[77] ? x[94] : x[93];
  assign t[191] = ~(t[198]);
  assign t[192] = ~(t[93]);
  assign t[193] = ~(t[226]);
  assign t[194] = t[28] ? x[96] : x[95];
  assign t[195] = t[243] ^ t[211];
  assign t[196] = t[244] ^ t[212];
  assign t[197] = t[81] ^ t[93];
  assign t[198] = t[95] ^ t[119];
  assign t[199] = t[28] ? x[98] : x[97];
  assign t[19] = ~(t[33] ^ t[34]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[245] ^ t[213];
  assign t[201] = t[214] & t[215];
  assign t[202] = ~(t[201] ^ t[216]);
  assign t[203] = t[144] ^ t[217];
  assign t[204] = t[77] ? x[100] : x[99];
  assign t[205] = t[77] ? x[102] : x[101];
  assign t[206] = ~(t[49]);
  assign t[207] = t[246] ^ t[218];
  assign t[208] = t[247] ^ t[219];
  assign t[209] = t[220] ? x[104] : x[103];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[206] ? x[106] : x[105];
  assign t[211] = t[28] ? x[108] : x[107];
  assign t[212] = t[28] ? x[110] : x[109];
  assign t[213] = t[220] ? x[112] : x[111];
  assign t[214] = ~(t[217]);
  assign t[215] = ~(t[181]);
  assign t[216] = t[131] ^ t[181];
  assign t[217] = t[185] ^ t[167];
  assign t[218] = t[220] ? x[114] : x[113];
  assign t[219] = t[220] ? x[116] : x[115];
  assign t[21] = t[37] ^ t[38];
  assign t[220] = ~(t[49]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[39] ^ t[40]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = (t[266]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (t[267]);
  assign t[241] = (t[268]);
  assign t[242] = (t[269]);
  assign t[243] = (t[270]);
  assign t[244] = (t[271]);
  assign t[245] = (t[272]);
  assign t[246] = (t[273]);
  assign t[247] = (t[274]);
  assign t[248] = t[275] ^ x[4];
  assign t[249] = t[276] ^ x[9];
  assign t[24] = ~(t[43] ^ t[21]);
  assign t[250] = t[277] ^ x[12];
  assign t[251] = t[278] ^ x[15];
  assign t[252] = t[279] ^ x[18];
  assign t[253] = t[280] ^ x[21];
  assign t[254] = t[281] ^ x[24];
  assign t[255] = t[282] ^ x[27];
  assign t[256] = t[283] ^ x[30];
  assign t[257] = t[284] ^ x[33];
  assign t[258] = t[285] ^ x[36];
  assign t[259] = t[286] ^ x[39];
  assign t[25] = t[44] ^ t[45];
  assign t[260] = t[287] ^ x[42];
  assign t[261] = t[288] ^ x[45];
  assign t[262] = t[289] ^ x[48];
  assign t[263] = t[290] ^ x[51];
  assign t[264] = t[291] ^ x[54];
  assign t[265] = t[292] ^ x[59];
  assign t[266] = t[293] ^ x[62];
  assign t[267] = t[294] ^ x[65];
  assign t[268] = t[295] ^ x[68];
  assign t[269] = t[296] ^ x[71];
  assign t[26] = ~(t[35] ^ t[46]);
  assign t[270] = t[297] ^ x[74];
  assign t[271] = t[298] ^ x[77];
  assign t[272] = t[299] ^ x[80];
  assign t[273] = t[300] ^ x[87];
  assign t[274] = t[301] ^ x[90];
  assign t[275] = (t[302] & ~t[303]);
  assign t[276] = (t[304] & ~t[305]);
  assign t[277] = (t[306] & ~t[307]);
  assign t[278] = (t[308] & ~t[309]);
  assign t[279] = (t[310] & ~t[311]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[312] & ~t[313]);
  assign t[281] = (t[314] & ~t[315]);
  assign t[282] = (t[316] & ~t[317]);
  assign t[283] = (t[318] & ~t[319]);
  assign t[284] = (t[320] & ~t[321]);
  assign t[285] = (t[322] & ~t[323]);
  assign t[286] = (t[324] & ~t[325]);
  assign t[287] = (t[326] & ~t[327]);
  assign t[288] = (t[328] & ~t[329]);
  assign t[289] = (t[330] & ~t[331]);
  assign t[28] = ~(t[49]);
  assign t[290] = (t[332] & ~t[333]);
  assign t[291] = (t[334] & ~t[335]);
  assign t[292] = (t[336] & ~t[337]);
  assign t[293] = (t[338] & ~t[339]);
  assign t[294] = (t[340] & ~t[341]);
  assign t[295] = (t[342] & ~t[343]);
  assign t[296] = (t[344] & ~t[345]);
  assign t[297] = (t[346] & ~t[347]);
  assign t[298] = (t[348] & ~t[349]);
  assign t[299] = (t[350] & ~t[351]);
  assign t[29] = ~(t[222]);
  assign t[2] = ~(t[5]);
  assign t[300] = (t[352] & ~t[353]);
  assign t[301] = (t[354] & ~t[355]);
  assign t[302] = t[356] ^ x[4];
  assign t[303] = t[357] ^ x[3];
  assign t[304] = t[358] ^ x[9];
  assign t[305] = t[359] ^ x[8];
  assign t[306] = t[360] ^ x[12];
  assign t[307] = t[361] ^ x[11];
  assign t[308] = t[362] ^ x[15];
  assign t[309] = t[363] ^ x[14];
  assign t[30] = ~(t[223]);
  assign t[310] = t[364] ^ x[18];
  assign t[311] = t[365] ^ x[17];
  assign t[312] = t[366] ^ x[21];
  assign t[313] = t[367] ^ x[20];
  assign t[314] = t[368] ^ x[24];
  assign t[315] = t[369] ^ x[23];
  assign t[316] = t[370] ^ x[27];
  assign t[317] = t[371] ^ x[26];
  assign t[318] = t[372] ^ x[30];
  assign t[319] = t[373] ^ x[29];
  assign t[31] = ~(t[224]);
  assign t[320] = t[374] ^ x[33];
  assign t[321] = t[375] ^ x[32];
  assign t[322] = t[376] ^ x[36];
  assign t[323] = t[377] ^ x[35];
  assign t[324] = t[378] ^ x[39];
  assign t[325] = t[379] ^ x[38];
  assign t[326] = t[380] ^ x[42];
  assign t[327] = t[381] ^ x[41];
  assign t[328] = t[382] ^ x[45];
  assign t[329] = t[383] ^ x[44];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[48];
  assign t[331] = t[385] ^ x[47];
  assign t[332] = t[386] ^ x[51];
  assign t[333] = t[387] ^ x[50];
  assign t[334] = t[388] ^ x[54];
  assign t[335] = t[389] ^ x[53];
  assign t[336] = t[390] ^ x[59];
  assign t[337] = t[391] ^ x[58];
  assign t[338] = t[392] ^ x[62];
  assign t[339] = t[393] ^ x[61];
  assign t[33] = t[52] ^ t[14];
  assign t[340] = t[394] ^ x[65];
  assign t[341] = t[395] ^ x[64];
  assign t[342] = t[396] ^ x[68];
  assign t[343] = t[397] ^ x[67];
  assign t[344] = t[398] ^ x[71];
  assign t[345] = t[399] ^ x[70];
  assign t[346] = t[400] ^ x[74];
  assign t[347] = t[401] ^ x[73];
  assign t[348] = t[402] ^ x[77];
  assign t[349] = t[403] ^ x[76];
  assign t[34] = ~(t[53] ^ t[43]);
  assign t[350] = t[404] ^ x[80];
  assign t[351] = t[405] ^ x[79];
  assign t[352] = t[406] ^ x[87];
  assign t[353] = t[407] ^ x[86];
  assign t[354] = t[408] ^ x[90];
  assign t[355] = t[409] ^ x[89];
  assign t[356] = (x[2]);
  assign t[357] = (x[2]);
  assign t[358] = (x[7]);
  assign t[359] = (x[7]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[10]);
  assign t[361] = (x[10]);
  assign t[362] = (x[13]);
  assign t[363] = (x[13]);
  assign t[364] = (x[16]);
  assign t[365] = (x[16]);
  assign t[366] = (x[19]);
  assign t[367] = (x[19]);
  assign t[368] = (x[22]);
  assign t[369] = (x[22]);
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[370] = (x[25]);
  assign t[371] = (x[25]);
  assign t[372] = (x[28]);
  assign t[373] = (x[28]);
  assign t[374] = (x[31]);
  assign t[375] = (x[31]);
  assign t[376] = (x[34]);
  assign t[377] = (x[34]);
  assign t[378] = (x[37]);
  assign t[379] = (x[37]);
  assign t[37] = t[225] ^ t[58];
  assign t[380] = (x[40]);
  assign t[381] = (x[40]);
  assign t[382] = (x[43]);
  assign t[383] = (x[43]);
  assign t[384] = (x[46]);
  assign t[385] = (x[46]);
  assign t[386] = (x[49]);
  assign t[387] = (x[49]);
  assign t[388] = (x[52]);
  assign t[389] = (x[52]);
  assign t[38] = t[59] ^ t[60];
  assign t[390] = (x[57]);
  assign t[391] = (x[57]);
  assign t[392] = (x[60]);
  assign t[393] = (x[60]);
  assign t[394] = (x[63]);
  assign t[395] = (x[63]);
  assign t[396] = (x[66]);
  assign t[397] = (x[66]);
  assign t[398] = (x[69]);
  assign t[399] = (x[69]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[72]);
  assign t[401] = (x[72]);
  assign t[402] = (x[75]);
  assign t[403] = (x[75]);
  assign t[404] = (x[78]);
  assign t[405] = (x[78]);
  assign t[406] = (x[85]);
  assign t[407] = (x[85]);
  assign t[408] = (x[88]);
  assign t[409] = (x[88]);
  assign t[40] = ~(t[41] ^ t[46]);
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[67] ^ t[35]);
  assign t[44] = ~(t[68] ^ t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] ^ t[73];
  assign t[47] = ~(t[74] & t[75]);
  assign t[48] = t[226] | t[76];
  assign t[49] = ~(t[77]);
  assign t[4] = t[8] ? t[9] : t[221];
  assign t[50] = ~(t[225]);
  assign t[51] = ~(t[78] & t[227]);
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] ^ t[37];
  assign t[55] = t[59] ^ t[84];
  assign t[56] = t[85] ^ t[44];
  assign t[57] = ~(t[21] ^ t[86]);
  assign t[58] = t[8] ? t[87] : t[228];
  assign t[59] = t[88] ^ t[80];
  assign t[5] = ~(t[10]);
  assign t[60] = t[89] & t[90];
  assign t[61] = t[21] ^ t[52];
  assign t[62] = ~(t[91] ^ t[92]);
  assign t[63] = t[93] ^ t[72];
  assign t[64] = t[94] & t[95];
  assign t[65] = t[96] ^ t[97];
  assign t[66] = t[98] ^ t[99];
  assign t[67] = ~(t[100] ^ t[101]);
  assign t[68] = t[102] ^ t[103];
  assign t[69] = ~(t[104] ^ t[105]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[106] ^ t[96];
  assign t[71] = t[107] & t[108];
  assign t[72] = t[109];
  assign t[73] = t[110] ^ t[111];
  assign t[74] = ~(t[76] & t[112]);
  assign t[75] = ~(t[229] ^ t[113]);
  assign t[76] = ~(t[114] & t[115]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[230]);
  assign t[79] = t[116] ^ t[37];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] & t[118];
  assign t[81] = t[119] ^ t[72];
  assign t[82] = t[110] ^ t[120];
  assign t[83] = t[224] ^ t[121];
  assign t[84] = t[122] & t[123];
  assign t[85] = ~(t[124] ^ t[125]);
  assign t[86] = t[126] ^ t[111];
  assign t[87] = t[228] ^ t[127];
  assign t[88] = t[128] & t[129];
  assign t[89] = ~(t[130] ^ t[59]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[54] ^ t[118];
  assign t[91] = ~(t[45] ^ t[105]);
  assign t[92] = t[131] ^ t[132];
  assign t[93] = t[133];
  assign t[94] = ~(t[119]);
  assign t[95] = t[134];
  assign t[96] = t[8] ? t[135] : t[231];
  assign t[97] = t[8] ? t[136] : t[232];
  assign t[98] = t[137] ^ t[138];
  assign t[99] = t[139] & t[140];
  assign t[9] = t[221] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [116:0] x;
 output y;

 wire [400:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[139] ^ t[132];
  assign t[101] = ~t[140];
  assign t[102] = t[141] ^ t[106];
  assign t[103] = t[142] & t[143];
  assign t[104] = t[8] ? t[144] : t[226];
  assign t[105] = t[123] ^ t[67];
  assign t[106] = t[145] & t[146];
  assign t[107] = t[217] ^ t[147];
  assign t[108] = t[119] ^ t[54];
  assign t[109] = t[148] ^ t[121];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[149] & t[150]);
  assign t[111] = t[151] ^ t[227];
  assign t[112] = ~(t[221]);
  assign t[113] = t[152] & t[151];
  assign t[114] = t[223] ^ t[153];
  assign t[115] = t[88] ? t[154] : t[228];
  assign t[116] = t[224] ^ t[155];
  assign t[117] = t[225] ^ t[156];
  assign t[118] = t[8] ? t[157] : t[229];
  assign t[119] = t[158] ^ t[159];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[222] ^ t[160];
  assign t[121] = t[8] ? t[161] : t[230];
  assign t[122] = t[162] & t[163];
  assign t[123] = t[164];
  assign t[124] = ~(t[86] ^ t[102]);
  assign t[125] = t[65] ^ t[146];
  assign t[126] = t[165] ? x[62] : x[61];
  assign t[127] = t[166] & t[167];
  assign t[128] = ~(t[135] ^ t[90]);
  assign t[129] = t[137] ^ t[79];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[75] ? x[64] : x[63];
  assign t[131] = t[168] & t[169];
  assign t[132] = t[170] & t[171];
  assign t[133] = ~(t[109] ^ t[93]);
  assign t[134] = t[84] ^ t[171];
  assign t[135] = t[77] ^ t[115];
  assign t[136] = t[172] & t[173];
  assign t[137] = t[115] ^ t[57];
  assign t[138] = t[90] ^ t[174];
  assign t[139] = t[148] ^ t[59];
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[8] ? t[175] : t[231];
  assign t[141] = t[176] & t[177];
  assign t[142] = ~(t[141] ^ t[178]);
  assign t[143] = t[105] ^ t[179];
  assign t[144] = t[226] ^ t[180];
  assign t[145] = ~(t[101]);
  assign t[146] = t[181];
  assign t[147] = t[8] ? t[182] : t[232];
  assign t[148] = t[8] ? t[183] : t[233];
  assign t[149] = ~(t[152] | t[151]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[184] | t[112]);
  assign t[151] = ~(t[234]);
  assign t[152] = ~(t[227]);
  assign t[153] = t[165] ? x[78] : x[77];
  assign t[154] = t[228] ^ t[185];
  assign t[155] = t[165] ? x[80] : x[79];
  assign t[156] = t[28] ? x[82] : x[81];
  assign t[157] = t[229] ^ t[186];
  assign t[158] = t[187] & t[188];
  assign t[159] = t[189] & t[120];
  assign t[15] = ~(t[27]);
  assign t[160] = t[8] ? t[190] : t[235];
  assign t[161] = t[230] ^ t[191];
  assign t[162] = ~(t[131] ^ t[192]);
  assign t[163] = t[139] ^ t[193];
  assign t[164] = t[8] ? t[194] : t[236];
  assign t[165] = ~(t[48]);
  assign t[166] = ~(t[195]);
  assign t[167] = ~(t[77]);
  assign t[168] = ~(t[193]);
  assign t[169] = ~(t[148]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[121]);
  assign t[171] = t[8] ? t[196] : t[237];
  assign t[172] = ~(t[158] ^ t[197]);
  assign t[173] = t[198] ^ t[199];
  assign t[174] = t[200] & t[201];
  assign t[175] = t[231] ^ t[202];
  assign t[176] = ~(t[179]);
  assign t[177] = ~(t[123]);
  assign t[178] = t[65] ^ t[123];
  assign t[179] = t[146] ^ t[101];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[75] ? x[93] : x[92];
  assign t[181] = t[8] ? t[203] : t[238];
  assign t[182] = t[232] ^ t[204];
  assign t[183] = t[233] ^ t[205];
  assign t[184] = ~(t[216]);
  assign t[185] = t[165] ? x[98] : x[97];
  assign t[186] = t[28] ? x[100] : x[99];
  assign t[187] = ~(t[199]);
  assign t[188] = ~(t[80]);
  assign t[189] = ~(t[81]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[235] ^ t[206];
  assign t[191] = t[207] ? x[102] : x[101];
  assign t[192] = t[84] ^ t[148];
  assign t[193] = t[171] ^ t[121];
  assign t[194] = t[236] ^ t[208];
  assign t[195] = t[79] ^ t[115];
  assign t[196] = t[237] ^ t[209];
  assign t[197] = t[97] ^ t[80];
  assign t[198] = t[80] ^ t[107];
  assign t[199] = t[120] ^ t[81];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[127] ^ t[210]);
  assign t[201] = t[51] ^ t[195];
  assign t[202] = t[28] ? x[104] : x[103];
  assign t[203] = t[238] ^ t[211];
  assign t[204] = t[28] ? x[106] : x[105];
  assign t[205] = t[207] ? x[108] : x[107];
  assign t[206] = t[28] ? x[110] : x[109];
  assign t[207] = ~(t[48]);
  assign t[208] = t[75] ? x[112] : x[111];
  assign t[209] = t[207] ? x[114] : x[113];
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = t[137] ^ t[77];
  assign t[211] = t[75] ? x[116] : x[115];
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[35]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[38] ^ t[39];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = t[266] ^ x[4];
  assign t[23] = t[22] ^ t[34];
  assign t[240] = t[267] ^ x[9];
  assign t[241] = t[268] ^ x[12];
  assign t[242] = t[269] ^ x[15];
  assign t[243] = t[270] ^ x[18];
  assign t[244] = t[271] ^ x[21];
  assign t[245] = t[272] ^ x[24];
  assign t[246] = t[273] ^ x[27];
  assign t[247] = t[274] ^ x[30];
  assign t[248] = t[275] ^ x[33];
  assign t[249] = t[276] ^ x[36];
  assign t[24] = ~(t[40] ^ t[41]);
  assign t[250] = t[277] ^ x[39];
  assign t[251] = t[278] ^ x[42];
  assign t[252] = t[279] ^ x[45];
  assign t[253] = t[280] ^ x[48];
  assign t[254] = t[281] ^ x[51];
  assign t[255] = t[282] ^ x[54];
  assign t[256] = t[283] ^ x[57];
  assign t[257] = t[284] ^ x[60];
  assign t[258] = t[285] ^ x[67];
  assign t[259] = t[286] ^ x[70];
  assign t[25] = ~(t[42] ^ t[43]);
  assign t[260] = t[287] ^ x[73];
  assign t[261] = t[288] ^ x[76];
  assign t[262] = t[289] ^ x[85];
  assign t[263] = t[290] ^ x[88];
  assign t[264] = t[291] ^ x[91];
  assign t[265] = t[292] ^ x[96];
  assign t[266] = (t[293] & ~t[294]);
  assign t[267] = (t[295] & ~t[296]);
  assign t[268] = (t[297] & ~t[298]);
  assign t[269] = (t[299] & ~t[300]);
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[270] = (t[301] & ~t[302]);
  assign t[271] = (t[303] & ~t[304]);
  assign t[272] = (t[305] & ~t[306]);
  assign t[273] = (t[307] & ~t[308]);
  assign t[274] = (t[309] & ~t[310]);
  assign t[275] = (t[311] & ~t[312]);
  assign t[276] = (t[313] & ~t[314]);
  assign t[277] = (t[315] & ~t[316]);
  assign t[278] = (t[317] & ~t[318]);
  assign t[279] = (t[319] & ~t[320]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = t[347] ^ x[4];
  assign t[294] = t[348] ^ x[3];
  assign t[295] = t[349] ^ x[9];
  assign t[296] = t[350] ^ x[8];
  assign t[297] = t[351] ^ x[12];
  assign t[298] = t[352] ^ x[11];
  assign t[299] = t[353] ^ x[15];
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[14];
  assign t[301] = t[355] ^ x[18];
  assign t[302] = t[356] ^ x[17];
  assign t[303] = t[357] ^ x[21];
  assign t[304] = t[358] ^ x[20];
  assign t[305] = t[359] ^ x[24];
  assign t[306] = t[360] ^ x[23];
  assign t[307] = t[361] ^ x[27];
  assign t[308] = t[362] ^ x[26];
  assign t[309] = t[363] ^ x[30];
  assign t[30] = ~(t[214]);
  assign t[310] = t[364] ^ x[29];
  assign t[311] = t[365] ^ x[33];
  assign t[312] = t[366] ^ x[32];
  assign t[313] = t[367] ^ x[36];
  assign t[314] = t[368] ^ x[35];
  assign t[315] = t[369] ^ x[39];
  assign t[316] = t[370] ^ x[38];
  assign t[317] = t[371] ^ x[42];
  assign t[318] = t[372] ^ x[41];
  assign t[319] = t[373] ^ x[45];
  assign t[31] = ~(t[215]);
  assign t[320] = t[374] ^ x[44];
  assign t[321] = t[375] ^ x[48];
  assign t[322] = t[376] ^ x[47];
  assign t[323] = t[377] ^ x[51];
  assign t[324] = t[378] ^ x[50];
  assign t[325] = t[379] ^ x[54];
  assign t[326] = t[380] ^ x[53];
  assign t[327] = t[381] ^ x[57];
  assign t[328] = t[382] ^ x[56];
  assign t[329] = t[383] ^ x[60];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[59];
  assign t[331] = t[385] ^ x[67];
  assign t[332] = t[386] ^ x[66];
  assign t[333] = t[387] ^ x[70];
  assign t[334] = t[388] ^ x[69];
  assign t[335] = t[389] ^ x[73];
  assign t[336] = t[390] ^ x[72];
  assign t[337] = t[391] ^ x[76];
  assign t[338] = t[392] ^ x[75];
  assign t[339] = t[393] ^ x[85];
  assign t[33] = t[51] ^ t[52];
  assign t[340] = t[394] ^ x[84];
  assign t[341] = t[395] ^ x[88];
  assign t[342] = t[396] ^ x[87];
  assign t[343] = t[397] ^ x[91];
  assign t[344] = t[398] ^ x[90];
  assign t[345] = t[399] ^ x[96];
  assign t[346] = t[400] ^ x[95];
  assign t[347] = (x[2]);
  assign t[348] = (x[2]);
  assign t[349] = (x[7]);
  assign t[34] = t[53] ^ t[54];
  assign t[350] = (x[7]);
  assign t[351] = (x[10]);
  assign t[352] = (x[10]);
  assign t[353] = (x[13]);
  assign t[354] = (x[13]);
  assign t[355] = (x[16]);
  assign t[356] = (x[16]);
  assign t[357] = (x[19]);
  assign t[358] = (x[19]);
  assign t[359] = (x[22]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[22]);
  assign t[361] = (x[25]);
  assign t[362] = (x[25]);
  assign t[363] = (x[28]);
  assign t[364] = (x[28]);
  assign t[365] = (x[31]);
  assign t[366] = (x[31]);
  assign t[367] = (x[34]);
  assign t[368] = (x[34]);
  assign t[369] = (x[37]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[37]);
  assign t[371] = (x[40]);
  assign t[372] = (x[40]);
  assign t[373] = (x[43]);
  assign t[374] = (x[43]);
  assign t[375] = (x[46]);
  assign t[376] = (x[46]);
  assign t[377] = (x[49]);
  assign t[378] = (x[49]);
  assign t[379] = (x[52]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[52]);
  assign t[381] = (x[55]);
  assign t[382] = (x[55]);
  assign t[383] = (x[58]);
  assign t[384] = (x[58]);
  assign t[385] = (x[65]);
  assign t[386] = (x[65]);
  assign t[387] = (x[68]);
  assign t[388] = (x[68]);
  assign t[389] = (x[71]);
  assign t[38] = ~(t[61] ^ t[62]);
  assign t[390] = (x[71]);
  assign t[391] = (x[74]);
  assign t[392] = (x[74]);
  assign t[393] = (x[83]);
  assign t[394] = (x[83]);
  assign t[395] = (x[86]);
  assign t[396] = (x[86]);
  assign t[397] = (x[89]);
  assign t[398] = (x[89]);
  assign t[399] = (x[94]);
  assign t[39] = ~(t[63] ^ t[64]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[94]);
  assign t[40] = t[65] ^ t[66];
  assign t[41] = t[67] ^ t[68];
  assign t[42] = t[69] ^ t[55];
  assign t[43] = ~(t[38] ^ t[70]);
  assign t[44] = t[11] ^ t[71];
  assign t[45] = ~(t[62] ^ t[41]);
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[216] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[217]);
  assign t[4] = t[8] ? t[9] : t[212];
  assign t[50] = ~(t[76] & t[218]);
  assign t[51] = t[77] ^ t[57];
  assign t[52] = t[78] & t[79];
  assign t[53] = t[80] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = t[84] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ? t[89] : t[219];
  assign t[58] = t[90] ^ t[91];
  assign t[59] = t[8] ? t[92] : t[220];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] ^ t[94];
  assign t[61] = ~(t[95] ^ t[96]);
  assign t[62] = t[97] ^ t[98];
  assign t[63] = t[99] ^ t[100];
  assign t[64] = ~(t[70] ^ t[41]);
  assign t[65] = t[101] ^ t[67];
  assign t[66] = t[102] ^ t[103];
  assign t[67] = t[104];
  assign t[68] = t[102] ^ t[87];
  assign t[69] = t[105] ^ t[106];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[107] ^ t[108];
  assign t[71] = t[109] ^ t[94];
  assign t[72] = ~(t[74] & t[110]);
  assign t[73] = ~(t[221] ^ t[111]);
  assign t[74] = ~(t[112] & t[113]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[222]);
  assign t[77] = t[88] ? t[114] : t[223];
  assign t[78] = ~(t[115]);
  assign t[79] = t[88] ? t[116] : t[224];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[117] : t[225];
  assign t[81] = t[215] ^ t[118];
  assign t[82] = ~(t[53] ^ t[119]);
  assign t[83] = t[97] ^ t[120];
  assign t[84] = t[121] ^ t[59];
  assign t[85] = t[93] ^ t[122];
  assign t[86] = t[123] ^ t[101];
  assign t[87] = t[124] & t[125];
  assign t[88] = ~(t[15]);
  assign t[89] = t[219] ^ t[126];
  assign t[8] = ~(t[15]);
  assign t[90] = t[127] ^ t[52];
  assign t[91] = t[128] & t[129];
  assign t[92] = t[220] ^ t[130];
  assign t[93] = t[131] ^ t[132];
  assign t[94] = t[133] & t[134];
  assign t[95] = t[40] ^ t[37];
  assign t[96] = t[135] ^ t[91];
  assign t[97] = t[81] ^ t[107];
  assign t[98] = t[119] ^ t[136];
  assign t[99] = t[137] ^ t[138];
  assign t[9] = t[212] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind141(x, y);
 input [116:0] x;
 output y;

 wire [400:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[139] ^ t[132];
  assign t[101] = ~t[140];
  assign t[102] = t[141] ^ t[106];
  assign t[103] = t[142] & t[143];
  assign t[104] = t[8] ? t[144] : t[226];
  assign t[105] = t[123] ^ t[67];
  assign t[106] = t[145] & t[146];
  assign t[107] = t[217] ^ t[147];
  assign t[108] = t[119] ^ t[54];
  assign t[109] = t[148] ^ t[121];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[149] & t[150]);
  assign t[111] = t[151] ^ t[227];
  assign t[112] = ~(t[221]);
  assign t[113] = t[152] & t[151];
  assign t[114] = t[223] ^ t[153];
  assign t[115] = t[88] ? t[154] : t[228];
  assign t[116] = t[224] ^ t[155];
  assign t[117] = t[225] ^ t[156];
  assign t[118] = t[8] ? t[157] : t[229];
  assign t[119] = t[158] ^ t[159];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[222] ^ t[160];
  assign t[121] = t[8] ? t[161] : t[230];
  assign t[122] = t[162] & t[163];
  assign t[123] = t[164];
  assign t[124] = ~(t[86] ^ t[102]);
  assign t[125] = t[65] ^ t[146];
  assign t[126] = t[165] ? x[62] : x[61];
  assign t[127] = t[166] & t[167];
  assign t[128] = ~(t[135] ^ t[90]);
  assign t[129] = t[137] ^ t[79];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[75] ? x[64] : x[63];
  assign t[131] = t[168] & t[169];
  assign t[132] = t[170] & t[171];
  assign t[133] = ~(t[109] ^ t[93]);
  assign t[134] = t[84] ^ t[171];
  assign t[135] = t[77] ^ t[115];
  assign t[136] = t[172] & t[173];
  assign t[137] = t[115] ^ t[57];
  assign t[138] = t[90] ^ t[174];
  assign t[139] = t[148] ^ t[59];
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[8] ? t[175] : t[231];
  assign t[141] = t[176] & t[177];
  assign t[142] = ~(t[141] ^ t[178]);
  assign t[143] = t[105] ^ t[179];
  assign t[144] = t[226] ^ t[180];
  assign t[145] = ~(t[101]);
  assign t[146] = t[181];
  assign t[147] = t[8] ? t[182] : t[232];
  assign t[148] = t[8] ? t[183] : t[233];
  assign t[149] = ~(t[152] | t[151]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[184] | t[112]);
  assign t[151] = ~(t[234]);
  assign t[152] = ~(t[227]);
  assign t[153] = t[165] ? x[78] : x[77];
  assign t[154] = t[228] ^ t[185];
  assign t[155] = t[165] ? x[80] : x[79];
  assign t[156] = t[28] ? x[82] : x[81];
  assign t[157] = t[229] ^ t[186];
  assign t[158] = t[187] & t[188];
  assign t[159] = t[189] & t[120];
  assign t[15] = ~(t[27]);
  assign t[160] = t[8] ? t[190] : t[235];
  assign t[161] = t[230] ^ t[191];
  assign t[162] = ~(t[131] ^ t[192]);
  assign t[163] = t[139] ^ t[193];
  assign t[164] = t[8] ? t[194] : t[236];
  assign t[165] = ~(t[48]);
  assign t[166] = ~(t[195]);
  assign t[167] = ~(t[77]);
  assign t[168] = ~(t[193]);
  assign t[169] = ~(t[148]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[121]);
  assign t[171] = t[8] ? t[196] : t[237];
  assign t[172] = ~(t[158] ^ t[197]);
  assign t[173] = t[198] ^ t[199];
  assign t[174] = t[200] & t[201];
  assign t[175] = t[231] ^ t[202];
  assign t[176] = ~(t[179]);
  assign t[177] = ~(t[123]);
  assign t[178] = t[65] ^ t[123];
  assign t[179] = t[146] ^ t[101];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[75] ? x[93] : x[92];
  assign t[181] = t[8] ? t[203] : t[238];
  assign t[182] = t[232] ^ t[204];
  assign t[183] = t[233] ^ t[205];
  assign t[184] = ~(t[216]);
  assign t[185] = t[165] ? x[98] : x[97];
  assign t[186] = t[28] ? x[100] : x[99];
  assign t[187] = ~(t[199]);
  assign t[188] = ~(t[80]);
  assign t[189] = ~(t[81]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[235] ^ t[206];
  assign t[191] = t[207] ? x[102] : x[101];
  assign t[192] = t[84] ^ t[148];
  assign t[193] = t[171] ^ t[121];
  assign t[194] = t[236] ^ t[208];
  assign t[195] = t[79] ^ t[115];
  assign t[196] = t[237] ^ t[209];
  assign t[197] = t[97] ^ t[80];
  assign t[198] = t[80] ^ t[107];
  assign t[199] = t[120] ^ t[81];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[127] ^ t[210]);
  assign t[201] = t[51] ^ t[195];
  assign t[202] = t[28] ? x[104] : x[103];
  assign t[203] = t[238] ^ t[211];
  assign t[204] = t[28] ? x[106] : x[105];
  assign t[205] = t[207] ? x[108] : x[107];
  assign t[206] = t[28] ? x[110] : x[109];
  assign t[207] = ~(t[48]);
  assign t[208] = t[75] ? x[112] : x[111];
  assign t[209] = t[207] ? x[114] : x[113];
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = t[137] ^ t[77];
  assign t[211] = t[75] ? x[116] : x[115];
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[35]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[38] ^ t[39];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = t[266] ^ x[4];
  assign t[23] = t[22] ^ t[34];
  assign t[240] = t[267] ^ x[9];
  assign t[241] = t[268] ^ x[12];
  assign t[242] = t[269] ^ x[15];
  assign t[243] = t[270] ^ x[18];
  assign t[244] = t[271] ^ x[21];
  assign t[245] = t[272] ^ x[24];
  assign t[246] = t[273] ^ x[27];
  assign t[247] = t[274] ^ x[30];
  assign t[248] = t[275] ^ x[33];
  assign t[249] = t[276] ^ x[36];
  assign t[24] = ~(t[40] ^ t[41]);
  assign t[250] = t[277] ^ x[39];
  assign t[251] = t[278] ^ x[42];
  assign t[252] = t[279] ^ x[45];
  assign t[253] = t[280] ^ x[48];
  assign t[254] = t[281] ^ x[51];
  assign t[255] = t[282] ^ x[54];
  assign t[256] = t[283] ^ x[57];
  assign t[257] = t[284] ^ x[60];
  assign t[258] = t[285] ^ x[67];
  assign t[259] = t[286] ^ x[70];
  assign t[25] = ~(t[42] ^ t[43]);
  assign t[260] = t[287] ^ x[73];
  assign t[261] = t[288] ^ x[76];
  assign t[262] = t[289] ^ x[85];
  assign t[263] = t[290] ^ x[88];
  assign t[264] = t[291] ^ x[91];
  assign t[265] = t[292] ^ x[96];
  assign t[266] = (t[293] & ~t[294]);
  assign t[267] = (t[295] & ~t[296]);
  assign t[268] = (t[297] & ~t[298]);
  assign t[269] = (t[299] & ~t[300]);
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[270] = (t[301] & ~t[302]);
  assign t[271] = (t[303] & ~t[304]);
  assign t[272] = (t[305] & ~t[306]);
  assign t[273] = (t[307] & ~t[308]);
  assign t[274] = (t[309] & ~t[310]);
  assign t[275] = (t[311] & ~t[312]);
  assign t[276] = (t[313] & ~t[314]);
  assign t[277] = (t[315] & ~t[316]);
  assign t[278] = (t[317] & ~t[318]);
  assign t[279] = (t[319] & ~t[320]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = t[347] ^ x[4];
  assign t[294] = t[348] ^ x[3];
  assign t[295] = t[349] ^ x[9];
  assign t[296] = t[350] ^ x[8];
  assign t[297] = t[351] ^ x[12];
  assign t[298] = t[352] ^ x[11];
  assign t[299] = t[353] ^ x[15];
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[14];
  assign t[301] = t[355] ^ x[18];
  assign t[302] = t[356] ^ x[17];
  assign t[303] = t[357] ^ x[21];
  assign t[304] = t[358] ^ x[20];
  assign t[305] = t[359] ^ x[24];
  assign t[306] = t[360] ^ x[23];
  assign t[307] = t[361] ^ x[27];
  assign t[308] = t[362] ^ x[26];
  assign t[309] = t[363] ^ x[30];
  assign t[30] = ~(t[214]);
  assign t[310] = t[364] ^ x[29];
  assign t[311] = t[365] ^ x[33];
  assign t[312] = t[366] ^ x[32];
  assign t[313] = t[367] ^ x[36];
  assign t[314] = t[368] ^ x[35];
  assign t[315] = t[369] ^ x[39];
  assign t[316] = t[370] ^ x[38];
  assign t[317] = t[371] ^ x[42];
  assign t[318] = t[372] ^ x[41];
  assign t[319] = t[373] ^ x[45];
  assign t[31] = ~(t[215]);
  assign t[320] = t[374] ^ x[44];
  assign t[321] = t[375] ^ x[48];
  assign t[322] = t[376] ^ x[47];
  assign t[323] = t[377] ^ x[51];
  assign t[324] = t[378] ^ x[50];
  assign t[325] = t[379] ^ x[54];
  assign t[326] = t[380] ^ x[53];
  assign t[327] = t[381] ^ x[57];
  assign t[328] = t[382] ^ x[56];
  assign t[329] = t[383] ^ x[60];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[59];
  assign t[331] = t[385] ^ x[67];
  assign t[332] = t[386] ^ x[66];
  assign t[333] = t[387] ^ x[70];
  assign t[334] = t[388] ^ x[69];
  assign t[335] = t[389] ^ x[73];
  assign t[336] = t[390] ^ x[72];
  assign t[337] = t[391] ^ x[76];
  assign t[338] = t[392] ^ x[75];
  assign t[339] = t[393] ^ x[85];
  assign t[33] = t[51] ^ t[52];
  assign t[340] = t[394] ^ x[84];
  assign t[341] = t[395] ^ x[88];
  assign t[342] = t[396] ^ x[87];
  assign t[343] = t[397] ^ x[91];
  assign t[344] = t[398] ^ x[90];
  assign t[345] = t[399] ^ x[96];
  assign t[346] = t[400] ^ x[95];
  assign t[347] = (x[2]);
  assign t[348] = (x[2]);
  assign t[349] = (x[7]);
  assign t[34] = t[53] ^ t[54];
  assign t[350] = (x[7]);
  assign t[351] = (x[10]);
  assign t[352] = (x[10]);
  assign t[353] = (x[13]);
  assign t[354] = (x[13]);
  assign t[355] = (x[16]);
  assign t[356] = (x[16]);
  assign t[357] = (x[19]);
  assign t[358] = (x[19]);
  assign t[359] = (x[22]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[22]);
  assign t[361] = (x[25]);
  assign t[362] = (x[25]);
  assign t[363] = (x[28]);
  assign t[364] = (x[28]);
  assign t[365] = (x[31]);
  assign t[366] = (x[31]);
  assign t[367] = (x[34]);
  assign t[368] = (x[34]);
  assign t[369] = (x[37]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[37]);
  assign t[371] = (x[40]);
  assign t[372] = (x[40]);
  assign t[373] = (x[43]);
  assign t[374] = (x[43]);
  assign t[375] = (x[46]);
  assign t[376] = (x[46]);
  assign t[377] = (x[49]);
  assign t[378] = (x[49]);
  assign t[379] = (x[52]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[52]);
  assign t[381] = (x[55]);
  assign t[382] = (x[55]);
  assign t[383] = (x[58]);
  assign t[384] = (x[58]);
  assign t[385] = (x[65]);
  assign t[386] = (x[65]);
  assign t[387] = (x[68]);
  assign t[388] = (x[68]);
  assign t[389] = (x[71]);
  assign t[38] = ~(t[61] ^ t[62]);
  assign t[390] = (x[71]);
  assign t[391] = (x[74]);
  assign t[392] = (x[74]);
  assign t[393] = (x[83]);
  assign t[394] = (x[83]);
  assign t[395] = (x[86]);
  assign t[396] = (x[86]);
  assign t[397] = (x[89]);
  assign t[398] = (x[89]);
  assign t[399] = (x[94]);
  assign t[39] = ~(t[63] ^ t[64]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[94]);
  assign t[40] = t[65] ^ t[66];
  assign t[41] = t[67] ^ t[68];
  assign t[42] = t[69] ^ t[55];
  assign t[43] = ~(t[38] ^ t[70]);
  assign t[44] = t[11] ^ t[71];
  assign t[45] = ~(t[62] ^ t[41]);
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[216] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[217]);
  assign t[4] = t[8] ? t[9] : t[212];
  assign t[50] = ~(t[76] & t[218]);
  assign t[51] = t[77] ^ t[57];
  assign t[52] = t[78] & t[79];
  assign t[53] = t[80] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = t[84] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ? t[89] : t[219];
  assign t[58] = t[90] ^ t[91];
  assign t[59] = t[8] ? t[92] : t[220];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] ^ t[94];
  assign t[61] = ~(t[95] ^ t[96]);
  assign t[62] = t[97] ^ t[98];
  assign t[63] = t[99] ^ t[100];
  assign t[64] = ~(t[70] ^ t[41]);
  assign t[65] = t[101] ^ t[67];
  assign t[66] = t[102] ^ t[103];
  assign t[67] = t[104];
  assign t[68] = t[102] ^ t[87];
  assign t[69] = t[105] ^ t[106];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[107] ^ t[108];
  assign t[71] = t[109] ^ t[94];
  assign t[72] = ~(t[74] & t[110]);
  assign t[73] = ~(t[221] ^ t[111]);
  assign t[74] = ~(t[112] & t[113]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[222]);
  assign t[77] = t[88] ? t[114] : t[223];
  assign t[78] = ~(t[115]);
  assign t[79] = t[88] ? t[116] : t[224];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[117] : t[225];
  assign t[81] = t[215] ^ t[118];
  assign t[82] = ~(t[53] ^ t[119]);
  assign t[83] = t[97] ^ t[120];
  assign t[84] = t[121] ^ t[59];
  assign t[85] = t[93] ^ t[122];
  assign t[86] = t[123] ^ t[101];
  assign t[87] = t[124] & t[125];
  assign t[88] = ~(t[15]);
  assign t[89] = t[219] ^ t[126];
  assign t[8] = ~(t[15]);
  assign t[90] = t[127] ^ t[52];
  assign t[91] = t[128] & t[129];
  assign t[92] = t[220] ^ t[130];
  assign t[93] = t[131] ^ t[132];
  assign t[94] = t[133] & t[134];
  assign t[95] = t[40] ^ t[37];
  assign t[96] = t[135] ^ t[91];
  assign t[97] = t[81] ^ t[107];
  assign t[98] = t[119] ^ t[136];
  assign t[99] = t[137] ^ t[138];
  assign t[9] = t[212] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[141] ^ t[142];
  assign t[101] = t[28] ? x[56] : x[55];
  assign t[102] = t[218] ^ t[143];
  assign t[103] = t[8] ? t[144] : t[227];
  assign t[104] = ~(t[145] & t[146]);
  assign t[105] = t[147] ^ t[228];
  assign t[106] = ~(t[220]);
  assign t[107] = t[148] & t[147];
  assign t[108] = t[87] ^ t[127];
  assign t[109] = t[149] & t[150];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[132] ? t[151] : t[229];
  assign t[111] = t[112] ^ t[62];
  assign t[112] = t[152] ^ t[153];
  assign t[113] = t[154] & t[155];
  assign t[114] = t[221] ^ t[156];
  assign t[115] = t[157] ^ t[59];
  assign t[116] = t[127] ^ t[78];
  assign t[117] = t[115] ^ t[158];
  assign t[118] = t[159] ^ t[129];
  assign t[119] = t[160] & t[161];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[63] ^ t[162];
  assign t[121] = t[141] ^ t[98];
  assign t[122] = t[159] ^ t[124];
  assign t[123] = t[163] & t[164];
  assign t[124] = t[165];
  assign t[125] = t[130] ^ t[119];
  assign t[126] = t[222] ^ t[166];
  assign t[127] = t[8] ? t[167] : t[230];
  assign t[128] = t[223] ^ t[168];
  assign t[129] = ~t[169];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[170] ^ t[123];
  assign t[131] = t[171] & t[172];
  assign t[132] = ~(t[15]);
  assign t[133] = t[224] ^ t[173];
  assign t[134] = t[225] ^ t[174];
  assign t[135] = t[132] ? t[175] : t[231];
  assign t[136] = t[226] ^ t[176];
  assign t[137] = ~(t[142]);
  assign t[138] = ~(t[42]);
  assign t[139] = ~(t[43]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[40] ^ t[42];
  assign t[141] = t[42] ^ t[63];
  assign t[142] = t[68] ^ t[43];
  assign t[143] = t[28] ? x[73] : x[72];
  assign t[144] = t[227] ^ t[177];
  assign t[145] = ~(t[148] | t[147]);
  assign t[146] = ~(t[178] | t[106]);
  assign t[147] = ~(t[232]);
  assign t[148] = ~(t[228]);
  assign t[149] = ~(t[108] ^ t[115]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[116] ^ t[89];
  assign t[151] = t[229] ^ t[179];
  assign t[152] = t[180] & t[181];
  assign t[153] = t[182] & t[135];
  assign t[154] = ~(t[152] ^ t[183]);
  assign t[155] = t[184] ^ t[185];
  assign t[156] = t[72] ? x[78] : x[77];
  assign t[157] = t[186] & t[187];
  assign t[158] = t[188] & t[189];
  assign t[159] = t[190];
  assign t[15] = ~(t[27]);
  assign t[160] = ~(t[118] ^ t[130]);
  assign t[161] = t[90] ^ t[164];
  assign t[162] = t[64] ^ t[26];
  assign t[163] = ~(t[129]);
  assign t[164] = t[191];
  assign t[165] = t[8] ? t[192] : t[233];
  assign t[166] = t[193] ? x[83] : x[82];
  assign t[167] = t[230] ^ t[194];
  assign t[168] = t[193] ? x[85] : x[84];
  assign t[169] = t[8] ? t[195] : t[234];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[196] & t[197];
  assign t[171] = ~(t[170] ^ t[198]);
  assign t[172] = t[122] ^ t[199];
  assign t[173] = t[200] ? x[90] : x[89];
  assign t[174] = t[200] ? x[92] : x[91];
  assign t[175] = t[231] ^ t[201];
  assign t[176] = t[28] ? x[94] : x[93];
  assign t[177] = t[28] ? x[96] : x[95];
  assign t[178] = ~(t[215]);
  assign t[179] = t[200] ? x[98] : x[97];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[185]);
  assign t[181] = ~(t[92]);
  assign t[182] = ~(t[93]);
  assign t[183] = t[76] ^ t[92];
  assign t[184] = t[92] ^ t[110];
  assign t[185] = t[135] ^ t[93];
  assign t[186] = ~(t[202]);
  assign t[187] = ~(t[87]);
  assign t[188] = ~(t[157] ^ t[203]);
  assign t[189] = t[58] ^ t[202];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[8] ? t[204] : t[235];
  assign t[191] = t[8] ? t[205] : t[236];
  assign t[192] = t[233] ^ t[206];
  assign t[193] = ~(t[48]);
  assign t[194] = t[193] ? x[106] : x[105];
  assign t[195] = t[234] ^ t[207];
  assign t[196] = ~(t[199]);
  assign t[197] = ~(t[159]);
  assign t[198] = t[90] ^ t[159];
  assign t[199] = t[164] ^ t[129];
  assign t[19] = ~(t[24] ^ t[33]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[48]);
  assign t[201] = t[200] ? x[108] : x[107];
  assign t[202] = t[89] ^ t[127];
  assign t[203] = t[116] ^ t[87];
  assign t[204] = t[235] ^ t[208];
  assign t[205] = t[236] ^ t[209];
  assign t[206] = t[72] ? x[110] : x[109];
  assign t[207] = t[28] ? x[112] : x[111];
  assign t[208] = t[72] ? x[114] : x[113];
  assign t[209] = t[72] ? x[116] : x[115];
  assign t[20] = ~(t[34] ^ t[35]);
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[38] ^ t[14]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[9];
  assign t[239] = t[266] ^ x[12];
  assign t[23] = ~(t[38] ^ t[39]);
  assign t[240] = t[267] ^ x[15];
  assign t[241] = t[268] ^ x[18];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = t[40] ^ t[41];
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[51];
  assign t[253] = t[280] ^ x[54];
  assign t[254] = t[281] ^ x[59];
  assign t[255] = t[282] ^ x[62];
  assign t[256] = t[283] ^ x[65];
  assign t[257] = t[284] ^ x[68];
  assign t[258] = t[285] ^ x[71];
  assign t[259] = t[286] ^ x[76];
  assign t[25] = t[42] ^ t[43];
  assign t[260] = t[287] ^ x[81];
  assign t[261] = t[288] ^ x[88];
  assign t[262] = t[289] ^ x[101];
  assign t[263] = t[290] ^ x[104];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = t[44] & t[45];
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[9];
  assign t[294] = t[348] ^ x[8];
  assign t[295] = t[349] ^ x[12];
  assign t[296] = t[350] ^ x[11];
  assign t[297] = t[351] ^ x[15];
  assign t[298] = t[352] ^ x[14];
  assign t[299] = t[353] ^ x[18];
  assign t[29] = ~(t[211]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[17];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = ~(t[212]);
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[213]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[51];
  assign t[322] = t[376] ^ x[50];
  assign t[323] = t[377] ^ x[54];
  assign t[324] = t[378] ^ x[53];
  assign t[325] = t[379] ^ x[59];
  assign t[326] = t[380] ^ x[58];
  assign t[327] = t[381] ^ x[62];
  assign t[328] = t[382] ^ x[61];
  assign t[329] = t[383] ^ x[65];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[64];
  assign t[331] = t[385] ^ x[68];
  assign t[332] = t[386] ^ x[67];
  assign t[333] = t[387] ^ x[71];
  assign t[334] = t[388] ^ x[70];
  assign t[335] = t[389] ^ x[76];
  assign t[336] = t[390] ^ x[75];
  assign t[337] = t[391] ^ x[81];
  assign t[338] = t[392] ^ x[80];
  assign t[339] = t[393] ^ x[88];
  assign t[33] = ~(t[51] ^ t[52]);
  assign t[340] = t[394] ^ x[87];
  assign t[341] = t[395] ^ x[101];
  assign t[342] = t[396] ^ x[100];
  assign t[343] = t[397] ^ x[104];
  assign t[344] = t[398] ^ x[103];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[7]);
  assign t[348] = (x[7]);
  assign t[349] = (x[10]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[10]);
  assign t[351] = (x[13]);
  assign t[352] = (x[13]);
  assign t[353] = (x[16]);
  assign t[354] = (x[16]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = t[13] ^ t[55];
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[49]);
  assign t[376] = (x[49]);
  assign t[377] = (x[52]);
  assign t[378] = (x[52]);
  assign t[379] = (x[57]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[57]);
  assign t[381] = (x[60]);
  assign t[382] = (x[60]);
  assign t[383] = (x[63]);
  assign t[384] = (x[63]);
  assign t[385] = (x[66]);
  assign t[386] = (x[66]);
  assign t[387] = (x[69]);
  assign t[388] = (x[69]);
  assign t[389] = (x[74]);
  assign t[38] = t[60] ^ t[53];
  assign t[390] = (x[74]);
  assign t[391] = (x[79]);
  assign t[392] = (x[79]);
  assign t[393] = (x[86]);
  assign t[394] = (x[86]);
  assign t[395] = (x[99]);
  assign t[396] = (x[99]);
  assign t[397] = (x[102]);
  assign t[398] = (x[102]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[43] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[8] ? t[66] : t[214];
  assign t[43] = t[213] ^ t[67];
  assign t[44] = ~(t[25] ^ t[64]);
  assign t[45] = t[40] ^ t[68];
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = t[215] | t[71];
  assign t[48] = ~(t[72]);
  assign t[49] = ~(t[216]);
  assign t[4] = t[8] ? t[9] : t[210];
  assign t[50] = ~(t[73] & t[217]);
  assign t[51] = ~(t[74] ^ t[75]);
  assign t[52] = t[76] ^ t[77];
  assign t[53] = t[78] ^ t[79];
  assign t[54] = t[80] ^ t[81];
  assign t[55] = ~(t[82] ^ t[83]);
  assign t[56] = t[84] ^ t[33];
  assign t[57] = ~(t[85] ^ t[86]);
  assign t[58] = t[87] ^ t[78];
  assign t[59] = t[88] & t[89];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92] ^ t[93];
  assign t[62] = t[94] & t[95];
  assign t[63] = t[216] ^ t[96];
  assign t[64] = t[97] ^ t[98];
  assign t[65] = t[99] & t[100];
  assign t[66] = t[214] ^ t[101];
  assign t[67] = t[8] ? t[102] : t[218];
  assign t[68] = t[219] ^ t[103];
  assign t[69] = ~(t[71] & t[104]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[220] ^ t[105]);
  assign t[71] = ~(t[106] & t[107]);
  assign t[72] = ~(t[47]);
  assign t[73] = ~(t[219]);
  assign t[74] = t[108] ^ t[109];
  assign t[75] = t[110] ^ t[111];
  assign t[76] = t[93] ^ t[110];
  assign t[77] = t[112] ^ t[113];
  assign t[78] = t[8] ? t[114] : t[221];
  assign t[79] = t[115] ^ t[109];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[116] ^ t[117];
  assign t[81] = t[118] ^ t[119];
  assign t[82] = t[52] ^ t[37];
  assign t[83] = ~(t[120] ^ t[86]);
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[122] ^ t[123];
  assign t[86] = t[124] ^ t[125];
  assign t[87] = t[8] ? t[126] : t[222];
  assign t[88] = ~(t[127]);
  assign t[89] = t[8] ? t[128] : t[223];
  assign t[8] = ~(t[15]);
  assign t[90] = t[129] ^ t[124];
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[132] ? t[133] : t[224];
  assign t[93] = t[132] ? t[134] : t[225];
  assign t[94] = ~(t[61] ^ t[112]);
  assign t[95] = t[76] ^ t[135];
  assign t[96] = t[8] ? t[136] : t[226];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[139] & t[68];
  assign t[99] = ~(t[97] ^ t[140]);
  assign t[9] = t[210] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[141] ^ t[142];
  assign t[101] = t[28] ? x[56] : x[55];
  assign t[102] = t[218] ^ t[143];
  assign t[103] = t[8] ? t[144] : t[227];
  assign t[104] = ~(t[145] & t[146]);
  assign t[105] = t[147] ^ t[228];
  assign t[106] = ~(t[220]);
  assign t[107] = t[148] & t[147];
  assign t[108] = t[87] ^ t[127];
  assign t[109] = t[149] & t[150];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[132] ? t[151] : t[229];
  assign t[111] = t[112] ^ t[62];
  assign t[112] = t[152] ^ t[153];
  assign t[113] = t[154] & t[155];
  assign t[114] = t[221] ^ t[156];
  assign t[115] = t[157] ^ t[59];
  assign t[116] = t[127] ^ t[78];
  assign t[117] = t[115] ^ t[158];
  assign t[118] = t[159] ^ t[129];
  assign t[119] = t[160] & t[161];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[63] ^ t[162];
  assign t[121] = t[141] ^ t[98];
  assign t[122] = t[159] ^ t[124];
  assign t[123] = t[163] & t[164];
  assign t[124] = t[165];
  assign t[125] = t[130] ^ t[119];
  assign t[126] = t[222] ^ t[166];
  assign t[127] = t[8] ? t[167] : t[230];
  assign t[128] = t[223] ^ t[168];
  assign t[129] = ~t[169];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[170] ^ t[123];
  assign t[131] = t[171] & t[172];
  assign t[132] = ~(t[15]);
  assign t[133] = t[224] ^ t[173];
  assign t[134] = t[225] ^ t[174];
  assign t[135] = t[132] ? t[175] : t[231];
  assign t[136] = t[226] ^ t[176];
  assign t[137] = ~(t[142]);
  assign t[138] = ~(t[42]);
  assign t[139] = ~(t[43]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[40] ^ t[42];
  assign t[141] = t[42] ^ t[63];
  assign t[142] = t[68] ^ t[43];
  assign t[143] = t[28] ? x[73] : x[72];
  assign t[144] = t[227] ^ t[177];
  assign t[145] = ~(t[148] | t[147]);
  assign t[146] = ~(t[178] | t[106]);
  assign t[147] = ~(t[232]);
  assign t[148] = ~(t[228]);
  assign t[149] = ~(t[108] ^ t[115]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[116] ^ t[89];
  assign t[151] = t[229] ^ t[179];
  assign t[152] = t[180] & t[181];
  assign t[153] = t[182] & t[135];
  assign t[154] = ~(t[152] ^ t[183]);
  assign t[155] = t[184] ^ t[185];
  assign t[156] = t[72] ? x[78] : x[77];
  assign t[157] = t[186] & t[187];
  assign t[158] = t[188] & t[189];
  assign t[159] = t[190];
  assign t[15] = ~(t[27]);
  assign t[160] = ~(t[118] ^ t[130]);
  assign t[161] = t[90] ^ t[164];
  assign t[162] = t[64] ^ t[26];
  assign t[163] = ~(t[129]);
  assign t[164] = t[191];
  assign t[165] = t[8] ? t[192] : t[233];
  assign t[166] = t[193] ? x[83] : x[82];
  assign t[167] = t[230] ^ t[194];
  assign t[168] = t[193] ? x[85] : x[84];
  assign t[169] = t[8] ? t[195] : t[234];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[196] & t[197];
  assign t[171] = ~(t[170] ^ t[198]);
  assign t[172] = t[122] ^ t[199];
  assign t[173] = t[200] ? x[90] : x[89];
  assign t[174] = t[200] ? x[92] : x[91];
  assign t[175] = t[231] ^ t[201];
  assign t[176] = t[28] ? x[94] : x[93];
  assign t[177] = t[28] ? x[96] : x[95];
  assign t[178] = ~(t[215]);
  assign t[179] = t[200] ? x[98] : x[97];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[185]);
  assign t[181] = ~(t[92]);
  assign t[182] = ~(t[93]);
  assign t[183] = t[76] ^ t[92];
  assign t[184] = t[92] ^ t[110];
  assign t[185] = t[135] ^ t[93];
  assign t[186] = ~(t[202]);
  assign t[187] = ~(t[87]);
  assign t[188] = ~(t[157] ^ t[203]);
  assign t[189] = t[58] ^ t[202];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[8] ? t[204] : t[235];
  assign t[191] = t[8] ? t[205] : t[236];
  assign t[192] = t[233] ^ t[206];
  assign t[193] = ~(t[48]);
  assign t[194] = t[193] ? x[106] : x[105];
  assign t[195] = t[234] ^ t[207];
  assign t[196] = ~(t[199]);
  assign t[197] = ~(t[159]);
  assign t[198] = t[90] ^ t[159];
  assign t[199] = t[164] ^ t[129];
  assign t[19] = ~(t[24] ^ t[33]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[48]);
  assign t[201] = t[200] ? x[108] : x[107];
  assign t[202] = t[89] ^ t[127];
  assign t[203] = t[116] ^ t[87];
  assign t[204] = t[235] ^ t[208];
  assign t[205] = t[236] ^ t[209];
  assign t[206] = t[72] ? x[110] : x[109];
  assign t[207] = t[28] ? x[112] : x[111];
  assign t[208] = t[72] ? x[114] : x[113];
  assign t[209] = t[72] ? x[116] : x[115];
  assign t[20] = ~(t[34] ^ t[35]);
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[38] ^ t[14]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[9];
  assign t[239] = t[266] ^ x[12];
  assign t[23] = ~(t[38] ^ t[39]);
  assign t[240] = t[267] ^ x[15];
  assign t[241] = t[268] ^ x[18];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = t[40] ^ t[41];
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[51];
  assign t[253] = t[280] ^ x[54];
  assign t[254] = t[281] ^ x[59];
  assign t[255] = t[282] ^ x[62];
  assign t[256] = t[283] ^ x[65];
  assign t[257] = t[284] ^ x[68];
  assign t[258] = t[285] ^ x[71];
  assign t[259] = t[286] ^ x[76];
  assign t[25] = t[42] ^ t[43];
  assign t[260] = t[287] ^ x[81];
  assign t[261] = t[288] ^ x[88];
  assign t[262] = t[289] ^ x[101];
  assign t[263] = t[290] ^ x[104];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = t[44] & t[45];
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[9];
  assign t[294] = t[348] ^ x[8];
  assign t[295] = t[349] ^ x[12];
  assign t[296] = t[350] ^ x[11];
  assign t[297] = t[351] ^ x[15];
  assign t[298] = t[352] ^ x[14];
  assign t[299] = t[353] ^ x[18];
  assign t[29] = ~(t[211]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[17];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = ~(t[212]);
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[213]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[51];
  assign t[322] = t[376] ^ x[50];
  assign t[323] = t[377] ^ x[54];
  assign t[324] = t[378] ^ x[53];
  assign t[325] = t[379] ^ x[59];
  assign t[326] = t[380] ^ x[58];
  assign t[327] = t[381] ^ x[62];
  assign t[328] = t[382] ^ x[61];
  assign t[329] = t[383] ^ x[65];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[64];
  assign t[331] = t[385] ^ x[68];
  assign t[332] = t[386] ^ x[67];
  assign t[333] = t[387] ^ x[71];
  assign t[334] = t[388] ^ x[70];
  assign t[335] = t[389] ^ x[76];
  assign t[336] = t[390] ^ x[75];
  assign t[337] = t[391] ^ x[81];
  assign t[338] = t[392] ^ x[80];
  assign t[339] = t[393] ^ x[88];
  assign t[33] = ~(t[51] ^ t[52]);
  assign t[340] = t[394] ^ x[87];
  assign t[341] = t[395] ^ x[101];
  assign t[342] = t[396] ^ x[100];
  assign t[343] = t[397] ^ x[104];
  assign t[344] = t[398] ^ x[103];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[7]);
  assign t[348] = (x[7]);
  assign t[349] = (x[10]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[10]);
  assign t[351] = (x[13]);
  assign t[352] = (x[13]);
  assign t[353] = (x[16]);
  assign t[354] = (x[16]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = t[13] ^ t[55];
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[49]);
  assign t[376] = (x[49]);
  assign t[377] = (x[52]);
  assign t[378] = (x[52]);
  assign t[379] = (x[57]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[57]);
  assign t[381] = (x[60]);
  assign t[382] = (x[60]);
  assign t[383] = (x[63]);
  assign t[384] = (x[63]);
  assign t[385] = (x[66]);
  assign t[386] = (x[66]);
  assign t[387] = (x[69]);
  assign t[388] = (x[69]);
  assign t[389] = (x[74]);
  assign t[38] = t[60] ^ t[53];
  assign t[390] = (x[74]);
  assign t[391] = (x[79]);
  assign t[392] = (x[79]);
  assign t[393] = (x[86]);
  assign t[394] = (x[86]);
  assign t[395] = (x[99]);
  assign t[396] = (x[99]);
  assign t[397] = (x[102]);
  assign t[398] = (x[102]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[43] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[8] ? t[66] : t[214];
  assign t[43] = t[213] ^ t[67];
  assign t[44] = ~(t[25] ^ t[64]);
  assign t[45] = t[40] ^ t[68];
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = t[215] | t[71];
  assign t[48] = ~(t[72]);
  assign t[49] = ~(t[216]);
  assign t[4] = t[8] ? t[9] : t[210];
  assign t[50] = ~(t[73] & t[217]);
  assign t[51] = ~(t[74] ^ t[75]);
  assign t[52] = t[76] ^ t[77];
  assign t[53] = t[78] ^ t[79];
  assign t[54] = t[80] ^ t[81];
  assign t[55] = ~(t[82] ^ t[83]);
  assign t[56] = t[84] ^ t[33];
  assign t[57] = ~(t[85] ^ t[86]);
  assign t[58] = t[87] ^ t[78];
  assign t[59] = t[88] & t[89];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92] ^ t[93];
  assign t[62] = t[94] & t[95];
  assign t[63] = t[216] ^ t[96];
  assign t[64] = t[97] ^ t[98];
  assign t[65] = t[99] & t[100];
  assign t[66] = t[214] ^ t[101];
  assign t[67] = t[8] ? t[102] : t[218];
  assign t[68] = t[219] ^ t[103];
  assign t[69] = ~(t[71] & t[104]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[220] ^ t[105]);
  assign t[71] = ~(t[106] & t[107]);
  assign t[72] = ~(t[47]);
  assign t[73] = ~(t[219]);
  assign t[74] = t[108] ^ t[109];
  assign t[75] = t[110] ^ t[111];
  assign t[76] = t[93] ^ t[110];
  assign t[77] = t[112] ^ t[113];
  assign t[78] = t[8] ? t[114] : t[221];
  assign t[79] = t[115] ^ t[109];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[116] ^ t[117];
  assign t[81] = t[118] ^ t[119];
  assign t[82] = t[52] ^ t[37];
  assign t[83] = ~(t[120] ^ t[86]);
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[122] ^ t[123];
  assign t[86] = t[124] ^ t[125];
  assign t[87] = t[8] ? t[126] : t[222];
  assign t[88] = ~(t[127]);
  assign t[89] = t[8] ? t[128] : t[223];
  assign t[8] = ~(t[15]);
  assign t[90] = t[129] ^ t[124];
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[132] ? t[133] : t[224];
  assign t[93] = t[132] ? t[134] : t[225];
  assign t[94] = ~(t[61] ^ t[112]);
  assign t[95] = t[76] ^ t[135];
  assign t[96] = t[8] ? t[136] : t[226];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[139] & t[68];
  assign t[99] = ~(t[97] ^ t[140]);
  assign t[9] = t[210] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [116:0] x;
 output y;

 wire [400:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[116] ^ t[142];
  assign t[101] = t[27] ? t[143] : t[226];
  assign t[102] = t[27] ? t[144] : t[227];
  assign t[103] = t[27] ? t[145] : t[228];
  assign t[104] = t[28] ? x[56] : x[55];
  assign t[105] = ~(t[117] ^ t[57]);
  assign t[106] = t[35] ^ t[127];
  assign t[107] = t[223] ^ t[146];
  assign t[108] = t[147] & t[148];
  assign t[109] = t[149] & t[150];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[93] ^ t[72]);
  assign t[111] = t[151] ^ t[150];
  assign t[112] = ~(t[152] & t[153]);
  assign t[113] = t[154] ^ t[229];
  assign t[114] = ~(t[224]);
  assign t[115] = t[155] & t[154];
  assign t[116] = t[156] ^ t[62];
  assign t[117] = t[157] ^ t[56];
  assign t[118] = t[122] ^ t[158];
  assign t[119] = t[63] ^ t[159];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[27] ? t[160] : t[230];
  assign t[121] = t[161] ^ t[42];
  assign t[122] = t[83] ^ t[66];
  assign t[123] = t[28] ? x[64] : x[63];
  assign t[124] = ~(t[130]);
  assign t[125] = ~(t[157]);
  assign t[126] = ~(t[56]);
  assign t[127] = t[8] ? t[162] : t[231];
  assign t[128] = t[35] ^ t[157];
  assign t[129] = t[157] ^ t[43];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[127] ^ t[56];
  assign t[131] = ~(t[163] ^ t[164]);
  assign t[132] = t[165] ^ t[166];
  assign t[133] = t[8] ? t[167] : t[232];
  assign t[134] = t[213] ^ t[168];
  assign t[135] = t[169] ? x[72] : x[71];
  assign t[136] = t[169] ? x[74] : x[73];
  assign t[137] = ~(t[142]);
  assign t[138] = ~(t[156]);
  assign t[139] = ~(t[61]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[94] ? t[170] : t[233];
  assign t[141] = t[39] ^ t[156];
  assign t[142] = t[140] ^ t[61];
  assign t[143] = t[226] ^ t[171];
  assign t[144] = t[227] ^ t[172];
  assign t[145] = t[228] ^ t[173];
  assign t[146] = t[77] ? x[79] : x[78];
  assign t[147] = ~(t[174]);
  assign t[148] = ~(t[133]);
  assign t[149] = ~(t[134]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[214] ^ t[175];
  assign t[151] = t[134] ^ t[45];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[176] | t[114]);
  assign t[154] = ~(t[234]);
  assign t[155] = ~(t[229]);
  assign t[156] = t[94] ? t[177] : t[235];
  assign t[157] = t[8] ? t[178] : t[236];
  assign t[158] = t[121] ^ t[179];
  assign t[159] = t[180] & t[181];
  assign t[15] = ~(t[27]);
  assign t[160] = t[230] ^ t[182];
  assign t[161] = t[183] & t[184];
  assign t[162] = t[231] ^ t[185];
  assign t[163] = t[186] ^ t[187];
  assign t[164] = ~(t[188] ^ t[26]);
  assign t[165] = t[151] ^ t[189];
  assign t[166] = t[66] ^ t[190];
  assign t[167] = t[232] ^ t[191];
  assign t[168] = t[27] ? t[192] : t[237];
  assign t[169] = ~(t[49]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[233] ^ t[193];
  assign t[171] = t[77] ? x[93] : x[92];
  assign t[172] = t[77] ? x[95] : x[94];
  assign t[173] = t[28] ? x[97] : x[96];
  assign t[174] = t[150] ^ t[134];
  assign t[175] = t[8] ? t[194] : t[238];
  assign t[176] = ~(t[218]);
  assign t[177] = t[235] ^ t[195];
  assign t[178] = t[236] ^ t[196];
  assign t[179] = t[197] & t[198];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[199] ^ t[63]);
  assign t[181] = t[39] ^ t[140];
  assign t[182] = t[200] ? x[102] : x[101];
  assign t[183] = ~(t[201]);
  assign t[184] = ~(t[65]);
  assign t[185] = t[28] ? x[104] : x[103];
  assign t[186] = t[25] ^ t[202];
  assign t[187] = ~(t[203] ^ t[23]);
  assign t[188] = t[204] ^ t[109];
  assign t[189] = t[72] ^ t[205];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[121] ^ t[55];
  assign t[191] = t[77] ? x[106] : x[105];
  assign t[192] = t[237] ^ t[206];
  assign t[193] = t[169] ? x[108] : x[107];
  assign t[194] = t[238] ^ t[207];
  assign t[195] = t[169] ? x[110] : x[109];
  assign t[196] = t[28] ? x[112] : x[111];
  assign t[197] = ~(t[161] ^ t[208]);
  assign t[198] = t[41] ^ t[201];
  assign t[199] = t[156] ^ t[61];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[49]);
  assign t[201] = t[68] ^ t[83];
  assign t[202] = t[129] ^ t[88];
  assign t[203] = ~(t[34] ^ t[82]);
  assign t[204] = t[133] ^ t[45];
  assign t[205] = t[209] & t[210];
  assign t[206] = t[200] ? x[114] : x[113];
  assign t[207] = t[200] ? x[116] : x[115];
  assign t[208] = t[122] ^ t[65];
  assign t[209] = ~(t[108] ^ t[211]);
  assign t[20] = ~(t[21] ^ t[26]);
  assign t[210] = t[204] ^ t[174];
  assign t[211] = t[151] ^ t[133];
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[35] ^ t[36];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[37] ^ t[38]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = t[266] ^ x[4];
  assign t[23] = t[39] ^ t[40];
  assign t[240] = t[267] ^ x[9];
  assign t[241] = t[268] ^ x[12];
  assign t[242] = t[269] ^ x[15];
  assign t[243] = t[270] ^ x[18];
  assign t[244] = t[271] ^ x[21];
  assign t[245] = t[272] ^ x[24];
  assign t[246] = t[273] ^ x[27];
  assign t[247] = t[274] ^ x[30];
  assign t[248] = t[275] ^ x[33];
  assign t[249] = t[276] ^ x[36];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[277] ^ x[39];
  assign t[251] = t[278] ^ x[42];
  assign t[252] = t[279] ^ x[45];
  assign t[253] = t[280] ^ x[48];
  assign t[254] = t[281] ^ x[51];
  assign t[255] = t[282] ^ x[54];
  assign t[256] = t[283] ^ x[59];
  assign t[257] = t[284] ^ x[62];
  assign t[258] = t[285] ^ x[67];
  assign t[259] = t[286] ^ x[70];
  assign t[25] = t[43] ^ t[44];
  assign t[260] = t[287] ^ x[77];
  assign t[261] = t[288] ^ x[82];
  assign t[262] = t[289] ^ x[85];
  assign t[263] = t[290] ^ x[88];
  assign t[264] = t[291] ^ x[91];
  assign t[265] = t[292] ^ x[100];
  assign t[266] = (t[293] & ~t[294]);
  assign t[267] = (t[295] & ~t[296]);
  assign t[268] = (t[297] & ~t[298]);
  assign t[269] = (t[299] & ~t[300]);
  assign t[26] = t[45] ^ t[46];
  assign t[270] = (t[301] & ~t[302]);
  assign t[271] = (t[303] & ~t[304]);
  assign t[272] = (t[305] & ~t[306]);
  assign t[273] = (t[307] & ~t[308]);
  assign t[274] = (t[309] & ~t[310]);
  assign t[275] = (t[311] & ~t[312]);
  assign t[276] = (t[313] & ~t[314]);
  assign t[277] = (t[315] & ~t[316]);
  assign t[278] = (t[317] & ~t[318]);
  assign t[279] = (t[319] & ~t[320]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = ~(t[49]);
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = t[347] ^ x[4];
  assign t[294] = t[348] ^ x[3];
  assign t[295] = t[349] ^ x[9];
  assign t[296] = t[350] ^ x[8];
  assign t[297] = t[351] ^ x[12];
  assign t[298] = t[352] ^ x[11];
  assign t[299] = t[353] ^ x[15];
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[14];
  assign t[301] = t[355] ^ x[18];
  assign t[302] = t[356] ^ x[17];
  assign t[303] = t[357] ^ x[21];
  assign t[304] = t[358] ^ x[20];
  assign t[305] = t[359] ^ x[24];
  assign t[306] = t[360] ^ x[23];
  assign t[307] = t[361] ^ x[27];
  assign t[308] = t[362] ^ x[26];
  assign t[309] = t[363] ^ x[30];
  assign t[30] = ~(t[214]);
  assign t[310] = t[364] ^ x[29];
  assign t[311] = t[365] ^ x[33];
  assign t[312] = t[366] ^ x[32];
  assign t[313] = t[367] ^ x[36];
  assign t[314] = t[368] ^ x[35];
  assign t[315] = t[369] ^ x[39];
  assign t[316] = t[370] ^ x[38];
  assign t[317] = t[371] ^ x[42];
  assign t[318] = t[372] ^ x[41];
  assign t[319] = t[373] ^ x[45];
  assign t[31] = ~(t[215]);
  assign t[320] = t[374] ^ x[44];
  assign t[321] = t[375] ^ x[48];
  assign t[322] = t[376] ^ x[47];
  assign t[323] = t[377] ^ x[51];
  assign t[324] = t[378] ^ x[50];
  assign t[325] = t[379] ^ x[54];
  assign t[326] = t[380] ^ x[53];
  assign t[327] = t[381] ^ x[59];
  assign t[328] = t[382] ^ x[58];
  assign t[329] = t[383] ^ x[62];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[61];
  assign t[331] = t[385] ^ x[67];
  assign t[332] = t[386] ^ x[66];
  assign t[333] = t[387] ^ x[70];
  assign t[334] = t[388] ^ x[69];
  assign t[335] = t[389] ^ x[77];
  assign t[336] = t[390] ^ x[76];
  assign t[337] = t[391] ^ x[82];
  assign t[338] = t[392] ^ x[81];
  assign t[339] = t[393] ^ x[85];
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[340] = t[394] ^ x[84];
  assign t[341] = t[395] ^ x[88];
  assign t[342] = t[396] ^ x[87];
  assign t[343] = t[397] ^ x[91];
  assign t[344] = t[398] ^ x[90];
  assign t[345] = t[399] ^ x[100];
  assign t[346] = t[400] ^ x[99];
  assign t[347] = (x[2]);
  assign t[348] = (x[2]);
  assign t[349] = (x[7]);
  assign t[34] = t[54] ^ t[55];
  assign t[350] = (x[7]);
  assign t[351] = (x[10]);
  assign t[352] = (x[10]);
  assign t[353] = (x[13]);
  assign t[354] = (x[13]);
  assign t[355] = (x[16]);
  assign t[356] = (x[16]);
  assign t[357] = (x[19]);
  assign t[358] = (x[19]);
  assign t[359] = (x[22]);
  assign t[35] = t[56] ^ t[43];
  assign t[360] = (x[22]);
  assign t[361] = (x[25]);
  assign t[362] = (x[25]);
  assign t[363] = (x[28]);
  assign t[364] = (x[28]);
  assign t[365] = (x[31]);
  assign t[366] = (x[31]);
  assign t[367] = (x[34]);
  assign t[368] = (x[34]);
  assign t[369] = (x[37]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[37]);
  assign t[371] = (x[40]);
  assign t[372] = (x[40]);
  assign t[373] = (x[43]);
  assign t[374] = (x[43]);
  assign t[375] = (x[46]);
  assign t[376] = (x[46]);
  assign t[377] = (x[49]);
  assign t[378] = (x[49]);
  assign t[379] = (x[52]);
  assign t[37] = t[59] ^ t[33];
  assign t[380] = (x[52]);
  assign t[381] = (x[57]);
  assign t[382] = (x[57]);
  assign t[383] = (x[60]);
  assign t[384] = (x[60]);
  assign t[385] = (x[65]);
  assign t[386] = (x[65]);
  assign t[387] = (x[68]);
  assign t[388] = (x[68]);
  assign t[389] = (x[75]);
  assign t[38] = ~(t[25] ^ t[60]);
  assign t[390] = (x[75]);
  assign t[391] = (x[80]);
  assign t[392] = (x[80]);
  assign t[393] = (x[83]);
  assign t[394] = (x[83]);
  assign t[395] = (x[86]);
  assign t[396] = (x[86]);
  assign t[397] = (x[89]);
  assign t[398] = (x[89]);
  assign t[399] = (x[98]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[98]);
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] & t[68];
  assign t[43] = t[8] ? t[69] : t[216];
  assign t[44] = t[57] ^ t[70];
  assign t[45] = t[217] ^ t[71];
  assign t[46] = t[72] ^ t[73];
  assign t[47] = ~(t[74] & t[75]);
  assign t[48] = t[218] | t[76];
  assign t[49] = ~(t[77]);
  assign t[4] = t[8] ? t[9] : t[212];
  assign t[50] = ~(t[219]);
  assign t[51] = ~(t[78] & t[217]);
  assign t[52] = t[79] ^ t[80];
  assign t[53] = ~(t[81] ^ t[82]);
  assign t[54] = t[65] ^ t[83];
  assign t[55] = t[84] & t[85];
  assign t[56] = t[8] ? t[86] : t[220];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] & t[90];
  assign t[59] = ~(t[91] ^ t[92]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] ^ t[73];
  assign t[61] = t[94] ? t[95] : t[221];
  assign t[62] = t[94] ? t[96] : t[222];
  assign t[63] = t[97] ^ t[98];
  assign t[64] = t[99] & t[100];
  assign t[65] = ~t[101];
  assign t[66] = ~t[102];
  assign t[67] = ~(t[83]);
  assign t[68] = t[103];
  assign t[69] = t[216] ^ t[104];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[105] & t[106];
  assign t[71] = t[8] ? t[107] : t[223];
  assign t[72] = t[108] ^ t[109];
  assign t[73] = t[110] & t[111];
  assign t[74] = ~(t[76] & t[112]);
  assign t[75] = ~(t[224] ^ t[113]);
  assign t[76] = ~(t[114] & t[115]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[225]);
  assign t[79] = t[116] ^ t[98];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] ^ t[70];
  assign t[81] = t[118] ^ t[60];
  assign t[82] = t[62] ^ t[119];
  assign t[83] = t[120];
  assign t[84] = ~(t[54] ^ t[121]);
  assign t[85] = t[122] ^ t[68];
  assign t[86] = t[220] ^ t[123];
  assign t[87] = t[124] & t[125];
  assign t[88] = t[126] & t[127];
  assign t[89] = ~(t[87] ^ t[128]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[131] ^ t[24];
  assign t[92] = ~(t[132] ^ t[80]);
  assign t[93] = t[133] ^ t[134];
  assign t[94] = ~(t[15]);
  assign t[95] = t[221] ^ t[135];
  assign t[96] = t[222] ^ t[136];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[139] & t[140];
  assign t[99] = ~(t[97] ^ t[141]);
  assign t[9] = t[212] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [116:0] x;
 output y;

 wire [400:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[116] ^ t[142];
  assign t[101] = t[27] ? t[143] : t[226];
  assign t[102] = t[27] ? t[144] : t[227];
  assign t[103] = t[27] ? t[145] : t[228];
  assign t[104] = t[28] ? x[56] : x[55];
  assign t[105] = ~(t[117] ^ t[57]);
  assign t[106] = t[35] ^ t[127];
  assign t[107] = t[223] ^ t[146];
  assign t[108] = t[147] & t[148];
  assign t[109] = t[149] & t[150];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[93] ^ t[72]);
  assign t[111] = t[151] ^ t[150];
  assign t[112] = ~(t[152] & t[153]);
  assign t[113] = t[154] ^ t[229];
  assign t[114] = ~(t[224]);
  assign t[115] = t[155] & t[154];
  assign t[116] = t[156] ^ t[62];
  assign t[117] = t[157] ^ t[56];
  assign t[118] = t[122] ^ t[158];
  assign t[119] = t[63] ^ t[159];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[27] ? t[160] : t[230];
  assign t[121] = t[161] ^ t[42];
  assign t[122] = t[83] ^ t[66];
  assign t[123] = t[28] ? x[64] : x[63];
  assign t[124] = ~(t[130]);
  assign t[125] = ~(t[157]);
  assign t[126] = ~(t[56]);
  assign t[127] = t[8] ? t[162] : t[231];
  assign t[128] = t[35] ^ t[157];
  assign t[129] = t[157] ^ t[43];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[127] ^ t[56];
  assign t[131] = ~(t[163] ^ t[164]);
  assign t[132] = t[165] ^ t[166];
  assign t[133] = t[8] ? t[167] : t[232];
  assign t[134] = t[213] ^ t[168];
  assign t[135] = t[169] ? x[72] : x[71];
  assign t[136] = t[169] ? x[74] : x[73];
  assign t[137] = ~(t[142]);
  assign t[138] = ~(t[156]);
  assign t[139] = ~(t[61]);
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[94] ? t[170] : t[233];
  assign t[141] = t[39] ^ t[156];
  assign t[142] = t[140] ^ t[61];
  assign t[143] = t[226] ^ t[171];
  assign t[144] = t[227] ^ t[172];
  assign t[145] = t[228] ^ t[173];
  assign t[146] = t[77] ? x[79] : x[78];
  assign t[147] = ~(t[174]);
  assign t[148] = ~(t[133]);
  assign t[149] = ~(t[134]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[214] ^ t[175];
  assign t[151] = t[134] ^ t[45];
  assign t[152] = ~(t[155] | t[154]);
  assign t[153] = ~(t[176] | t[114]);
  assign t[154] = ~(t[234]);
  assign t[155] = ~(t[229]);
  assign t[156] = t[94] ? t[177] : t[235];
  assign t[157] = t[8] ? t[178] : t[236];
  assign t[158] = t[121] ^ t[179];
  assign t[159] = t[180] & t[181];
  assign t[15] = ~(t[27]);
  assign t[160] = t[230] ^ t[182];
  assign t[161] = t[183] & t[184];
  assign t[162] = t[231] ^ t[185];
  assign t[163] = t[186] ^ t[187];
  assign t[164] = ~(t[188] ^ t[26]);
  assign t[165] = t[151] ^ t[189];
  assign t[166] = t[66] ^ t[190];
  assign t[167] = t[232] ^ t[191];
  assign t[168] = t[27] ? t[192] : t[237];
  assign t[169] = ~(t[49]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[233] ^ t[193];
  assign t[171] = t[77] ? x[93] : x[92];
  assign t[172] = t[77] ? x[95] : x[94];
  assign t[173] = t[28] ? x[97] : x[96];
  assign t[174] = t[150] ^ t[134];
  assign t[175] = t[8] ? t[194] : t[238];
  assign t[176] = ~(t[218]);
  assign t[177] = t[235] ^ t[195];
  assign t[178] = t[236] ^ t[196];
  assign t[179] = t[197] & t[198];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = ~(t[199] ^ t[63]);
  assign t[181] = t[39] ^ t[140];
  assign t[182] = t[200] ? x[102] : x[101];
  assign t[183] = ~(t[201]);
  assign t[184] = ~(t[65]);
  assign t[185] = t[28] ? x[104] : x[103];
  assign t[186] = t[25] ^ t[202];
  assign t[187] = ~(t[203] ^ t[23]);
  assign t[188] = t[204] ^ t[109];
  assign t[189] = t[72] ^ t[205];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[121] ^ t[55];
  assign t[191] = t[77] ? x[106] : x[105];
  assign t[192] = t[237] ^ t[206];
  assign t[193] = t[169] ? x[108] : x[107];
  assign t[194] = t[238] ^ t[207];
  assign t[195] = t[169] ? x[110] : x[109];
  assign t[196] = t[28] ? x[112] : x[111];
  assign t[197] = ~(t[161] ^ t[208]);
  assign t[198] = t[41] ^ t[201];
  assign t[199] = t[156] ^ t[61];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[49]);
  assign t[201] = t[68] ^ t[83];
  assign t[202] = t[129] ^ t[88];
  assign t[203] = ~(t[34] ^ t[82]);
  assign t[204] = t[133] ^ t[45];
  assign t[205] = t[209] & t[210];
  assign t[206] = t[200] ? x[114] : x[113];
  assign t[207] = t[200] ? x[116] : x[115];
  assign t[208] = t[122] ^ t[65];
  assign t[209] = ~(t[108] ^ t[211]);
  assign t[20] = ~(t[21] ^ t[26]);
  assign t[210] = t[204] ^ t[174];
  assign t[211] = t[151] ^ t[133];
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[35] ^ t[36];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[37] ^ t[38]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = t[266] ^ x[4];
  assign t[23] = t[39] ^ t[40];
  assign t[240] = t[267] ^ x[9];
  assign t[241] = t[268] ^ x[12];
  assign t[242] = t[269] ^ x[15];
  assign t[243] = t[270] ^ x[18];
  assign t[244] = t[271] ^ x[21];
  assign t[245] = t[272] ^ x[24];
  assign t[246] = t[273] ^ x[27];
  assign t[247] = t[274] ^ x[30];
  assign t[248] = t[275] ^ x[33];
  assign t[249] = t[276] ^ x[36];
  assign t[24] = t[41] ^ t[42];
  assign t[250] = t[277] ^ x[39];
  assign t[251] = t[278] ^ x[42];
  assign t[252] = t[279] ^ x[45];
  assign t[253] = t[280] ^ x[48];
  assign t[254] = t[281] ^ x[51];
  assign t[255] = t[282] ^ x[54];
  assign t[256] = t[283] ^ x[59];
  assign t[257] = t[284] ^ x[62];
  assign t[258] = t[285] ^ x[67];
  assign t[259] = t[286] ^ x[70];
  assign t[25] = t[43] ^ t[44];
  assign t[260] = t[287] ^ x[77];
  assign t[261] = t[288] ^ x[82];
  assign t[262] = t[289] ^ x[85];
  assign t[263] = t[290] ^ x[88];
  assign t[264] = t[291] ^ x[91];
  assign t[265] = t[292] ^ x[100];
  assign t[266] = (t[293] & ~t[294]);
  assign t[267] = (t[295] & ~t[296]);
  assign t[268] = (t[297] & ~t[298]);
  assign t[269] = (t[299] & ~t[300]);
  assign t[26] = t[45] ^ t[46];
  assign t[270] = (t[301] & ~t[302]);
  assign t[271] = (t[303] & ~t[304]);
  assign t[272] = (t[305] & ~t[306]);
  assign t[273] = (t[307] & ~t[308]);
  assign t[274] = (t[309] & ~t[310]);
  assign t[275] = (t[311] & ~t[312]);
  assign t[276] = (t[313] & ~t[314]);
  assign t[277] = (t[315] & ~t[316]);
  assign t[278] = (t[317] & ~t[318]);
  assign t[279] = (t[319] & ~t[320]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = ~(t[49]);
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = t[347] ^ x[4];
  assign t[294] = t[348] ^ x[3];
  assign t[295] = t[349] ^ x[9];
  assign t[296] = t[350] ^ x[8];
  assign t[297] = t[351] ^ x[12];
  assign t[298] = t[352] ^ x[11];
  assign t[299] = t[353] ^ x[15];
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[14];
  assign t[301] = t[355] ^ x[18];
  assign t[302] = t[356] ^ x[17];
  assign t[303] = t[357] ^ x[21];
  assign t[304] = t[358] ^ x[20];
  assign t[305] = t[359] ^ x[24];
  assign t[306] = t[360] ^ x[23];
  assign t[307] = t[361] ^ x[27];
  assign t[308] = t[362] ^ x[26];
  assign t[309] = t[363] ^ x[30];
  assign t[30] = ~(t[214]);
  assign t[310] = t[364] ^ x[29];
  assign t[311] = t[365] ^ x[33];
  assign t[312] = t[366] ^ x[32];
  assign t[313] = t[367] ^ x[36];
  assign t[314] = t[368] ^ x[35];
  assign t[315] = t[369] ^ x[39];
  assign t[316] = t[370] ^ x[38];
  assign t[317] = t[371] ^ x[42];
  assign t[318] = t[372] ^ x[41];
  assign t[319] = t[373] ^ x[45];
  assign t[31] = ~(t[215]);
  assign t[320] = t[374] ^ x[44];
  assign t[321] = t[375] ^ x[48];
  assign t[322] = t[376] ^ x[47];
  assign t[323] = t[377] ^ x[51];
  assign t[324] = t[378] ^ x[50];
  assign t[325] = t[379] ^ x[54];
  assign t[326] = t[380] ^ x[53];
  assign t[327] = t[381] ^ x[59];
  assign t[328] = t[382] ^ x[58];
  assign t[329] = t[383] ^ x[62];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[61];
  assign t[331] = t[385] ^ x[67];
  assign t[332] = t[386] ^ x[66];
  assign t[333] = t[387] ^ x[70];
  assign t[334] = t[388] ^ x[69];
  assign t[335] = t[389] ^ x[77];
  assign t[336] = t[390] ^ x[76];
  assign t[337] = t[391] ^ x[82];
  assign t[338] = t[392] ^ x[81];
  assign t[339] = t[393] ^ x[85];
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[340] = t[394] ^ x[84];
  assign t[341] = t[395] ^ x[88];
  assign t[342] = t[396] ^ x[87];
  assign t[343] = t[397] ^ x[91];
  assign t[344] = t[398] ^ x[90];
  assign t[345] = t[399] ^ x[100];
  assign t[346] = t[400] ^ x[99];
  assign t[347] = (x[2]);
  assign t[348] = (x[2]);
  assign t[349] = (x[7]);
  assign t[34] = t[54] ^ t[55];
  assign t[350] = (x[7]);
  assign t[351] = (x[10]);
  assign t[352] = (x[10]);
  assign t[353] = (x[13]);
  assign t[354] = (x[13]);
  assign t[355] = (x[16]);
  assign t[356] = (x[16]);
  assign t[357] = (x[19]);
  assign t[358] = (x[19]);
  assign t[359] = (x[22]);
  assign t[35] = t[56] ^ t[43];
  assign t[360] = (x[22]);
  assign t[361] = (x[25]);
  assign t[362] = (x[25]);
  assign t[363] = (x[28]);
  assign t[364] = (x[28]);
  assign t[365] = (x[31]);
  assign t[366] = (x[31]);
  assign t[367] = (x[34]);
  assign t[368] = (x[34]);
  assign t[369] = (x[37]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[37]);
  assign t[371] = (x[40]);
  assign t[372] = (x[40]);
  assign t[373] = (x[43]);
  assign t[374] = (x[43]);
  assign t[375] = (x[46]);
  assign t[376] = (x[46]);
  assign t[377] = (x[49]);
  assign t[378] = (x[49]);
  assign t[379] = (x[52]);
  assign t[37] = t[59] ^ t[33];
  assign t[380] = (x[52]);
  assign t[381] = (x[57]);
  assign t[382] = (x[57]);
  assign t[383] = (x[60]);
  assign t[384] = (x[60]);
  assign t[385] = (x[65]);
  assign t[386] = (x[65]);
  assign t[387] = (x[68]);
  assign t[388] = (x[68]);
  assign t[389] = (x[75]);
  assign t[38] = ~(t[25] ^ t[60]);
  assign t[390] = (x[75]);
  assign t[391] = (x[80]);
  assign t[392] = (x[80]);
  assign t[393] = (x[83]);
  assign t[394] = (x[83]);
  assign t[395] = (x[86]);
  assign t[396] = (x[86]);
  assign t[397] = (x[89]);
  assign t[398] = (x[89]);
  assign t[399] = (x[98]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[98]);
  assign t[40] = t[63] ^ t[64];
  assign t[41] = t[65] ^ t[66];
  assign t[42] = t[67] & t[68];
  assign t[43] = t[8] ? t[69] : t[216];
  assign t[44] = t[57] ^ t[70];
  assign t[45] = t[217] ^ t[71];
  assign t[46] = t[72] ^ t[73];
  assign t[47] = ~(t[74] & t[75]);
  assign t[48] = t[218] | t[76];
  assign t[49] = ~(t[77]);
  assign t[4] = t[8] ? t[9] : t[212];
  assign t[50] = ~(t[219]);
  assign t[51] = ~(t[78] & t[217]);
  assign t[52] = t[79] ^ t[80];
  assign t[53] = ~(t[81] ^ t[82]);
  assign t[54] = t[65] ^ t[83];
  assign t[55] = t[84] & t[85];
  assign t[56] = t[8] ? t[86] : t[220];
  assign t[57] = t[87] ^ t[88];
  assign t[58] = t[89] & t[90];
  assign t[59] = ~(t[91] ^ t[92]);
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] ^ t[73];
  assign t[61] = t[94] ? t[95] : t[221];
  assign t[62] = t[94] ? t[96] : t[222];
  assign t[63] = t[97] ^ t[98];
  assign t[64] = t[99] & t[100];
  assign t[65] = ~t[101];
  assign t[66] = ~t[102];
  assign t[67] = ~(t[83]);
  assign t[68] = t[103];
  assign t[69] = t[216] ^ t[104];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[105] & t[106];
  assign t[71] = t[8] ? t[107] : t[223];
  assign t[72] = t[108] ^ t[109];
  assign t[73] = t[110] & t[111];
  assign t[74] = ~(t[76] & t[112]);
  assign t[75] = ~(t[224] ^ t[113]);
  assign t[76] = ~(t[114] & t[115]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[225]);
  assign t[79] = t[116] ^ t[98];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] ^ t[70];
  assign t[81] = t[118] ^ t[60];
  assign t[82] = t[62] ^ t[119];
  assign t[83] = t[120];
  assign t[84] = ~(t[54] ^ t[121]);
  assign t[85] = t[122] ^ t[68];
  assign t[86] = t[220] ^ t[123];
  assign t[87] = t[124] & t[125];
  assign t[88] = t[126] & t[127];
  assign t[89] = ~(t[87] ^ t[128]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[129] ^ t[130];
  assign t[91] = t[131] ^ t[24];
  assign t[92] = ~(t[132] ^ t[80]);
  assign t[93] = t[133] ^ t[134];
  assign t[94] = ~(t[15]);
  assign t[95] = t[221] ^ t[135];
  assign t[96] = t[222] ^ t[136];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[139] & t[140];
  assign t[99] = ~(t[97] ^ t[141]);
  assign t[9] = t[212] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind146(x, y);
 input [116:0] x;
 output y;

 wire [409:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[53] ^ t[140];
  assign t[101] = t[141] ^ t[142];
  assign t[102] = t[143] ^ t[144];
  assign t[103] = t[129] ^ t[60];
  assign t[104] = t[42] ^ t[86];
  assign t[105] = t[145] ^ t[146];
  assign t[106] = ~t[147];
  assign t[107] = ~(t[70] ^ t[98]);
  assign t[108] = t[65] ^ t[148];
  assign t[109] = t[8] ? t[149] : t[233];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[150] ^ t[64];
  assign t[111] = t[151] & t[152];
  assign t[112] = ~(t[153] & t[154]);
  assign t[113] = t[155] ^ t[234];
  assign t[114] = ~(t[229]);
  assign t[115] = t[156] & t[155];
  assign t[116] = t[8] ? t[157] : t[235];
  assign t[117] = ~(t[83]);
  assign t[118] = t[8] ? t[158] : t[236];
  assign t[119] = t[222] ^ t[159];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[160] & t[161];
  assign t[121] = t[231] ^ t[162];
  assign t[122] = ~(t[88] ^ t[163]);
  assign t[123] = t[79] ^ t[164];
  assign t[124] = t[22] ^ t[165];
  assign t[125] = ~(t[100] ^ t[103]);
  assign t[126] = t[93] ^ t[119];
  assign t[127] = ~(t[164]);
  assign t[128] = ~(t[116]);
  assign t[129] = t[116] ^ t[83];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[166] ^ t[145];
  assign t[131] = t[167] ^ t[168];
  assign t[132] = t[232] ^ t[169];
  assign t[133] = t[8] ? t[170] : t[237];
  assign t[134] = t[27] ? t[171] : t[238];
  assign t[135] = t[27] ? t[172] : t[239];
  assign t[136] = t[173] & t[174];
  assign t[137] = t[175] & t[148];
  assign t[138] = ~(t[136] ^ t[176]);
  assign t[139] = t[177] ^ t[178];
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[97] ^ t[179];
  assign t[141] = t[180] ^ t[166];
  assign t[142] = t[181] & t[182];
  assign t[143] = t[180] ^ t[145];
  assign t[144] = t[183] & t[184];
  assign t[145] = t[185] ? t[186] : t[240];
  assign t[146] = t[167] ^ t[142];
  assign t[147] = t[27] ? t[187] : t[241];
  assign t[148] = t[188];
  assign t[149] = t[233] ^ t[189];
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[190] & t[191];
  assign t[151] = ~(t[126] ^ t[110]);
  assign t[152] = t[81] ^ t[95];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[192] | t[114]);
  assign t[155] = ~(t[242]);
  assign t[156] = ~(t[234]);
  assign t[157] = t[235] ^ t[193];
  assign t[158] = t[236] ^ t[194];
  assign t[159] = t[27] ? t[195] : t[243];
  assign t[15] = ~(t[27]);
  assign t[160] = ~(t[150] ^ t[196]);
  assign t[161] = t[63] ^ t[197];
  assign t[162] = t[28] ? x[76] : x[75];
  assign t[163] = t[54] ^ t[116];
  assign t[164] = t[118] ^ t[83];
  assign t[165] = t[177] ^ t[137];
  assign t[166] = t[185] ? t[198] : t[244];
  assign t[167] = t[199] ^ t[144];
  assign t[168] = t[200] & t[201];
  assign t[169] = t[77] ? x[81] : x[80];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[237] ^ t[202];
  assign t[171] = t[238] ^ t[203];
  assign t[172] = t[239] ^ t[204];
  assign t[173] = ~(t[178]);
  assign t[174] = ~(t[106]);
  assign t[175] = ~(t[96]);
  assign t[176] = t[65] ^ t[106];
  assign t[177] = t[106] ^ t[97];
  assign t[178] = t[148] ^ t[96];
  assign t[179] = t[98] ^ t[71];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[185] ? t[205] : t[245];
  assign t[181] = ~(t[141] ^ t[167]);
  assign t[182] = t[130] ^ t[184];
  assign t[183] = ~(t[166]);
  assign t[184] = t[185] ? t[206] : t[246];
  assign t[185] = ~(t[15]);
  assign t[186] = t[240] ^ t[207];
  assign t[187] = t[241] ^ t[208];
  assign t[188] = t[27] ? t[209] : t[247];
  assign t[189] = t[77] ? x[92] : x[91];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = ~(t[197]);
  assign t[191] = ~(t[93]);
  assign t[192] = ~(t[226]);
  assign t[193] = t[28] ? x[94] : x[93];
  assign t[194] = t[28] ? x[96] : x[95];
  assign t[195] = t[243] ^ t[210];
  assign t[196] = t[81] ^ t[93];
  assign t[197] = t[95] ^ t[119];
  assign t[198] = t[244] ^ t[211];
  assign t[199] = t[212] & t[213];
  assign t[19] = ~(t[33] ^ t[34]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[199] ^ t[214]);
  assign t[201] = t[143] ^ t[215];
  assign t[202] = t[216] ? x[98] : x[97];
  assign t[203] = t[216] ? x[100] : x[99];
  assign t[204] = t[77] ? x[102] : x[101];
  assign t[205] = t[245] ^ t[217];
  assign t[206] = t[246] ^ t[218];
  assign t[207] = t[219] ? x[104] : x[103];
  assign t[208] = t[77] ? x[106] : x[105];
  assign t[209] = t[247] ^ t[220];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[216] ? x[108] : x[107];
  assign t[211] = t[219] ? x[110] : x[109];
  assign t[212] = ~(t[215]);
  assign t[213] = ~(t[180]);
  assign t[214] = t[130] ^ t[180];
  assign t[215] = t[184] ^ t[166];
  assign t[216] = ~(t[49]);
  assign t[217] = t[219] ? x[112] : x[111];
  assign t[218] = t[219] ? x[114] : x[113];
  assign t[219] = ~(t[49]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[28] ? x[116] : x[115];
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[39] ^ t[40]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = (t[266]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (t[267]);
  assign t[241] = (t[268]);
  assign t[242] = (t[269]);
  assign t[243] = (t[270]);
  assign t[244] = (t[271]);
  assign t[245] = (t[272]);
  assign t[246] = (t[273]);
  assign t[247] = (t[274]);
  assign t[248] = t[275] ^ x[4];
  assign t[249] = t[276] ^ x[9];
  assign t[24] = ~(t[43] ^ t[21]);
  assign t[250] = t[277] ^ x[12];
  assign t[251] = t[278] ^ x[15];
  assign t[252] = t[279] ^ x[18];
  assign t[253] = t[280] ^ x[21];
  assign t[254] = t[281] ^ x[24];
  assign t[255] = t[282] ^ x[27];
  assign t[256] = t[283] ^ x[30];
  assign t[257] = t[284] ^ x[33];
  assign t[258] = t[285] ^ x[36];
  assign t[259] = t[286] ^ x[41];
  assign t[25] = t[44] ^ t[45];
  assign t[260] = t[287] ^ x[44];
  assign t[261] = t[288] ^ x[47];
  assign t[262] = t[289] ^ x[50];
  assign t[263] = t[290] ^ x[53];
  assign t[264] = t[291] ^ x[56];
  assign t[265] = t[292] ^ x[59];
  assign t[266] = t[293] ^ x[62];
  assign t[267] = t[294] ^ x[65];
  assign t[268] = t[295] ^ x[68];
  assign t[269] = t[296] ^ x[71];
  assign t[26] = ~(t[35] ^ t[46]);
  assign t[270] = t[297] ^ x[74];
  assign t[271] = t[298] ^ x[79];
  assign t[272] = t[299] ^ x[84];
  assign t[273] = t[300] ^ x[87];
  assign t[274] = t[301] ^ x[90];
  assign t[275] = (t[302] & ~t[303]);
  assign t[276] = (t[304] & ~t[305]);
  assign t[277] = (t[306] & ~t[307]);
  assign t[278] = (t[308] & ~t[309]);
  assign t[279] = (t[310] & ~t[311]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[312] & ~t[313]);
  assign t[281] = (t[314] & ~t[315]);
  assign t[282] = (t[316] & ~t[317]);
  assign t[283] = (t[318] & ~t[319]);
  assign t[284] = (t[320] & ~t[321]);
  assign t[285] = (t[322] & ~t[323]);
  assign t[286] = (t[324] & ~t[325]);
  assign t[287] = (t[326] & ~t[327]);
  assign t[288] = (t[328] & ~t[329]);
  assign t[289] = (t[330] & ~t[331]);
  assign t[28] = ~(t[49]);
  assign t[290] = (t[332] & ~t[333]);
  assign t[291] = (t[334] & ~t[335]);
  assign t[292] = (t[336] & ~t[337]);
  assign t[293] = (t[338] & ~t[339]);
  assign t[294] = (t[340] & ~t[341]);
  assign t[295] = (t[342] & ~t[343]);
  assign t[296] = (t[344] & ~t[345]);
  assign t[297] = (t[346] & ~t[347]);
  assign t[298] = (t[348] & ~t[349]);
  assign t[299] = (t[350] & ~t[351]);
  assign t[29] = ~(t[222]);
  assign t[2] = ~(t[5]);
  assign t[300] = (t[352] & ~t[353]);
  assign t[301] = (t[354] & ~t[355]);
  assign t[302] = t[356] ^ x[4];
  assign t[303] = t[357] ^ x[3];
  assign t[304] = t[358] ^ x[9];
  assign t[305] = t[359] ^ x[8];
  assign t[306] = t[360] ^ x[12];
  assign t[307] = t[361] ^ x[11];
  assign t[308] = t[362] ^ x[15];
  assign t[309] = t[363] ^ x[14];
  assign t[30] = ~(t[223]);
  assign t[310] = t[364] ^ x[18];
  assign t[311] = t[365] ^ x[17];
  assign t[312] = t[366] ^ x[21];
  assign t[313] = t[367] ^ x[20];
  assign t[314] = t[368] ^ x[24];
  assign t[315] = t[369] ^ x[23];
  assign t[316] = t[370] ^ x[27];
  assign t[317] = t[371] ^ x[26];
  assign t[318] = t[372] ^ x[30];
  assign t[319] = t[373] ^ x[29];
  assign t[31] = ~(t[224]);
  assign t[320] = t[374] ^ x[33];
  assign t[321] = t[375] ^ x[32];
  assign t[322] = t[376] ^ x[36];
  assign t[323] = t[377] ^ x[35];
  assign t[324] = t[378] ^ x[41];
  assign t[325] = t[379] ^ x[40];
  assign t[326] = t[380] ^ x[44];
  assign t[327] = t[381] ^ x[43];
  assign t[328] = t[382] ^ x[47];
  assign t[329] = t[383] ^ x[46];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[50];
  assign t[331] = t[385] ^ x[49];
  assign t[332] = t[386] ^ x[53];
  assign t[333] = t[387] ^ x[52];
  assign t[334] = t[388] ^ x[56];
  assign t[335] = t[389] ^ x[55];
  assign t[336] = t[390] ^ x[59];
  assign t[337] = t[391] ^ x[58];
  assign t[338] = t[392] ^ x[62];
  assign t[339] = t[393] ^ x[61];
  assign t[33] = t[52] ^ t[14];
  assign t[340] = t[394] ^ x[65];
  assign t[341] = t[395] ^ x[64];
  assign t[342] = t[396] ^ x[68];
  assign t[343] = t[397] ^ x[67];
  assign t[344] = t[398] ^ x[71];
  assign t[345] = t[399] ^ x[70];
  assign t[346] = t[400] ^ x[74];
  assign t[347] = t[401] ^ x[73];
  assign t[348] = t[402] ^ x[79];
  assign t[349] = t[403] ^ x[78];
  assign t[34] = ~(t[53] ^ t[43]);
  assign t[350] = t[404] ^ x[84];
  assign t[351] = t[405] ^ x[83];
  assign t[352] = t[406] ^ x[87];
  assign t[353] = t[407] ^ x[86];
  assign t[354] = t[408] ^ x[90];
  assign t[355] = t[409] ^ x[89];
  assign t[356] = (x[2]);
  assign t[357] = (x[2]);
  assign t[358] = (x[7]);
  assign t[359] = (x[7]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[10]);
  assign t[361] = (x[10]);
  assign t[362] = (x[13]);
  assign t[363] = (x[13]);
  assign t[364] = (x[16]);
  assign t[365] = (x[16]);
  assign t[366] = (x[19]);
  assign t[367] = (x[19]);
  assign t[368] = (x[22]);
  assign t[369] = (x[22]);
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[370] = (x[25]);
  assign t[371] = (x[25]);
  assign t[372] = (x[28]);
  assign t[373] = (x[28]);
  assign t[374] = (x[31]);
  assign t[375] = (x[31]);
  assign t[376] = (x[34]);
  assign t[377] = (x[34]);
  assign t[378] = (x[39]);
  assign t[379] = (x[39]);
  assign t[37] = t[8] ? t[58] : t[225];
  assign t[380] = (x[42]);
  assign t[381] = (x[42]);
  assign t[382] = (x[45]);
  assign t[383] = (x[45]);
  assign t[384] = (x[48]);
  assign t[385] = (x[48]);
  assign t[386] = (x[51]);
  assign t[387] = (x[51]);
  assign t[388] = (x[54]);
  assign t[389] = (x[54]);
  assign t[38] = t[59] ^ t[60];
  assign t[390] = (x[57]);
  assign t[391] = (x[57]);
  assign t[392] = (x[60]);
  assign t[393] = (x[60]);
  assign t[394] = (x[63]);
  assign t[395] = (x[63]);
  assign t[396] = (x[66]);
  assign t[397] = (x[66]);
  assign t[398] = (x[69]);
  assign t[399] = (x[69]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[72]);
  assign t[401] = (x[72]);
  assign t[402] = (x[77]);
  assign t[403] = (x[77]);
  assign t[404] = (x[82]);
  assign t[405] = (x[82]);
  assign t[406] = (x[85]);
  assign t[407] = (x[85]);
  assign t[408] = (x[88]);
  assign t[409] = (x[88]);
  assign t[40] = ~(t[41] ^ t[46]);
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[67] ^ t[35]);
  assign t[44] = ~(t[68] ^ t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] ^ t[73];
  assign t[47] = ~(t[74] & t[75]);
  assign t[48] = t[226] | t[76];
  assign t[49] = ~(t[77]);
  assign t[4] = t[8] ? t[9] : t[221];
  assign t[50] = ~(t[227]);
  assign t[51] = ~(t[78] & t[228]);
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] ^ t[37];
  assign t[55] = t[59] ^ t[84];
  assign t[56] = t[85] ^ t[44];
  assign t[57] = ~(t[21] ^ t[86]);
  assign t[58] = t[225] ^ t[87];
  assign t[59] = t[88] ^ t[80];
  assign t[5] = ~(t[10]);
  assign t[60] = t[89] & t[90];
  assign t[61] = t[21] ^ t[52];
  assign t[62] = ~(t[91] ^ t[92]);
  assign t[63] = t[93] ^ t[72];
  assign t[64] = t[94] & t[95];
  assign t[65] = t[96] ^ t[97];
  assign t[66] = t[98] ^ t[99];
  assign t[67] = ~(t[100] ^ t[101]);
  assign t[68] = t[102] ^ t[103];
  assign t[69] = ~(t[104] ^ t[105]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[106] ^ t[96];
  assign t[71] = t[107] & t[108];
  assign t[72] = t[228] ^ t[109];
  assign t[73] = t[110] ^ t[111];
  assign t[74] = ~(t[76] & t[112]);
  assign t[75] = ~(t[229] ^ t[113]);
  assign t[76] = ~(t[114] & t[115]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[230]);
  assign t[79] = t[116] ^ t[37];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] & t[118];
  assign t[81] = t[119] ^ t[72];
  assign t[82] = t[110] ^ t[120];
  assign t[83] = t[8] ? t[121] : t[231];
  assign t[84] = t[122] & t[123];
  assign t[85] = ~(t[124] ^ t[125]);
  assign t[86] = t[126] ^ t[111];
  assign t[87] = t[28] ? x[38] : x[37];
  assign t[88] = t[127] & t[128];
  assign t[89] = ~(t[129] ^ t[59]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[54] ^ t[118];
  assign t[91] = ~(t[45] ^ t[105]);
  assign t[92] = t[130] ^ t[131];
  assign t[93] = t[8] ? t[132] : t[232];
  assign t[94] = ~(t[119]);
  assign t[95] = t[223] ^ t[133];
  assign t[96] = t[134];
  assign t[97] = ~t[135];
  assign t[98] = t[136] ^ t[137];
  assign t[99] = t[138] & t[139];
  assign t[9] = t[221] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [116:0] x;
 output y;

 wire [409:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[53] ^ t[140];
  assign t[101] = t[141] ^ t[142];
  assign t[102] = t[143] ^ t[144];
  assign t[103] = t[129] ^ t[60];
  assign t[104] = t[42] ^ t[86];
  assign t[105] = t[145] ^ t[146];
  assign t[106] = ~t[147];
  assign t[107] = ~(t[70] ^ t[98]);
  assign t[108] = t[65] ^ t[148];
  assign t[109] = t[8] ? t[149] : t[233];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[150] ^ t[64];
  assign t[111] = t[151] & t[152];
  assign t[112] = ~(t[153] & t[154]);
  assign t[113] = t[155] ^ t[234];
  assign t[114] = ~(t[229]);
  assign t[115] = t[156] & t[155];
  assign t[116] = t[8] ? t[157] : t[235];
  assign t[117] = ~(t[83]);
  assign t[118] = t[8] ? t[158] : t[236];
  assign t[119] = t[222] ^ t[159];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[160] & t[161];
  assign t[121] = t[231] ^ t[162];
  assign t[122] = ~(t[88] ^ t[163]);
  assign t[123] = t[79] ^ t[164];
  assign t[124] = t[22] ^ t[165];
  assign t[125] = ~(t[100] ^ t[103]);
  assign t[126] = t[93] ^ t[119];
  assign t[127] = ~(t[164]);
  assign t[128] = ~(t[116]);
  assign t[129] = t[116] ^ t[83];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[166] ^ t[145];
  assign t[131] = t[167] ^ t[168];
  assign t[132] = t[232] ^ t[169];
  assign t[133] = t[8] ? t[170] : t[237];
  assign t[134] = t[27] ? t[171] : t[238];
  assign t[135] = t[27] ? t[172] : t[239];
  assign t[136] = t[173] & t[174];
  assign t[137] = t[175] & t[148];
  assign t[138] = ~(t[136] ^ t[176]);
  assign t[139] = t[177] ^ t[178];
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[97] ^ t[179];
  assign t[141] = t[180] ^ t[166];
  assign t[142] = t[181] & t[182];
  assign t[143] = t[180] ^ t[145];
  assign t[144] = t[183] & t[184];
  assign t[145] = t[185] ? t[186] : t[240];
  assign t[146] = t[167] ^ t[142];
  assign t[147] = t[27] ? t[187] : t[241];
  assign t[148] = t[188];
  assign t[149] = t[233] ^ t[189];
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = t[190] & t[191];
  assign t[151] = ~(t[126] ^ t[110]);
  assign t[152] = t[81] ^ t[95];
  assign t[153] = ~(t[156] | t[155]);
  assign t[154] = ~(t[192] | t[114]);
  assign t[155] = ~(t[242]);
  assign t[156] = ~(t[234]);
  assign t[157] = t[235] ^ t[193];
  assign t[158] = t[236] ^ t[194];
  assign t[159] = t[27] ? t[195] : t[243];
  assign t[15] = ~(t[27]);
  assign t[160] = ~(t[150] ^ t[196]);
  assign t[161] = t[63] ^ t[197];
  assign t[162] = t[28] ? x[76] : x[75];
  assign t[163] = t[54] ^ t[116];
  assign t[164] = t[118] ^ t[83];
  assign t[165] = t[177] ^ t[137];
  assign t[166] = t[185] ? t[198] : t[244];
  assign t[167] = t[199] ^ t[144];
  assign t[168] = t[200] & t[201];
  assign t[169] = t[77] ? x[81] : x[80];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = t[237] ^ t[202];
  assign t[171] = t[238] ^ t[203];
  assign t[172] = t[239] ^ t[204];
  assign t[173] = ~(t[178]);
  assign t[174] = ~(t[106]);
  assign t[175] = ~(t[96]);
  assign t[176] = t[65] ^ t[106];
  assign t[177] = t[106] ^ t[97];
  assign t[178] = t[148] ^ t[96];
  assign t[179] = t[98] ^ t[71];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[185] ? t[205] : t[245];
  assign t[181] = ~(t[141] ^ t[167]);
  assign t[182] = t[130] ^ t[184];
  assign t[183] = ~(t[166]);
  assign t[184] = t[185] ? t[206] : t[246];
  assign t[185] = ~(t[15]);
  assign t[186] = t[240] ^ t[207];
  assign t[187] = t[241] ^ t[208];
  assign t[188] = t[27] ? t[209] : t[247];
  assign t[189] = t[77] ? x[92] : x[91];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = ~(t[197]);
  assign t[191] = ~(t[93]);
  assign t[192] = ~(t[226]);
  assign t[193] = t[28] ? x[94] : x[93];
  assign t[194] = t[28] ? x[96] : x[95];
  assign t[195] = t[243] ^ t[210];
  assign t[196] = t[81] ^ t[93];
  assign t[197] = t[95] ^ t[119];
  assign t[198] = t[244] ^ t[211];
  assign t[199] = t[212] & t[213];
  assign t[19] = ~(t[33] ^ t[34]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[199] ^ t[214]);
  assign t[201] = t[143] ^ t[215];
  assign t[202] = t[216] ? x[98] : x[97];
  assign t[203] = t[216] ? x[100] : x[99];
  assign t[204] = t[77] ? x[102] : x[101];
  assign t[205] = t[245] ^ t[217];
  assign t[206] = t[246] ^ t[218];
  assign t[207] = t[219] ? x[104] : x[103];
  assign t[208] = t[77] ? x[106] : x[105];
  assign t[209] = t[247] ^ t[220];
  assign t[20] = t[35] ^ t[36];
  assign t[210] = t[216] ? x[108] : x[107];
  assign t[211] = t[219] ? x[110] : x[109];
  assign t[212] = ~(t[215]);
  assign t[213] = ~(t[180]);
  assign t[214] = t[130] ^ t[180];
  assign t[215] = t[184] ^ t[166];
  assign t[216] = ~(t[49]);
  assign t[217] = t[219] ? x[112] : x[111];
  assign t[218] = t[219] ? x[114] : x[113];
  assign t[219] = ~(t[49]);
  assign t[21] = t[37] ^ t[38];
  assign t[220] = t[28] ? x[116] : x[115];
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[39] ^ t[40]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = (t[266]);
  assign t[23] = t[41] ^ t[42];
  assign t[240] = (t[267]);
  assign t[241] = (t[268]);
  assign t[242] = (t[269]);
  assign t[243] = (t[270]);
  assign t[244] = (t[271]);
  assign t[245] = (t[272]);
  assign t[246] = (t[273]);
  assign t[247] = (t[274]);
  assign t[248] = t[275] ^ x[4];
  assign t[249] = t[276] ^ x[9];
  assign t[24] = ~(t[43] ^ t[21]);
  assign t[250] = t[277] ^ x[12];
  assign t[251] = t[278] ^ x[15];
  assign t[252] = t[279] ^ x[18];
  assign t[253] = t[280] ^ x[21];
  assign t[254] = t[281] ^ x[24];
  assign t[255] = t[282] ^ x[27];
  assign t[256] = t[283] ^ x[30];
  assign t[257] = t[284] ^ x[33];
  assign t[258] = t[285] ^ x[36];
  assign t[259] = t[286] ^ x[41];
  assign t[25] = t[44] ^ t[45];
  assign t[260] = t[287] ^ x[44];
  assign t[261] = t[288] ^ x[47];
  assign t[262] = t[289] ^ x[50];
  assign t[263] = t[290] ^ x[53];
  assign t[264] = t[291] ^ x[56];
  assign t[265] = t[292] ^ x[59];
  assign t[266] = t[293] ^ x[62];
  assign t[267] = t[294] ^ x[65];
  assign t[268] = t[295] ^ x[68];
  assign t[269] = t[296] ^ x[71];
  assign t[26] = ~(t[35] ^ t[46]);
  assign t[270] = t[297] ^ x[74];
  assign t[271] = t[298] ^ x[79];
  assign t[272] = t[299] ^ x[84];
  assign t[273] = t[300] ^ x[87];
  assign t[274] = t[301] ^ x[90];
  assign t[275] = (t[302] & ~t[303]);
  assign t[276] = (t[304] & ~t[305]);
  assign t[277] = (t[306] & ~t[307]);
  assign t[278] = (t[308] & ~t[309]);
  assign t[279] = (t[310] & ~t[311]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[280] = (t[312] & ~t[313]);
  assign t[281] = (t[314] & ~t[315]);
  assign t[282] = (t[316] & ~t[317]);
  assign t[283] = (t[318] & ~t[319]);
  assign t[284] = (t[320] & ~t[321]);
  assign t[285] = (t[322] & ~t[323]);
  assign t[286] = (t[324] & ~t[325]);
  assign t[287] = (t[326] & ~t[327]);
  assign t[288] = (t[328] & ~t[329]);
  assign t[289] = (t[330] & ~t[331]);
  assign t[28] = ~(t[49]);
  assign t[290] = (t[332] & ~t[333]);
  assign t[291] = (t[334] & ~t[335]);
  assign t[292] = (t[336] & ~t[337]);
  assign t[293] = (t[338] & ~t[339]);
  assign t[294] = (t[340] & ~t[341]);
  assign t[295] = (t[342] & ~t[343]);
  assign t[296] = (t[344] & ~t[345]);
  assign t[297] = (t[346] & ~t[347]);
  assign t[298] = (t[348] & ~t[349]);
  assign t[299] = (t[350] & ~t[351]);
  assign t[29] = ~(t[222]);
  assign t[2] = ~(t[5]);
  assign t[300] = (t[352] & ~t[353]);
  assign t[301] = (t[354] & ~t[355]);
  assign t[302] = t[356] ^ x[4];
  assign t[303] = t[357] ^ x[3];
  assign t[304] = t[358] ^ x[9];
  assign t[305] = t[359] ^ x[8];
  assign t[306] = t[360] ^ x[12];
  assign t[307] = t[361] ^ x[11];
  assign t[308] = t[362] ^ x[15];
  assign t[309] = t[363] ^ x[14];
  assign t[30] = ~(t[223]);
  assign t[310] = t[364] ^ x[18];
  assign t[311] = t[365] ^ x[17];
  assign t[312] = t[366] ^ x[21];
  assign t[313] = t[367] ^ x[20];
  assign t[314] = t[368] ^ x[24];
  assign t[315] = t[369] ^ x[23];
  assign t[316] = t[370] ^ x[27];
  assign t[317] = t[371] ^ x[26];
  assign t[318] = t[372] ^ x[30];
  assign t[319] = t[373] ^ x[29];
  assign t[31] = ~(t[224]);
  assign t[320] = t[374] ^ x[33];
  assign t[321] = t[375] ^ x[32];
  assign t[322] = t[376] ^ x[36];
  assign t[323] = t[377] ^ x[35];
  assign t[324] = t[378] ^ x[41];
  assign t[325] = t[379] ^ x[40];
  assign t[326] = t[380] ^ x[44];
  assign t[327] = t[381] ^ x[43];
  assign t[328] = t[382] ^ x[47];
  assign t[329] = t[383] ^ x[46];
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = t[384] ^ x[50];
  assign t[331] = t[385] ^ x[49];
  assign t[332] = t[386] ^ x[53];
  assign t[333] = t[387] ^ x[52];
  assign t[334] = t[388] ^ x[56];
  assign t[335] = t[389] ^ x[55];
  assign t[336] = t[390] ^ x[59];
  assign t[337] = t[391] ^ x[58];
  assign t[338] = t[392] ^ x[62];
  assign t[339] = t[393] ^ x[61];
  assign t[33] = t[52] ^ t[14];
  assign t[340] = t[394] ^ x[65];
  assign t[341] = t[395] ^ x[64];
  assign t[342] = t[396] ^ x[68];
  assign t[343] = t[397] ^ x[67];
  assign t[344] = t[398] ^ x[71];
  assign t[345] = t[399] ^ x[70];
  assign t[346] = t[400] ^ x[74];
  assign t[347] = t[401] ^ x[73];
  assign t[348] = t[402] ^ x[79];
  assign t[349] = t[403] ^ x[78];
  assign t[34] = ~(t[53] ^ t[43]);
  assign t[350] = t[404] ^ x[84];
  assign t[351] = t[405] ^ x[83];
  assign t[352] = t[406] ^ x[87];
  assign t[353] = t[407] ^ x[86];
  assign t[354] = t[408] ^ x[90];
  assign t[355] = t[409] ^ x[89];
  assign t[356] = (x[2]);
  assign t[357] = (x[2]);
  assign t[358] = (x[7]);
  assign t[359] = (x[7]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[10]);
  assign t[361] = (x[10]);
  assign t[362] = (x[13]);
  assign t[363] = (x[13]);
  assign t[364] = (x[16]);
  assign t[365] = (x[16]);
  assign t[366] = (x[19]);
  assign t[367] = (x[19]);
  assign t[368] = (x[22]);
  assign t[369] = (x[22]);
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[370] = (x[25]);
  assign t[371] = (x[25]);
  assign t[372] = (x[28]);
  assign t[373] = (x[28]);
  assign t[374] = (x[31]);
  assign t[375] = (x[31]);
  assign t[376] = (x[34]);
  assign t[377] = (x[34]);
  assign t[378] = (x[39]);
  assign t[379] = (x[39]);
  assign t[37] = t[8] ? t[58] : t[225];
  assign t[380] = (x[42]);
  assign t[381] = (x[42]);
  assign t[382] = (x[45]);
  assign t[383] = (x[45]);
  assign t[384] = (x[48]);
  assign t[385] = (x[48]);
  assign t[386] = (x[51]);
  assign t[387] = (x[51]);
  assign t[388] = (x[54]);
  assign t[389] = (x[54]);
  assign t[38] = t[59] ^ t[60];
  assign t[390] = (x[57]);
  assign t[391] = (x[57]);
  assign t[392] = (x[60]);
  assign t[393] = (x[60]);
  assign t[394] = (x[63]);
  assign t[395] = (x[63]);
  assign t[396] = (x[66]);
  assign t[397] = (x[66]);
  assign t[398] = (x[69]);
  assign t[399] = (x[69]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[72]);
  assign t[401] = (x[72]);
  assign t[402] = (x[77]);
  assign t[403] = (x[77]);
  assign t[404] = (x[82]);
  assign t[405] = (x[82]);
  assign t[406] = (x[85]);
  assign t[407] = (x[85]);
  assign t[408] = (x[88]);
  assign t[409] = (x[88]);
  assign t[40] = ~(t[41] ^ t[46]);
  assign t[41] = t[63] ^ t[64];
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[67] ^ t[35]);
  assign t[44] = ~(t[68] ^ t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = t[72] ^ t[73];
  assign t[47] = ~(t[74] & t[75]);
  assign t[48] = t[226] | t[76];
  assign t[49] = ~(t[77]);
  assign t[4] = t[8] ? t[9] : t[221];
  assign t[50] = ~(t[227]);
  assign t[51] = ~(t[78] & t[228]);
  assign t[52] = t[79] ^ t[80];
  assign t[53] = t[81] ^ t[82];
  assign t[54] = t[83] ^ t[37];
  assign t[55] = t[59] ^ t[84];
  assign t[56] = t[85] ^ t[44];
  assign t[57] = ~(t[21] ^ t[86]);
  assign t[58] = t[225] ^ t[87];
  assign t[59] = t[88] ^ t[80];
  assign t[5] = ~(t[10]);
  assign t[60] = t[89] & t[90];
  assign t[61] = t[21] ^ t[52];
  assign t[62] = ~(t[91] ^ t[92]);
  assign t[63] = t[93] ^ t[72];
  assign t[64] = t[94] & t[95];
  assign t[65] = t[96] ^ t[97];
  assign t[66] = t[98] ^ t[99];
  assign t[67] = ~(t[100] ^ t[101]);
  assign t[68] = t[102] ^ t[103];
  assign t[69] = ~(t[104] ^ t[105]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[106] ^ t[96];
  assign t[71] = t[107] & t[108];
  assign t[72] = t[228] ^ t[109];
  assign t[73] = t[110] ^ t[111];
  assign t[74] = ~(t[76] & t[112]);
  assign t[75] = ~(t[229] ^ t[113]);
  assign t[76] = ~(t[114] & t[115]);
  assign t[77] = ~(t[48]);
  assign t[78] = ~(t[230]);
  assign t[79] = t[116] ^ t[37];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[117] & t[118];
  assign t[81] = t[119] ^ t[72];
  assign t[82] = t[110] ^ t[120];
  assign t[83] = t[8] ? t[121] : t[231];
  assign t[84] = t[122] & t[123];
  assign t[85] = ~(t[124] ^ t[125]);
  assign t[86] = t[126] ^ t[111];
  assign t[87] = t[28] ? x[38] : x[37];
  assign t[88] = t[127] & t[128];
  assign t[89] = ~(t[129] ^ t[59]);
  assign t[8] = ~(t[15]);
  assign t[90] = t[54] ^ t[118];
  assign t[91] = ~(t[45] ^ t[105]);
  assign t[92] = t[130] ^ t[131];
  assign t[93] = t[8] ? t[132] : t[232];
  assign t[94] = ~(t[119]);
  assign t[95] = t[223] ^ t[133];
  assign t[96] = t[134];
  assign t[97] = ~t[135];
  assign t[98] = t[136] ^ t[137];
  assign t[99] = t[138] & t[139];
  assign t[9] = t[221] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [116:0] x;
 output y;

 wire [400:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[139] ^ t[132];
  assign t[101] = t[213] ^ t[140];
  assign t[102] = t[141] ^ t[106];
  assign t[103] = t[142] & t[143];
  assign t[104] = t[8] ? t[144] : t[227];
  assign t[105] = t[123] ^ t[67];
  assign t[106] = t[145] & t[146];
  assign t[107] = t[8] ? t[147] : t[228];
  assign t[108] = t[119] ^ t[54];
  assign t[109] = t[148] ^ t[121];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[149] & t[150]);
  assign t[111] = t[151] ^ t[229];
  assign t[112] = ~(t[220]);
  assign t[113] = t[152] & t[151];
  assign t[114] = t[222] ^ t[153];
  assign t[115] = t[88] ? t[154] : t[230];
  assign t[116] = t[223] ^ t[155];
  assign t[117] = t[224] ^ t[156];
  assign t[118] = t[225] ^ t[157];
  assign t[119] = t[158] ^ t[159];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[8] ? t[160] : t[231];
  assign t[121] = t[161];
  assign t[122] = t[162] & t[163];
  assign t[123] = t[8] ? t[164] : t[232];
  assign t[124] = ~(t[86] ^ t[102]);
  assign t[125] = t[65] ^ t[146];
  assign t[126] = t[165] ? x[68] : x[67];
  assign t[127] = t[166] & t[167];
  assign t[128] = ~(t[135] ^ t[90]);
  assign t[129] = t[137] ^ t[79];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[226] ^ t[168];
  assign t[131] = t[169] & t[170];
  assign t[132] = t[171] & t[172];
  assign t[133] = ~(t[109] ^ t[93]);
  assign t[134] = t[84] ^ t[172];
  assign t[135] = t[77] ^ t[115];
  assign t[136] = t[173] & t[174];
  assign t[137] = t[115] ^ t[57];
  assign t[138] = t[90] ^ t[175];
  assign t[139] = t[148] ^ t[59];
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[27] ? t[176] : t[233];
  assign t[141] = t[177] & t[178];
  assign t[142] = ~(t[141] ^ t[179]);
  assign t[143] = t[105] ^ t[180];
  assign t[144] = t[227] ^ t[181];
  assign t[145] = ~(t[101]);
  assign t[146] = t[214] ^ t[182];
  assign t[147] = t[228] ^ t[183];
  assign t[148] = ~t[184];
  assign t[149] = ~(t[152] | t[151]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[185] | t[112]);
  assign t[151] = ~(t[234]);
  assign t[152] = ~(t[229]);
  assign t[153] = t[165] ? x[76] : x[75];
  assign t[154] = t[230] ^ t[186];
  assign t[155] = t[165] ? x[78] : x[77];
  assign t[156] = t[28] ? x[80] : x[79];
  assign t[157] = t[28] ? x[82] : x[81];
  assign t[158] = t[187] & t[188];
  assign t[159] = t[189] & t[120];
  assign t[15] = ~(t[27]);
  assign t[160] = t[231] ^ t[190];
  assign t[161] = t[27] ? t[191] : t[235];
  assign t[162] = ~(t[131] ^ t[192]);
  assign t[163] = t[139] ^ t[193];
  assign t[164] = t[232] ^ t[194];
  assign t[165] = ~(t[48]);
  assign t[166] = ~(t[195]);
  assign t[167] = ~(t[77]);
  assign t[168] = t[75] ? x[87] : x[86];
  assign t[169] = ~(t[193]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[148]);
  assign t[171] = ~(t[121]);
  assign t[172] = t[196];
  assign t[173] = ~(t[158] ^ t[197]);
  assign t[174] = t[198] ^ t[199];
  assign t[175] = t[200] & t[201];
  assign t[176] = t[233] ^ t[202];
  assign t[177] = ~(t[180]);
  assign t[178] = ~(t[123]);
  assign t[179] = t[65] ^ t[123];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[146] ^ t[101];
  assign t[181] = t[75] ? x[89] : x[88];
  assign t[182] = t[8] ? t[203] : t[236];
  assign t[183] = t[28] ? x[94] : x[93];
  assign t[184] = t[27] ? t[204] : t[237];
  assign t[185] = ~(t[216]);
  assign t[186] = t[165] ? x[99] : x[98];
  assign t[187] = ~(t[199]);
  assign t[188] = ~(t[80]);
  assign t[189] = ~(t[81]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[28] ? x[101] : x[100];
  assign t[191] = t[235] ^ t[205];
  assign t[192] = t[84] ^ t[148];
  assign t[193] = t[172] ^ t[121];
  assign t[194] = t[75] ? x[103] : x[102];
  assign t[195] = t[79] ^ t[115];
  assign t[196] = t[27] ? t[206] : t[238];
  assign t[197] = t[97] ^ t[80];
  assign t[198] = t[80] ^ t[107];
  assign t[199] = t[120] ^ t[81];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[127] ^ t[207]);
  assign t[201] = t[51] ^ t[195];
  assign t[202] = t[208] ? x[108] : x[107];
  assign t[203] = t[236] ^ t[209];
  assign t[204] = t[237] ^ t[210];
  assign t[205] = t[208] ? x[110] : x[109];
  assign t[206] = t[238] ^ t[211];
  assign t[207] = t[137] ^ t[77];
  assign t[208] = ~(t[48]);
  assign t[209] = t[208] ? x[112] : x[111];
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = t[75] ? x[114] : x[113];
  assign t[211] = t[28] ? x[116] : x[115];
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[35]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[38] ^ t[39];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = t[266] ^ x[4];
  assign t[23] = t[22] ^ t[34];
  assign t[240] = t[267] ^ x[9];
  assign t[241] = t[268] ^ x[12];
  assign t[242] = t[269] ^ x[15];
  assign t[243] = t[270] ^ x[18];
  assign t[244] = t[271] ^ x[21];
  assign t[245] = t[272] ^ x[24];
  assign t[246] = t[273] ^ x[27];
  assign t[247] = t[274] ^ x[30];
  assign t[248] = t[275] ^ x[33];
  assign t[249] = t[276] ^ x[36];
  assign t[24] = ~(t[40] ^ t[41]);
  assign t[250] = t[277] ^ x[39];
  assign t[251] = t[278] ^ x[42];
  assign t[252] = t[279] ^ x[45];
  assign t[253] = t[280] ^ x[48];
  assign t[254] = t[281] ^ x[51];
  assign t[255] = t[282] ^ x[54];
  assign t[256] = t[283] ^ x[57];
  assign t[257] = t[284] ^ x[60];
  assign t[258] = t[285] ^ x[63];
  assign t[259] = t[286] ^ x[66];
  assign t[25] = ~(t[42] ^ t[43]);
  assign t[260] = t[287] ^ x[71];
  assign t[261] = t[288] ^ x[74];
  assign t[262] = t[289] ^ x[85];
  assign t[263] = t[290] ^ x[92];
  assign t[264] = t[291] ^ x[97];
  assign t[265] = t[292] ^ x[106];
  assign t[266] = (t[293] & ~t[294]);
  assign t[267] = (t[295] & ~t[296]);
  assign t[268] = (t[297] & ~t[298]);
  assign t[269] = (t[299] & ~t[300]);
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[270] = (t[301] & ~t[302]);
  assign t[271] = (t[303] & ~t[304]);
  assign t[272] = (t[305] & ~t[306]);
  assign t[273] = (t[307] & ~t[308]);
  assign t[274] = (t[309] & ~t[310]);
  assign t[275] = (t[311] & ~t[312]);
  assign t[276] = (t[313] & ~t[314]);
  assign t[277] = (t[315] & ~t[316]);
  assign t[278] = (t[317] & ~t[318]);
  assign t[279] = (t[319] & ~t[320]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = t[347] ^ x[4];
  assign t[294] = t[348] ^ x[3];
  assign t[295] = t[349] ^ x[9];
  assign t[296] = t[350] ^ x[8];
  assign t[297] = t[351] ^ x[12];
  assign t[298] = t[352] ^ x[11];
  assign t[299] = t[353] ^ x[15];
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[14];
  assign t[301] = t[355] ^ x[18];
  assign t[302] = t[356] ^ x[17];
  assign t[303] = t[357] ^ x[21];
  assign t[304] = t[358] ^ x[20];
  assign t[305] = t[359] ^ x[24];
  assign t[306] = t[360] ^ x[23];
  assign t[307] = t[361] ^ x[27];
  assign t[308] = t[362] ^ x[26];
  assign t[309] = t[363] ^ x[30];
  assign t[30] = ~(t[214]);
  assign t[310] = t[364] ^ x[29];
  assign t[311] = t[365] ^ x[33];
  assign t[312] = t[366] ^ x[32];
  assign t[313] = t[367] ^ x[36];
  assign t[314] = t[368] ^ x[35];
  assign t[315] = t[369] ^ x[39];
  assign t[316] = t[370] ^ x[38];
  assign t[317] = t[371] ^ x[42];
  assign t[318] = t[372] ^ x[41];
  assign t[319] = t[373] ^ x[45];
  assign t[31] = ~(t[215]);
  assign t[320] = t[374] ^ x[44];
  assign t[321] = t[375] ^ x[48];
  assign t[322] = t[376] ^ x[47];
  assign t[323] = t[377] ^ x[51];
  assign t[324] = t[378] ^ x[50];
  assign t[325] = t[379] ^ x[54];
  assign t[326] = t[380] ^ x[53];
  assign t[327] = t[381] ^ x[57];
  assign t[328] = t[382] ^ x[56];
  assign t[329] = t[383] ^ x[60];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[59];
  assign t[331] = t[385] ^ x[63];
  assign t[332] = t[386] ^ x[62];
  assign t[333] = t[387] ^ x[66];
  assign t[334] = t[388] ^ x[65];
  assign t[335] = t[389] ^ x[71];
  assign t[336] = t[390] ^ x[70];
  assign t[337] = t[391] ^ x[74];
  assign t[338] = t[392] ^ x[73];
  assign t[339] = t[393] ^ x[85];
  assign t[33] = t[51] ^ t[52];
  assign t[340] = t[394] ^ x[84];
  assign t[341] = t[395] ^ x[92];
  assign t[342] = t[396] ^ x[91];
  assign t[343] = t[397] ^ x[97];
  assign t[344] = t[398] ^ x[96];
  assign t[345] = t[399] ^ x[106];
  assign t[346] = t[400] ^ x[105];
  assign t[347] = (x[2]);
  assign t[348] = (x[2]);
  assign t[349] = (x[7]);
  assign t[34] = t[53] ^ t[54];
  assign t[350] = (x[7]);
  assign t[351] = (x[10]);
  assign t[352] = (x[10]);
  assign t[353] = (x[13]);
  assign t[354] = (x[13]);
  assign t[355] = (x[16]);
  assign t[356] = (x[16]);
  assign t[357] = (x[19]);
  assign t[358] = (x[19]);
  assign t[359] = (x[22]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[22]);
  assign t[361] = (x[25]);
  assign t[362] = (x[25]);
  assign t[363] = (x[28]);
  assign t[364] = (x[28]);
  assign t[365] = (x[31]);
  assign t[366] = (x[31]);
  assign t[367] = (x[34]);
  assign t[368] = (x[34]);
  assign t[369] = (x[37]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[37]);
  assign t[371] = (x[40]);
  assign t[372] = (x[40]);
  assign t[373] = (x[43]);
  assign t[374] = (x[43]);
  assign t[375] = (x[46]);
  assign t[376] = (x[46]);
  assign t[377] = (x[49]);
  assign t[378] = (x[49]);
  assign t[379] = (x[52]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[52]);
  assign t[381] = (x[55]);
  assign t[382] = (x[55]);
  assign t[383] = (x[58]);
  assign t[384] = (x[58]);
  assign t[385] = (x[61]);
  assign t[386] = (x[61]);
  assign t[387] = (x[64]);
  assign t[388] = (x[64]);
  assign t[389] = (x[69]);
  assign t[38] = ~(t[61] ^ t[62]);
  assign t[390] = (x[69]);
  assign t[391] = (x[72]);
  assign t[392] = (x[72]);
  assign t[393] = (x[83]);
  assign t[394] = (x[83]);
  assign t[395] = (x[90]);
  assign t[396] = (x[90]);
  assign t[397] = (x[95]);
  assign t[398] = (x[95]);
  assign t[399] = (x[104]);
  assign t[39] = ~(t[63] ^ t[64]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[104]);
  assign t[40] = t[65] ^ t[66];
  assign t[41] = t[67] ^ t[68];
  assign t[42] = t[69] ^ t[55];
  assign t[43] = ~(t[38] ^ t[70]);
  assign t[44] = t[11] ^ t[71];
  assign t[45] = ~(t[62] ^ t[41]);
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[216] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[217]);
  assign t[4] = t[8] ? t[9] : t[212];
  assign t[50] = ~(t[76] & t[218]);
  assign t[51] = t[77] ^ t[57];
  assign t[52] = t[78] & t[79];
  assign t[53] = t[80] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = t[84] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ? t[89] : t[219];
  assign t[58] = t[90] ^ t[91];
  assign t[59] = ~t[92];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] ^ t[94];
  assign t[61] = ~(t[95] ^ t[96]);
  assign t[62] = t[97] ^ t[98];
  assign t[63] = t[99] ^ t[100];
  assign t[64] = ~(t[70] ^ t[41]);
  assign t[65] = t[101] ^ t[67];
  assign t[66] = t[102] ^ t[103];
  assign t[67] = t[218] ^ t[104];
  assign t[68] = t[102] ^ t[87];
  assign t[69] = t[105] ^ t[106];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[107] ^ t[108];
  assign t[71] = t[109] ^ t[94];
  assign t[72] = ~(t[74] & t[110]);
  assign t[73] = ~(t[220] ^ t[111]);
  assign t[74] = ~(t[112] & t[113]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[221]);
  assign t[77] = t[88] ? t[114] : t[222];
  assign t[78] = ~(t[115]);
  assign t[79] = t[88] ? t[116] : t[223];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[117] : t[224];
  assign t[81] = t[8] ? t[118] : t[225];
  assign t[82] = ~(t[53] ^ t[119]);
  assign t[83] = t[97] ^ t[120];
  assign t[84] = t[121] ^ t[59];
  assign t[85] = t[93] ^ t[122];
  assign t[86] = t[123] ^ t[101];
  assign t[87] = t[124] & t[125];
  assign t[88] = ~(t[15]);
  assign t[89] = t[219] ^ t[126];
  assign t[8] = ~(t[15]);
  assign t[90] = t[127] ^ t[52];
  assign t[91] = t[128] & t[129];
  assign t[92] = t[27] ? t[130] : t[226];
  assign t[93] = t[131] ^ t[132];
  assign t[94] = t[133] & t[134];
  assign t[95] = t[40] ^ t[37];
  assign t[96] = t[135] ^ t[91];
  assign t[97] = t[81] ^ t[107];
  assign t[98] = t[119] ^ t[136];
  assign t[99] = t[137] ^ t[138];
  assign t[9] = t[212] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [116:0] x;
 output y;

 wire [400:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[139] ^ t[132];
  assign t[101] = t[213] ^ t[140];
  assign t[102] = t[141] ^ t[106];
  assign t[103] = t[142] & t[143];
  assign t[104] = t[8] ? t[144] : t[227];
  assign t[105] = t[123] ^ t[67];
  assign t[106] = t[145] & t[146];
  assign t[107] = t[8] ? t[147] : t[228];
  assign t[108] = t[119] ^ t[54];
  assign t[109] = t[148] ^ t[121];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = ~(t[149] & t[150]);
  assign t[111] = t[151] ^ t[229];
  assign t[112] = ~(t[220]);
  assign t[113] = t[152] & t[151];
  assign t[114] = t[222] ^ t[153];
  assign t[115] = t[88] ? t[154] : t[230];
  assign t[116] = t[223] ^ t[155];
  assign t[117] = t[224] ^ t[156];
  assign t[118] = t[225] ^ t[157];
  assign t[119] = t[158] ^ t[159];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[8] ? t[160] : t[231];
  assign t[121] = t[161];
  assign t[122] = t[162] & t[163];
  assign t[123] = t[8] ? t[164] : t[232];
  assign t[124] = ~(t[86] ^ t[102]);
  assign t[125] = t[65] ^ t[146];
  assign t[126] = t[165] ? x[68] : x[67];
  assign t[127] = t[166] & t[167];
  assign t[128] = ~(t[135] ^ t[90]);
  assign t[129] = t[137] ^ t[79];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[226] ^ t[168];
  assign t[131] = t[169] & t[170];
  assign t[132] = t[171] & t[172];
  assign t[133] = ~(t[109] ^ t[93]);
  assign t[134] = t[84] ^ t[172];
  assign t[135] = t[77] ^ t[115];
  assign t[136] = t[173] & t[174];
  assign t[137] = t[115] ^ t[57];
  assign t[138] = t[90] ^ t[175];
  assign t[139] = t[148] ^ t[59];
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[27] ? t[176] : t[233];
  assign t[141] = t[177] & t[178];
  assign t[142] = ~(t[141] ^ t[179]);
  assign t[143] = t[105] ^ t[180];
  assign t[144] = t[227] ^ t[181];
  assign t[145] = ~(t[101]);
  assign t[146] = t[214] ^ t[182];
  assign t[147] = t[228] ^ t[183];
  assign t[148] = ~t[184];
  assign t[149] = ~(t[152] | t[151]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[150] = ~(t[185] | t[112]);
  assign t[151] = ~(t[234]);
  assign t[152] = ~(t[229]);
  assign t[153] = t[165] ? x[76] : x[75];
  assign t[154] = t[230] ^ t[186];
  assign t[155] = t[165] ? x[78] : x[77];
  assign t[156] = t[28] ? x[80] : x[79];
  assign t[157] = t[28] ? x[82] : x[81];
  assign t[158] = t[187] & t[188];
  assign t[159] = t[189] & t[120];
  assign t[15] = ~(t[27]);
  assign t[160] = t[231] ^ t[190];
  assign t[161] = t[27] ? t[191] : t[235];
  assign t[162] = ~(t[131] ^ t[192]);
  assign t[163] = t[139] ^ t[193];
  assign t[164] = t[232] ^ t[194];
  assign t[165] = ~(t[48]);
  assign t[166] = ~(t[195]);
  assign t[167] = ~(t[77]);
  assign t[168] = t[75] ? x[87] : x[86];
  assign t[169] = ~(t[193]);
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[148]);
  assign t[171] = ~(t[121]);
  assign t[172] = t[196];
  assign t[173] = ~(t[158] ^ t[197]);
  assign t[174] = t[198] ^ t[199];
  assign t[175] = t[200] & t[201];
  assign t[176] = t[233] ^ t[202];
  assign t[177] = ~(t[180]);
  assign t[178] = ~(t[123]);
  assign t[179] = t[65] ^ t[123];
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[146] ^ t[101];
  assign t[181] = t[75] ? x[89] : x[88];
  assign t[182] = t[8] ? t[203] : t[236];
  assign t[183] = t[28] ? x[94] : x[93];
  assign t[184] = t[27] ? t[204] : t[237];
  assign t[185] = ~(t[216]);
  assign t[186] = t[165] ? x[99] : x[98];
  assign t[187] = ~(t[199]);
  assign t[188] = ~(t[80]);
  assign t[189] = ~(t[81]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[28] ? x[101] : x[100];
  assign t[191] = t[235] ^ t[205];
  assign t[192] = t[84] ^ t[148];
  assign t[193] = t[172] ^ t[121];
  assign t[194] = t[75] ? x[103] : x[102];
  assign t[195] = t[79] ^ t[115];
  assign t[196] = t[27] ? t[206] : t[238];
  assign t[197] = t[97] ^ t[80];
  assign t[198] = t[80] ^ t[107];
  assign t[199] = t[120] ^ t[81];
  assign t[19] = t[33] ^ t[34];
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = ~(t[127] ^ t[207]);
  assign t[201] = t[51] ^ t[195];
  assign t[202] = t[208] ? x[108] : x[107];
  assign t[203] = t[236] ^ t[209];
  assign t[204] = t[237] ^ t[210];
  assign t[205] = t[208] ? x[110] : x[109];
  assign t[206] = t[238] ^ t[211];
  assign t[207] = t[137] ^ t[77];
  assign t[208] = ~(t[48]);
  assign t[209] = t[208] ? x[112] : x[111];
  assign t[20] = ~(t[35] ^ t[36]);
  assign t[210] = t[75] ? x[114] : x[113];
  assign t[211] = t[28] ? x[116] : x[115];
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = ~(t[37] ^ t[35]);
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = t[38] ^ t[39];
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = (t[264]);
  assign t[238] = (t[265]);
  assign t[239] = t[266] ^ x[4];
  assign t[23] = t[22] ^ t[34];
  assign t[240] = t[267] ^ x[9];
  assign t[241] = t[268] ^ x[12];
  assign t[242] = t[269] ^ x[15];
  assign t[243] = t[270] ^ x[18];
  assign t[244] = t[271] ^ x[21];
  assign t[245] = t[272] ^ x[24];
  assign t[246] = t[273] ^ x[27];
  assign t[247] = t[274] ^ x[30];
  assign t[248] = t[275] ^ x[33];
  assign t[249] = t[276] ^ x[36];
  assign t[24] = ~(t[40] ^ t[41]);
  assign t[250] = t[277] ^ x[39];
  assign t[251] = t[278] ^ x[42];
  assign t[252] = t[279] ^ x[45];
  assign t[253] = t[280] ^ x[48];
  assign t[254] = t[281] ^ x[51];
  assign t[255] = t[282] ^ x[54];
  assign t[256] = t[283] ^ x[57];
  assign t[257] = t[284] ^ x[60];
  assign t[258] = t[285] ^ x[63];
  assign t[259] = t[286] ^ x[66];
  assign t[25] = ~(t[42] ^ t[43]);
  assign t[260] = t[287] ^ x[71];
  assign t[261] = t[288] ^ x[74];
  assign t[262] = t[289] ^ x[85];
  assign t[263] = t[290] ^ x[92];
  assign t[264] = t[291] ^ x[97];
  assign t[265] = t[292] ^ x[106];
  assign t[266] = (t[293] & ~t[294]);
  assign t[267] = (t[295] & ~t[296]);
  assign t[268] = (t[297] & ~t[298]);
  assign t[269] = (t[299] & ~t[300]);
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[270] = (t[301] & ~t[302]);
  assign t[271] = (t[303] & ~t[304]);
  assign t[272] = (t[305] & ~t[306]);
  assign t[273] = (t[307] & ~t[308]);
  assign t[274] = (t[309] & ~t[310]);
  assign t[275] = (t[311] & ~t[312]);
  assign t[276] = (t[313] & ~t[314]);
  assign t[277] = (t[315] & ~t[316]);
  assign t[278] = (t[317] & ~t[318]);
  assign t[279] = (t[319] & ~t[320]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[321] & ~t[322]);
  assign t[281] = (t[323] & ~t[324]);
  assign t[282] = (t[325] & ~t[326]);
  assign t[283] = (t[327] & ~t[328]);
  assign t[284] = (t[329] & ~t[330]);
  assign t[285] = (t[331] & ~t[332]);
  assign t[286] = (t[333] & ~t[334]);
  assign t[287] = (t[335] & ~t[336]);
  assign t[288] = (t[337] & ~t[338]);
  assign t[289] = (t[339] & ~t[340]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[341] & ~t[342]);
  assign t[291] = (t[343] & ~t[344]);
  assign t[292] = (t[345] & ~t[346]);
  assign t[293] = t[347] ^ x[4];
  assign t[294] = t[348] ^ x[3];
  assign t[295] = t[349] ^ x[9];
  assign t[296] = t[350] ^ x[8];
  assign t[297] = t[351] ^ x[12];
  assign t[298] = t[352] ^ x[11];
  assign t[299] = t[353] ^ x[15];
  assign t[29] = ~(t[213]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[14];
  assign t[301] = t[355] ^ x[18];
  assign t[302] = t[356] ^ x[17];
  assign t[303] = t[357] ^ x[21];
  assign t[304] = t[358] ^ x[20];
  assign t[305] = t[359] ^ x[24];
  assign t[306] = t[360] ^ x[23];
  assign t[307] = t[361] ^ x[27];
  assign t[308] = t[362] ^ x[26];
  assign t[309] = t[363] ^ x[30];
  assign t[30] = ~(t[214]);
  assign t[310] = t[364] ^ x[29];
  assign t[311] = t[365] ^ x[33];
  assign t[312] = t[366] ^ x[32];
  assign t[313] = t[367] ^ x[36];
  assign t[314] = t[368] ^ x[35];
  assign t[315] = t[369] ^ x[39];
  assign t[316] = t[370] ^ x[38];
  assign t[317] = t[371] ^ x[42];
  assign t[318] = t[372] ^ x[41];
  assign t[319] = t[373] ^ x[45];
  assign t[31] = ~(t[215]);
  assign t[320] = t[374] ^ x[44];
  assign t[321] = t[375] ^ x[48];
  assign t[322] = t[376] ^ x[47];
  assign t[323] = t[377] ^ x[51];
  assign t[324] = t[378] ^ x[50];
  assign t[325] = t[379] ^ x[54];
  assign t[326] = t[380] ^ x[53];
  assign t[327] = t[381] ^ x[57];
  assign t[328] = t[382] ^ x[56];
  assign t[329] = t[383] ^ x[60];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[59];
  assign t[331] = t[385] ^ x[63];
  assign t[332] = t[386] ^ x[62];
  assign t[333] = t[387] ^ x[66];
  assign t[334] = t[388] ^ x[65];
  assign t[335] = t[389] ^ x[71];
  assign t[336] = t[390] ^ x[70];
  assign t[337] = t[391] ^ x[74];
  assign t[338] = t[392] ^ x[73];
  assign t[339] = t[393] ^ x[85];
  assign t[33] = t[51] ^ t[52];
  assign t[340] = t[394] ^ x[84];
  assign t[341] = t[395] ^ x[92];
  assign t[342] = t[396] ^ x[91];
  assign t[343] = t[397] ^ x[97];
  assign t[344] = t[398] ^ x[96];
  assign t[345] = t[399] ^ x[106];
  assign t[346] = t[400] ^ x[105];
  assign t[347] = (x[2]);
  assign t[348] = (x[2]);
  assign t[349] = (x[7]);
  assign t[34] = t[53] ^ t[54];
  assign t[350] = (x[7]);
  assign t[351] = (x[10]);
  assign t[352] = (x[10]);
  assign t[353] = (x[13]);
  assign t[354] = (x[13]);
  assign t[355] = (x[16]);
  assign t[356] = (x[16]);
  assign t[357] = (x[19]);
  assign t[358] = (x[19]);
  assign t[359] = (x[22]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[22]);
  assign t[361] = (x[25]);
  assign t[362] = (x[25]);
  assign t[363] = (x[28]);
  assign t[364] = (x[28]);
  assign t[365] = (x[31]);
  assign t[366] = (x[31]);
  assign t[367] = (x[34]);
  assign t[368] = (x[34]);
  assign t[369] = (x[37]);
  assign t[36] = t[57] ^ t[58];
  assign t[370] = (x[37]);
  assign t[371] = (x[40]);
  assign t[372] = (x[40]);
  assign t[373] = (x[43]);
  assign t[374] = (x[43]);
  assign t[375] = (x[46]);
  assign t[376] = (x[46]);
  assign t[377] = (x[49]);
  assign t[378] = (x[49]);
  assign t[379] = (x[52]);
  assign t[37] = t[59] ^ t[60];
  assign t[380] = (x[52]);
  assign t[381] = (x[55]);
  assign t[382] = (x[55]);
  assign t[383] = (x[58]);
  assign t[384] = (x[58]);
  assign t[385] = (x[61]);
  assign t[386] = (x[61]);
  assign t[387] = (x[64]);
  assign t[388] = (x[64]);
  assign t[389] = (x[69]);
  assign t[38] = ~(t[61] ^ t[62]);
  assign t[390] = (x[69]);
  assign t[391] = (x[72]);
  assign t[392] = (x[72]);
  assign t[393] = (x[83]);
  assign t[394] = (x[83]);
  assign t[395] = (x[90]);
  assign t[396] = (x[90]);
  assign t[397] = (x[95]);
  assign t[398] = (x[95]);
  assign t[399] = (x[104]);
  assign t[39] = ~(t[63] ^ t[64]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[400] = (x[104]);
  assign t[40] = t[65] ^ t[66];
  assign t[41] = t[67] ^ t[68];
  assign t[42] = t[69] ^ t[55];
  assign t[43] = ~(t[38] ^ t[70]);
  assign t[44] = t[11] ^ t[71];
  assign t[45] = ~(t[62] ^ t[41]);
  assign t[46] = ~(t[72] & t[73]);
  assign t[47] = t[216] | t[74];
  assign t[48] = ~(t[75]);
  assign t[49] = ~(t[217]);
  assign t[4] = t[8] ? t[9] : t[212];
  assign t[50] = ~(t[76] & t[218]);
  assign t[51] = t[77] ^ t[57];
  assign t[52] = t[78] & t[79];
  assign t[53] = t[80] ^ t[81];
  assign t[54] = t[82] & t[83];
  assign t[55] = t[84] ^ t[85];
  assign t[56] = t[86] ^ t[87];
  assign t[57] = t[88] ? t[89] : t[219];
  assign t[58] = t[90] ^ t[91];
  assign t[59] = ~t[92];
  assign t[5] = ~(t[10]);
  assign t[60] = t[93] ^ t[94];
  assign t[61] = ~(t[95] ^ t[96]);
  assign t[62] = t[97] ^ t[98];
  assign t[63] = t[99] ^ t[100];
  assign t[64] = ~(t[70] ^ t[41]);
  assign t[65] = t[101] ^ t[67];
  assign t[66] = t[102] ^ t[103];
  assign t[67] = t[218] ^ t[104];
  assign t[68] = t[102] ^ t[87];
  assign t[69] = t[105] ^ t[106];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[107] ^ t[108];
  assign t[71] = t[109] ^ t[94];
  assign t[72] = ~(t[74] & t[110]);
  assign t[73] = ~(t[220] ^ t[111]);
  assign t[74] = ~(t[112] & t[113]);
  assign t[75] = ~(t[47]);
  assign t[76] = ~(t[221]);
  assign t[77] = t[88] ? t[114] : t[222];
  assign t[78] = ~(t[115]);
  assign t[79] = t[88] ? t[116] : t[223];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[8] ? t[117] : t[224];
  assign t[81] = t[8] ? t[118] : t[225];
  assign t[82] = ~(t[53] ^ t[119]);
  assign t[83] = t[97] ^ t[120];
  assign t[84] = t[121] ^ t[59];
  assign t[85] = t[93] ^ t[122];
  assign t[86] = t[123] ^ t[101];
  assign t[87] = t[124] & t[125];
  assign t[88] = ~(t[15]);
  assign t[89] = t[219] ^ t[126];
  assign t[8] = ~(t[15]);
  assign t[90] = t[127] ^ t[52];
  assign t[91] = t[128] & t[129];
  assign t[92] = t[27] ? t[130] : t[226];
  assign t[93] = t[131] ^ t[132];
  assign t[94] = t[133] & t[134];
  assign t[95] = t[40] ^ t[37];
  assign t[96] = t[135] ^ t[91];
  assign t[97] = t[81] ^ t[107];
  assign t[98] = t[119] ^ t[136];
  assign t[99] = t[137] ^ t[138];
  assign t[9] = t[212] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[141] ^ t[142];
  assign t[101] = t[28] ? x[50] : x[49];
  assign t[102] = t[28] ? x[52] : x[51];
  assign t[103] = t[220] ^ t[143];
  assign t[104] = ~(t[144] & t[145]);
  assign t[105] = t[146] ^ t[225];
  assign t[106] = ~(t[221]);
  assign t[107] = t[147] & t[146];
  assign t[108] = t[87] ^ t[127];
  assign t[109] = t[148] & t[149];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[132] ? t[150] : t[226];
  assign t[111] = t[112] ^ t[62];
  assign t[112] = t[151] ^ t[152];
  assign t[113] = t[153] & t[154];
  assign t[114] = t[27] ? t[155] : t[227];
  assign t[115] = t[156] ^ t[59];
  assign t[116] = t[127] ^ t[78];
  assign t[117] = t[115] ^ t[157];
  assign t[118] = t[158] ^ t[129];
  assign t[119] = t[159] & t[160];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[63] ^ t[161];
  assign t[121] = t[141] ^ t[98];
  assign t[122] = t[158] ^ t[124];
  assign t[123] = t[162] & t[163];
  assign t[124] = t[218] ^ t[164];
  assign t[125] = t[130] ^ t[119];
  assign t[126] = t[27] ? t[165] : t[228];
  assign t[127] = t[166];
  assign t[128] = t[27] ? t[167] : t[229];
  assign t[129] = t[211] ^ t[168];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[169] ^ t[123];
  assign t[131] = t[170] & t[171];
  assign t[132] = ~(t[15]);
  assign t[133] = t[223] ^ t[172];
  assign t[134] = t[224] ^ t[173];
  assign t[135] = t[132] ? t[174] : t[230];
  assign t[136] = t[28] ? x[72] : x[71];
  assign t[137] = ~(t[142]);
  assign t[138] = ~(t[42]);
  assign t[139] = ~(t[43]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[40] ^ t[42];
  assign t[141] = t[42] ^ t[63];
  assign t[142] = t[68] ^ t[43];
  assign t[143] = t[28] ? x[74] : x[73];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[175] | t[106]);
  assign t[146] = ~(t[231]);
  assign t[147] = ~(t[225]);
  assign t[148] = ~(t[108] ^ t[115]);
  assign t[149] = t[116] ^ t[89];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[226] ^ t[176];
  assign t[151] = t[177] & t[178];
  assign t[152] = t[179] & t[135];
  assign t[153] = ~(t[151] ^ t[180]);
  assign t[154] = t[181] ^ t[182];
  assign t[155] = t[227] ^ t[183];
  assign t[156] = t[184] & t[185];
  assign t[157] = t[186] & t[187];
  assign t[158] = t[8] ? t[188] : t[232];
  assign t[159] = ~(t[118] ^ t[130]);
  assign t[15] = ~(t[27]);
  assign t[160] = t[90] ^ t[163];
  assign t[161] = t[64] ^ t[26];
  assign t[162] = ~(t[129]);
  assign t[163] = t[212] ^ t[189];
  assign t[164] = t[8] ? t[190] : t[233];
  assign t[165] = t[228] ^ t[191];
  assign t[166] = t[27] ? t[192] : t[234];
  assign t[167] = t[229] ^ t[193];
  assign t[168] = t[27] ? t[194] : t[235];
  assign t[169] = t[195] & t[196];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[169] ^ t[197]);
  assign t[171] = t[122] ^ t[198];
  assign t[172] = t[199] ? x[91] : x[90];
  assign t[173] = t[199] ? x[93] : x[92];
  assign t[174] = t[230] ^ t[200];
  assign t[175] = ~(t[216]);
  assign t[176] = t[199] ? x[95] : x[94];
  assign t[177] = ~(t[182]);
  assign t[178] = ~(t[92]);
  assign t[179] = ~(t[93]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[76] ^ t[92];
  assign t[181] = t[92] ^ t[110];
  assign t[182] = t[135] ^ t[93];
  assign t[183] = t[72] ? x[97] : x[96];
  assign t[184] = ~(t[201]);
  assign t[185] = ~(t[87]);
  assign t[186] = ~(t[156] ^ t[202]);
  assign t[187] = t[58] ^ t[201];
  assign t[188] = t[232] ^ t[203];
  assign t[189] = t[8] ? t[204] : t[236];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[233] ^ t[205];
  assign t[191] = t[72] ? x[102] : x[101];
  assign t[192] = t[234] ^ t[206];
  assign t[193] = t[28] ? x[104] : x[103];
  assign t[194] = t[235] ^ t[207];
  assign t[195] = ~(t[198]);
  assign t[196] = ~(t[158]);
  assign t[197] = t[90] ^ t[158];
  assign t[198] = t[163] ^ t[129];
  assign t[199] = ~(t[48]);
  assign t[19] = ~(t[24] ^ t[33]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[199] ? x[106] : x[105];
  assign t[201] = t[89] ^ t[127];
  assign t[202] = t[116] ^ t[87];
  assign t[203] = t[72] ? x[108] : x[107];
  assign t[204] = t[236] ^ t[208];
  assign t[205] = t[72] ? x[110] : x[109];
  assign t[206] = t[209] ? x[112] : x[111];
  assign t[207] = t[209] ? x[114] : x[113];
  assign t[208] = t[209] ? x[116] : x[115];
  assign t[209] = ~(t[48]);
  assign t[20] = ~(t[34] ^ t[35]);
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[38] ^ t[14]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[9];
  assign t[239] = t[266] ^ x[12];
  assign t[23] = ~(t[38] ^ t[39]);
  assign t[240] = t[267] ^ x[15];
  assign t[241] = t[268] ^ x[18];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = t[40] ^ t[41];
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[55];
  assign t[253] = t[280] ^ x[58];
  assign t[254] = t[281] ^ x[61];
  assign t[255] = t[282] ^ x[64];
  assign t[256] = t[283] ^ x[67];
  assign t[257] = t[284] ^ x[70];
  assign t[258] = t[285] ^ x[77];
  assign t[259] = t[286] ^ x[80];
  assign t[25] = t[42] ^ t[43];
  assign t[260] = t[287] ^ x[83];
  assign t[261] = t[288] ^ x[86];
  assign t[262] = t[289] ^ x[89];
  assign t[263] = t[290] ^ x[100];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = t[44] & t[45];
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[9];
  assign t[294] = t[348] ^ x[8];
  assign t[295] = t[349] ^ x[12];
  assign t[296] = t[350] ^ x[11];
  assign t[297] = t[351] ^ x[15];
  assign t[298] = t[352] ^ x[14];
  assign t[299] = t[353] ^ x[18];
  assign t[29] = ~(t[211]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[17];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = ~(t[212]);
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[213]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[55];
  assign t[322] = t[376] ^ x[54];
  assign t[323] = t[377] ^ x[58];
  assign t[324] = t[378] ^ x[57];
  assign t[325] = t[379] ^ x[61];
  assign t[326] = t[380] ^ x[60];
  assign t[327] = t[381] ^ x[64];
  assign t[328] = t[382] ^ x[63];
  assign t[329] = t[383] ^ x[67];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[66];
  assign t[331] = t[385] ^ x[70];
  assign t[332] = t[386] ^ x[69];
  assign t[333] = t[387] ^ x[77];
  assign t[334] = t[388] ^ x[76];
  assign t[335] = t[389] ^ x[80];
  assign t[336] = t[390] ^ x[79];
  assign t[337] = t[391] ^ x[83];
  assign t[338] = t[392] ^ x[82];
  assign t[339] = t[393] ^ x[86];
  assign t[33] = ~(t[51] ^ t[52]);
  assign t[340] = t[394] ^ x[85];
  assign t[341] = t[395] ^ x[89];
  assign t[342] = t[396] ^ x[88];
  assign t[343] = t[397] ^ x[100];
  assign t[344] = t[398] ^ x[99];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[7]);
  assign t[348] = (x[7]);
  assign t[349] = (x[10]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[10]);
  assign t[351] = (x[13]);
  assign t[352] = (x[13]);
  assign t[353] = (x[16]);
  assign t[354] = (x[16]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = t[13] ^ t[55];
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[53]);
  assign t[376] = (x[53]);
  assign t[377] = (x[56]);
  assign t[378] = (x[56]);
  assign t[379] = (x[59]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[59]);
  assign t[381] = (x[62]);
  assign t[382] = (x[62]);
  assign t[383] = (x[65]);
  assign t[384] = (x[65]);
  assign t[385] = (x[68]);
  assign t[386] = (x[68]);
  assign t[387] = (x[75]);
  assign t[388] = (x[75]);
  assign t[389] = (x[78]);
  assign t[38] = t[60] ^ t[53];
  assign t[390] = (x[78]);
  assign t[391] = (x[81]);
  assign t[392] = (x[81]);
  assign t[393] = (x[84]);
  assign t[394] = (x[84]);
  assign t[395] = (x[87]);
  assign t[396] = (x[87]);
  assign t[397] = (x[98]);
  assign t[398] = (x[98]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[43] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[8] ? t[66] : t[214];
  assign t[43] = t[8] ? t[67] : t[215];
  assign t[44] = ~(t[25] ^ t[64]);
  assign t[45] = t[40] ^ t[68];
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = t[216] | t[71];
  assign t[48] = ~(t[72]);
  assign t[49] = ~(t[217]);
  assign t[4] = t[8] ? t[9] : t[210];
  assign t[50] = ~(t[73] & t[218]);
  assign t[51] = ~(t[74] ^ t[75]);
  assign t[52] = t[76] ^ t[77];
  assign t[53] = t[78] ^ t[79];
  assign t[54] = t[80] ^ t[81];
  assign t[55] = ~(t[82] ^ t[83]);
  assign t[56] = t[84] ^ t[33];
  assign t[57] = ~(t[85] ^ t[86]);
  assign t[58] = t[87] ^ t[78];
  assign t[59] = t[88] & t[89];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92] ^ t[93];
  assign t[62] = t[94] & t[95];
  assign t[63] = t[8] ? t[96] : t[219];
  assign t[64] = t[97] ^ t[98];
  assign t[65] = t[99] & t[100];
  assign t[66] = t[214] ^ t[101];
  assign t[67] = t[215] ^ t[102];
  assign t[68] = t[8] ? t[103] : t[220];
  assign t[69] = ~(t[71] & t[104]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[221] ^ t[105]);
  assign t[71] = ~(t[106] & t[107]);
  assign t[72] = ~(t[47]);
  assign t[73] = ~(t[222]);
  assign t[74] = t[108] ^ t[109];
  assign t[75] = t[110] ^ t[111];
  assign t[76] = t[93] ^ t[110];
  assign t[77] = t[112] ^ t[113];
  assign t[78] = ~t[114];
  assign t[79] = t[115] ^ t[109];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[116] ^ t[117];
  assign t[81] = t[118] ^ t[119];
  assign t[82] = t[52] ^ t[37];
  assign t[83] = ~(t[120] ^ t[86]);
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[122] ^ t[123];
  assign t[86] = t[124] ^ t[125];
  assign t[87] = ~t[126];
  assign t[88] = ~(t[127]);
  assign t[89] = t[128];
  assign t[8] = ~(t[15]);
  assign t[90] = t[129] ^ t[124];
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[132] ? t[133] : t[223];
  assign t[93] = t[132] ? t[134] : t[224];
  assign t[94] = ~(t[61] ^ t[112]);
  assign t[95] = t[76] ^ t[135];
  assign t[96] = t[219] ^ t[136];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[139] & t[68];
  assign t[99] = ~(t[97] ^ t[140]);
  assign t[9] = t[210] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind151(x, y);
 input [116:0] x;
 output y;

 wire [398:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[141] ^ t[142];
  assign t[101] = t[28] ? x[50] : x[49];
  assign t[102] = t[28] ? x[52] : x[51];
  assign t[103] = t[220] ^ t[143];
  assign t[104] = ~(t[144] & t[145]);
  assign t[105] = t[146] ^ t[225];
  assign t[106] = ~(t[221]);
  assign t[107] = t[147] & t[146];
  assign t[108] = t[87] ^ t[127];
  assign t[109] = t[148] & t[149];
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = t[132] ? t[150] : t[226];
  assign t[111] = t[112] ^ t[62];
  assign t[112] = t[151] ^ t[152];
  assign t[113] = t[153] & t[154];
  assign t[114] = t[27] ? t[155] : t[227];
  assign t[115] = t[156] ^ t[59];
  assign t[116] = t[127] ^ t[78];
  assign t[117] = t[115] ^ t[157];
  assign t[118] = t[158] ^ t[129];
  assign t[119] = t[159] & t[160];
  assign t[11] = ~(t[19] ^ t[20]);
  assign t[120] = t[63] ^ t[161];
  assign t[121] = t[141] ^ t[98];
  assign t[122] = t[158] ^ t[124];
  assign t[123] = t[162] & t[163];
  assign t[124] = t[218] ^ t[164];
  assign t[125] = t[130] ^ t[119];
  assign t[126] = t[27] ? t[165] : t[228];
  assign t[127] = t[166];
  assign t[128] = t[27] ? t[167] : t[229];
  assign t[129] = t[211] ^ t[168];
  assign t[12] = ~(t[21] ^ t[22]);
  assign t[130] = t[169] ^ t[123];
  assign t[131] = t[170] & t[171];
  assign t[132] = ~(t[15]);
  assign t[133] = t[223] ^ t[172];
  assign t[134] = t[224] ^ t[173];
  assign t[135] = t[132] ? t[174] : t[230];
  assign t[136] = t[28] ? x[72] : x[71];
  assign t[137] = ~(t[142]);
  assign t[138] = ~(t[42]);
  assign t[139] = ~(t[43]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[140] = t[40] ^ t[42];
  assign t[141] = t[42] ^ t[63];
  assign t[142] = t[68] ^ t[43];
  assign t[143] = t[28] ? x[74] : x[73];
  assign t[144] = ~(t[147] | t[146]);
  assign t[145] = ~(t[175] | t[106]);
  assign t[146] = ~(t[231]);
  assign t[147] = ~(t[225]);
  assign t[148] = ~(t[108] ^ t[115]);
  assign t[149] = t[116] ^ t[89];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[226] ^ t[176];
  assign t[151] = t[177] & t[178];
  assign t[152] = t[179] & t[135];
  assign t[153] = ~(t[151] ^ t[180]);
  assign t[154] = t[181] ^ t[182];
  assign t[155] = t[227] ^ t[183];
  assign t[156] = t[184] & t[185];
  assign t[157] = t[186] & t[187];
  assign t[158] = t[8] ? t[188] : t[232];
  assign t[159] = ~(t[118] ^ t[130]);
  assign t[15] = ~(t[27]);
  assign t[160] = t[90] ^ t[163];
  assign t[161] = t[64] ^ t[26];
  assign t[162] = ~(t[129]);
  assign t[163] = t[212] ^ t[189];
  assign t[164] = t[8] ? t[190] : t[233];
  assign t[165] = t[228] ^ t[191];
  assign t[166] = t[27] ? t[192] : t[234];
  assign t[167] = t[229] ^ t[193];
  assign t[168] = t[27] ? t[194] : t[235];
  assign t[169] = t[195] & t[196];
  assign t[16] = t[28] ? x[6] : x[5];
  assign t[170] = ~(t[169] ^ t[197]);
  assign t[171] = t[122] ^ t[198];
  assign t[172] = t[199] ? x[91] : x[90];
  assign t[173] = t[199] ? x[93] : x[92];
  assign t[174] = t[230] ^ t[200];
  assign t[175] = ~(t[216]);
  assign t[176] = t[199] ? x[95] : x[94];
  assign t[177] = ~(t[182]);
  assign t[178] = ~(t[92]);
  assign t[179] = ~(t[93]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[180] = t[76] ^ t[92];
  assign t[181] = t[92] ^ t[110];
  assign t[182] = t[135] ^ t[93];
  assign t[183] = t[72] ? x[97] : x[96];
  assign t[184] = ~(t[201]);
  assign t[185] = ~(t[87]);
  assign t[186] = ~(t[156] ^ t[202]);
  assign t[187] = t[58] ^ t[201];
  assign t[188] = t[232] ^ t[203];
  assign t[189] = t[8] ? t[204] : t[236];
  assign t[18] = ~(t[31] & t[32]);
  assign t[190] = t[233] ^ t[205];
  assign t[191] = t[72] ? x[102] : x[101];
  assign t[192] = t[234] ^ t[206];
  assign t[193] = t[28] ? x[104] : x[103];
  assign t[194] = t[235] ^ t[207];
  assign t[195] = ~(t[198]);
  assign t[196] = ~(t[158]);
  assign t[197] = t[90] ^ t[158];
  assign t[198] = t[163] ^ t[129];
  assign t[199] = ~(t[48]);
  assign t[19] = ~(t[24] ^ t[33]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[200] = t[199] ? x[106] : x[105];
  assign t[201] = t[89] ^ t[127];
  assign t[202] = t[116] ^ t[87];
  assign t[203] = t[72] ? x[108] : x[107];
  assign t[204] = t[236] ^ t[208];
  assign t[205] = t[72] ? x[110] : x[109];
  assign t[206] = t[209] ? x[112] : x[111];
  assign t[207] = t[209] ? x[114] : x[113];
  assign t[208] = t[209] ? x[116] : x[115];
  assign t[209] = ~(t[48]);
  assign t[20] = ~(t[34] ^ t[35]);
  assign t[210] = (t[237]);
  assign t[211] = (t[238]);
  assign t[212] = (t[239]);
  assign t[213] = (t[240]);
  assign t[214] = (t[241]);
  assign t[215] = (t[242]);
  assign t[216] = (t[243]);
  assign t[217] = (t[244]);
  assign t[218] = (t[245]);
  assign t[219] = (t[246]);
  assign t[21] = t[36] ^ t[37];
  assign t[220] = (t[247]);
  assign t[221] = (t[248]);
  assign t[222] = (t[249]);
  assign t[223] = (t[250]);
  assign t[224] = (t[251]);
  assign t[225] = (t[252]);
  assign t[226] = (t[253]);
  assign t[227] = (t[254]);
  assign t[228] = (t[255]);
  assign t[229] = (t[256]);
  assign t[22] = ~(t[38] ^ t[14]);
  assign t[230] = (t[257]);
  assign t[231] = (t[258]);
  assign t[232] = (t[259]);
  assign t[233] = (t[260]);
  assign t[234] = (t[261]);
  assign t[235] = (t[262]);
  assign t[236] = (t[263]);
  assign t[237] = t[264] ^ x[4];
  assign t[238] = t[265] ^ x[9];
  assign t[239] = t[266] ^ x[12];
  assign t[23] = ~(t[38] ^ t[39]);
  assign t[240] = t[267] ^ x[15];
  assign t[241] = t[268] ^ x[18];
  assign t[242] = t[269] ^ x[21];
  assign t[243] = t[270] ^ x[24];
  assign t[244] = t[271] ^ x[27];
  assign t[245] = t[272] ^ x[30];
  assign t[246] = t[273] ^ x[33];
  assign t[247] = t[274] ^ x[36];
  assign t[248] = t[275] ^ x[39];
  assign t[249] = t[276] ^ x[42];
  assign t[24] = t[40] ^ t[41];
  assign t[250] = t[277] ^ x[45];
  assign t[251] = t[278] ^ x[48];
  assign t[252] = t[279] ^ x[55];
  assign t[253] = t[280] ^ x[58];
  assign t[254] = t[281] ^ x[61];
  assign t[255] = t[282] ^ x[64];
  assign t[256] = t[283] ^ x[67];
  assign t[257] = t[284] ^ x[70];
  assign t[258] = t[285] ^ x[77];
  assign t[259] = t[286] ^ x[80];
  assign t[25] = t[42] ^ t[43];
  assign t[260] = t[287] ^ x[83];
  assign t[261] = t[288] ^ x[86];
  assign t[262] = t[289] ^ x[89];
  assign t[263] = t[290] ^ x[100];
  assign t[264] = (t[291] & ~t[292]);
  assign t[265] = (t[293] & ~t[294]);
  assign t[266] = (t[295] & ~t[296]);
  assign t[267] = (t[297] & ~t[298]);
  assign t[268] = (t[299] & ~t[300]);
  assign t[269] = (t[301] & ~t[302]);
  assign t[26] = t[44] & t[45];
  assign t[270] = (t[303] & ~t[304]);
  assign t[271] = (t[305] & ~t[306]);
  assign t[272] = (t[307] & ~t[308]);
  assign t[273] = (t[309] & ~t[310]);
  assign t[274] = (t[311] & ~t[312]);
  assign t[275] = (t[313] & ~t[314]);
  assign t[276] = (t[315] & ~t[316]);
  assign t[277] = (t[317] & ~t[318]);
  assign t[278] = (t[319] & ~t[320]);
  assign t[279] = (t[321] & ~t[322]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[280] = (t[323] & ~t[324]);
  assign t[281] = (t[325] & ~t[326]);
  assign t[282] = (t[327] & ~t[328]);
  assign t[283] = (t[329] & ~t[330]);
  assign t[284] = (t[331] & ~t[332]);
  assign t[285] = (t[333] & ~t[334]);
  assign t[286] = (t[335] & ~t[336]);
  assign t[287] = (t[337] & ~t[338]);
  assign t[288] = (t[339] & ~t[340]);
  assign t[289] = (t[341] & ~t[342]);
  assign t[28] = ~(t[48]);
  assign t[290] = (t[343] & ~t[344]);
  assign t[291] = t[345] ^ x[4];
  assign t[292] = t[346] ^ x[3];
  assign t[293] = t[347] ^ x[9];
  assign t[294] = t[348] ^ x[8];
  assign t[295] = t[349] ^ x[12];
  assign t[296] = t[350] ^ x[11];
  assign t[297] = t[351] ^ x[15];
  assign t[298] = t[352] ^ x[14];
  assign t[299] = t[353] ^ x[18];
  assign t[29] = ~(t[211]);
  assign t[2] = ~(t[5]);
  assign t[300] = t[354] ^ x[17];
  assign t[301] = t[355] ^ x[21];
  assign t[302] = t[356] ^ x[20];
  assign t[303] = t[357] ^ x[24];
  assign t[304] = t[358] ^ x[23];
  assign t[305] = t[359] ^ x[27];
  assign t[306] = t[360] ^ x[26];
  assign t[307] = t[361] ^ x[30];
  assign t[308] = t[362] ^ x[29];
  assign t[309] = t[363] ^ x[33];
  assign t[30] = ~(t[212]);
  assign t[310] = t[364] ^ x[32];
  assign t[311] = t[365] ^ x[36];
  assign t[312] = t[366] ^ x[35];
  assign t[313] = t[367] ^ x[39];
  assign t[314] = t[368] ^ x[38];
  assign t[315] = t[369] ^ x[42];
  assign t[316] = t[370] ^ x[41];
  assign t[317] = t[371] ^ x[45];
  assign t[318] = t[372] ^ x[44];
  assign t[319] = t[373] ^ x[48];
  assign t[31] = ~(t[213]);
  assign t[320] = t[374] ^ x[47];
  assign t[321] = t[375] ^ x[55];
  assign t[322] = t[376] ^ x[54];
  assign t[323] = t[377] ^ x[58];
  assign t[324] = t[378] ^ x[57];
  assign t[325] = t[379] ^ x[61];
  assign t[326] = t[380] ^ x[60];
  assign t[327] = t[381] ^ x[64];
  assign t[328] = t[382] ^ x[63];
  assign t[329] = t[383] ^ x[67];
  assign t[32] = ~(t[49] | t[50]);
  assign t[330] = t[384] ^ x[66];
  assign t[331] = t[385] ^ x[70];
  assign t[332] = t[386] ^ x[69];
  assign t[333] = t[387] ^ x[77];
  assign t[334] = t[388] ^ x[76];
  assign t[335] = t[389] ^ x[80];
  assign t[336] = t[390] ^ x[79];
  assign t[337] = t[391] ^ x[83];
  assign t[338] = t[392] ^ x[82];
  assign t[339] = t[393] ^ x[86];
  assign t[33] = ~(t[51] ^ t[52]);
  assign t[340] = t[394] ^ x[85];
  assign t[341] = t[395] ^ x[89];
  assign t[342] = t[396] ^ x[88];
  assign t[343] = t[397] ^ x[100];
  assign t[344] = t[398] ^ x[99];
  assign t[345] = (x[2]);
  assign t[346] = (x[2]);
  assign t[347] = (x[7]);
  assign t[348] = (x[7]);
  assign t[349] = (x[10]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[350] = (x[10]);
  assign t[351] = (x[13]);
  assign t[352] = (x[13]);
  assign t[353] = (x[16]);
  assign t[354] = (x[16]);
  assign t[355] = (x[19]);
  assign t[356] = (x[19]);
  assign t[357] = (x[22]);
  assign t[358] = (x[22]);
  assign t[359] = (x[25]);
  assign t[35] = t[13] ^ t[55];
  assign t[360] = (x[25]);
  assign t[361] = (x[28]);
  assign t[362] = (x[28]);
  assign t[363] = (x[31]);
  assign t[364] = (x[31]);
  assign t[365] = (x[34]);
  assign t[366] = (x[34]);
  assign t[367] = (x[37]);
  assign t[368] = (x[37]);
  assign t[369] = (x[40]);
  assign t[36] = ~(t[56] ^ t[57]);
  assign t[370] = (x[40]);
  assign t[371] = (x[43]);
  assign t[372] = (x[43]);
  assign t[373] = (x[46]);
  assign t[374] = (x[46]);
  assign t[375] = (x[53]);
  assign t[376] = (x[53]);
  assign t[377] = (x[56]);
  assign t[378] = (x[56]);
  assign t[379] = (x[59]);
  assign t[37] = t[58] ^ t[59];
  assign t[380] = (x[59]);
  assign t[381] = (x[62]);
  assign t[382] = (x[62]);
  assign t[383] = (x[65]);
  assign t[384] = (x[65]);
  assign t[385] = (x[68]);
  assign t[386] = (x[68]);
  assign t[387] = (x[75]);
  assign t[388] = (x[75]);
  assign t[389] = (x[78]);
  assign t[38] = t[60] ^ t[53];
  assign t[390] = (x[78]);
  assign t[391] = (x[81]);
  assign t[392] = (x[81]);
  assign t[393] = (x[84]);
  assign t[394] = (x[84]);
  assign t[395] = (x[87]);
  assign t[396] = (x[87]);
  assign t[397] = (x[98]);
  assign t[398] = (x[98]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[43] ^ t[63];
  assign t[41] = t[64] ^ t[65];
  assign t[42] = t[8] ? t[66] : t[214];
  assign t[43] = t[8] ? t[67] : t[215];
  assign t[44] = ~(t[25] ^ t[64]);
  assign t[45] = t[40] ^ t[68];
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = t[216] | t[71];
  assign t[48] = ~(t[72]);
  assign t[49] = ~(t[217]);
  assign t[4] = t[8] ? t[9] : t[210];
  assign t[50] = ~(t[73] & t[218]);
  assign t[51] = ~(t[74] ^ t[75]);
  assign t[52] = t[76] ^ t[77];
  assign t[53] = t[78] ^ t[79];
  assign t[54] = t[80] ^ t[81];
  assign t[55] = ~(t[82] ^ t[83]);
  assign t[56] = t[84] ^ t[33];
  assign t[57] = ~(t[85] ^ t[86]);
  assign t[58] = t[87] ^ t[78];
  assign t[59] = t[88] & t[89];
  assign t[5] = ~(t[10]);
  assign t[60] = t[90] ^ t[91];
  assign t[61] = t[92] ^ t[93];
  assign t[62] = t[94] & t[95];
  assign t[63] = t[8] ? t[96] : t[219];
  assign t[64] = t[97] ^ t[98];
  assign t[65] = t[99] & t[100];
  assign t[66] = t[214] ^ t[101];
  assign t[67] = t[215] ^ t[102];
  assign t[68] = t[8] ? t[103] : t[220];
  assign t[69] = ~(t[71] & t[104]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[221] ^ t[105]);
  assign t[71] = ~(t[106] & t[107]);
  assign t[72] = ~(t[47]);
  assign t[73] = ~(t[222]);
  assign t[74] = t[108] ^ t[109];
  assign t[75] = t[110] ^ t[111];
  assign t[76] = t[93] ^ t[110];
  assign t[77] = t[112] ^ t[113];
  assign t[78] = ~t[114];
  assign t[79] = t[115] ^ t[109];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[116] ^ t[117];
  assign t[81] = t[118] ^ t[119];
  assign t[82] = t[52] ^ t[37];
  assign t[83] = ~(t[120] ^ t[86]);
  assign t[84] = t[120] ^ t[121];
  assign t[85] = t[122] ^ t[123];
  assign t[86] = t[124] ^ t[125];
  assign t[87] = ~t[126];
  assign t[88] = ~(t[127]);
  assign t[89] = t[128];
  assign t[8] = ~(t[15]);
  assign t[90] = t[129] ^ t[124];
  assign t[91] = t[130] ^ t[131];
  assign t[92] = t[132] ? t[133] : t[223];
  assign t[93] = t[132] ? t[134] : t[224];
  assign t[94] = ~(t[61] ^ t[112]);
  assign t[95] = t[76] ^ t[135];
  assign t[96] = t[219] ^ t[136];
  assign t[97] = t[137] & t[138];
  assign t[98] = t[139] & t[68];
  assign t[99] = ~(t[97] ^ t[140]);
  assign t[9] = t[210] ^ t[16];
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [417:0] x;
 output [151:0] y;

  R2ind0 R2ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[2], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[2], x[1], x[0], x[3]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[2], x[1], x[0], x[3]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[12], x[11], x[10], x[18], x[17], x[16], x[3]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[12], x[11], x[10], x[18], x[17], x[16], x[3]}), .y(y[5]));
  R2ind6 R2ind6_inst(.x({x[15], x[14], x[13], x[3]}), .y(y[6]));
  R2ind7 R2ind7_inst(.x({x[15], x[14], x[13], x[3]}), .y(y[7]));
  R2ind8 R2ind8_inst(.x({x[21], x[20], x[19], x[3]}), .y(y[8]));
  R2ind9 R2ind9_inst(.x({x[21], x[20], x[19], x[3]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[6], x[5], x[4], x[3]}), .y(y[10]));
  R2ind11 R2ind11_inst(.x({x[6], x[5], x[4], x[3]}), .y(y[11]));
  R2ind12 R2ind12_inst(.x({x[9], x[8], x[7], x[3]}), .y(y[12]));
  R2ind13 R2ind13_inst(.x({x[9], x[8], x[7], x[3]}), .y(y[13]));
  R2ind14 R2ind14_inst(.x({x[18], x[17], x[16], x[3]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[18], x[17], x[16], x[3]}), .y(y[15]));
  R2ind16 R2ind16_inst(.x({x[3], x[24], x[23], x[22]}), .y(y[16]));
  R2ind17 R2ind17_inst(.x({x[3], x[24], x[23], x[22]}), .y(y[17]));
  R2ind18 R2ind18_inst(.x({x[27], x[26], x[25], x[3]}), .y(y[18]));
  R2ind19 R2ind19_inst(.x({x[27], x[26], x[25], x[3]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[30], x[29], x[28], x[3]}), .y(y[20]));
  R2ind21 R2ind21_inst(.x({x[30], x[29], x[28], x[3]}), .y(y[21]));
  R2ind22 R2ind22_inst(.x({x[33], x[32], x[31], x[3]}), .y(y[22]));
  R2ind23 R2ind23_inst(.x({x[33], x[32], x[31], x[3]}), .y(y[23]));
  R2ind24 R2ind24_inst(.x({x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[27], x[26], x[25], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[9], x[8], x[7], x[30], x[29], x[28], x[6], x[5], x[4], x[15], x[14], x[13], x[48], x[47], x[46], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[24], x[23], x[22], x[37], x[36], x[35], x[34], x[3]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[27], x[26], x[25], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[9], x[8], x[7], x[30], x[29], x[28], x[6], x[5], x[4], x[15], x[14], x[13], x[48], x[47], x[46], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[24], x[23], x[22], x[37], x[36], x[35], x[34], x[3]}), .y(y[25]));
  R2ind26 R2ind26_inst(.x({x[114], x[113], x[79], x[78], x[104], x[103], x[81], x[80], x[96], x[95], x[94], x[54], x[53], x[52], x[98], x[97], x[77], x[76], x[75], x[39], x[38], x[57], x[56], x[55], x[63], x[62], x[108], x[107], x[112], x[111], x[66], x[65], x[64], x[100], x[99], x[106], x[105], x[102], x[101], x[110], x[109], x[37], x[36], x[35], x[48], x[47], x[46], x[87], x[86], x[85], x[59], x[58], x[6], x[5], x[4], x[27], x[26], x[25], x[61], x[60], x[93], x[92], x[91], x[69], x[68], x[67], x[84], x[83], x[82], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[72], x[71], x[70], x[90], x[89], x[88], x[42], x[41], x[40], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[45], x[44], x[43], x[74], x[73], x[24], x[23], x[22], x[51], x[50], x[49], x[115], x[3]}), .y(y[26]));
  R2ind27 R2ind27_inst(.x({x[114], x[113], x[79], x[78], x[104], x[103], x[81], x[80], x[96], x[95], x[94], x[54], x[53], x[52], x[98], x[97], x[77], x[76], x[75], x[39], x[38], x[57], x[56], x[55], x[63], x[62], x[108], x[107], x[112], x[111], x[66], x[65], x[64], x[100], x[99], x[106], x[105], x[102], x[101], x[110], x[109], x[37], x[36], x[35], x[48], x[47], x[46], x[87], x[86], x[85], x[59], x[58], x[6], x[5], x[4], x[27], x[26], x[25], x[61], x[60], x[93], x[92], x[91], x[69], x[68], x[67], x[84], x[83], x[82], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[72], x[71], x[70], x[90], x[89], x[88], x[42], x[41], x[40], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[45], x[44], x[43], x[74], x[73], x[24], x[23], x[22], x[51], x[50], x[49], x[115], x[3]}), .y(y[27]));
  R2ind28 R2ind28_inst(.x({x[81], x[80], x[63], x[62], x[61], x[60], x[102], x[101], x[57], x[56], x[55], x[48], x[47], x[46], x[79], x[78], x[98], x[97], x[59], x[58], x[74], x[73], x[45], x[44], x[43], x[112], x[111], x[110], x[109], x[100], x[99], x[114], x[113], x[39], x[38], x[72], x[71], x[70], x[54], x[53], x[52], x[66], x[65], x[64], x[42], x[41], x[40], x[108], x[107], x[106], x[105], x[51], x[50], x[49], x[6], x[5], x[4], x[27], x[26], x[25], x[93], x[92], x[91], x[90], x[89], x[88], x[69], x[68], x[67], x[96], x[95], x[94], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[37], x[36], x[35], x[87], x[86], x[85], x[84], x[83], x[82], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[104], x[103], x[24], x[23], x[22], x[77], x[76], x[75], x[116], x[3]}), .y(y[28]));
  R2ind29 R2ind29_inst(.x({x[81], x[80], x[63], x[62], x[61], x[60], x[102], x[101], x[57], x[56], x[55], x[48], x[47], x[46], x[79], x[78], x[98], x[97], x[59], x[58], x[74], x[73], x[45], x[44], x[43], x[112], x[111], x[110], x[109], x[100], x[99], x[114], x[113], x[39], x[38], x[72], x[71], x[70], x[54], x[53], x[52], x[66], x[65], x[64], x[42], x[41], x[40], x[108], x[107], x[106], x[105], x[51], x[50], x[49], x[6], x[5], x[4], x[27], x[26], x[25], x[93], x[92], x[91], x[90], x[89], x[88], x[69], x[68], x[67], x[96], x[95], x[94], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[37], x[36], x[35], x[87], x[86], x[85], x[84], x[83], x[82], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[104], x[103], x[24], x[23], x[22], x[77], x[76], x[75], x[116], x[3]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[98], x[97], x[81], x[80], x[63], x[62], x[110], x[109], x[39], x[38], x[66], x[65], x[64], x[102], x[101], x[106], x[105], x[104], x[103], x[57], x[56], x[55], x[48], x[47], x[46], x[90], x[89], x[88], x[100], x[99], x[37], x[36], x[35], x[74], x[73], x[79], x[78], x[72], x[71], x[70], x[61], x[60], x[112], x[111], x[84], x[83], x[82], x[77], x[76], x[75], x[6], x[5], x[4], x[27], x[26], x[25], x[69], x[68], x[67], x[59], x[58], x[108], x[107], x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[93], x[92], x[91], x[9], x[8], x[7], x[30], x[29], x[28], x[15], x[14], x[13], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[42], x[41], x[40], x[87], x[86], x[85], x[114], x[113], x[24], x[23], x[22], x[96], x[95], x[94], x[117], x[3]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[98], x[97], x[81], x[80], x[63], x[62], x[110], x[109], x[39], x[38], x[66], x[65], x[64], x[102], x[101], x[106], x[105], x[104], x[103], x[57], x[56], x[55], x[48], x[47], x[46], x[90], x[89], x[88], x[100], x[99], x[37], x[36], x[35], x[74], x[73], x[79], x[78], x[72], x[71], x[70], x[61], x[60], x[112], x[111], x[84], x[83], x[82], x[77], x[76], x[75], x[6], x[5], x[4], x[27], x[26], x[25], x[69], x[68], x[67], x[59], x[58], x[108], x[107], x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[93], x[92], x[91], x[9], x[8], x[7], x[30], x[29], x[28], x[15], x[14], x[13], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[42], x[41], x[40], x[87], x[86], x[85], x[114], x[113], x[24], x[23], x[22], x[96], x[95], x[94], x[117], x[3]}), .y(y[31]));
  R2ind32 R2ind32_inst(.x({x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[27], x[26], x[25], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[30], x[29], x[28], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[6], x[5], x[4], x[33], x[32], x[31], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[15], x[14], x[13], x[24], x[23], x[22], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[9], x[8], x[7], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[3]}), .y(y[32]));
  R2ind33 R2ind33_inst(.x({x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[27], x[26], x[25], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[30], x[29], x[28], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[6], x[5], x[4], x[33], x[32], x[31], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[15], x[14], x[13], x[24], x[23], x[22], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[9], x[8], x[7], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[3]}), .y(y[33]));
  R2ind34 R2ind34_inst(.x({x[188], x[187], x[186], x[185], x[150], x[149], x[152], x[151], x[198], x[197], x[165], x[164], x[163], x[162], x[161], x[160], x[123], x[122], x[132], x[131], x[130], x[167], x[166], x[148], x[147], x[190], x[189], x[196], x[195], x[27], x[26], x[25], x[194], x[193], x[135], x[134], x[133], x[182], x[181], x[180], x[154], x[153], x[30], x[29], x[28], x[184], x[183], x[192], x[191], x[121], x[120], x[119], x[144], x[143], x[142], x[129], x[128], x[127], x[170], x[169], x[168], x[179], x[178], x[177], x[6], x[5], x[4], x[33], x[32], x[31], x[146], x[145], x[176], x[175], x[174], x[138], x[137], x[136], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[157], x[156], x[155], x[173], x[172], x[171], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[126], x[125], x[124], x[159], x[158], x[141], x[140], x[139], x[199], x[3]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[188], x[187], x[186], x[185], x[150], x[149], x[152], x[151], x[198], x[197], x[165], x[164], x[163], x[162], x[161], x[160], x[123], x[122], x[132], x[131], x[130], x[167], x[166], x[148], x[147], x[190], x[189], x[196], x[195], x[27], x[26], x[25], x[194], x[193], x[135], x[134], x[133], x[182], x[181], x[180], x[154], x[153], x[30], x[29], x[28], x[184], x[183], x[192], x[191], x[121], x[120], x[119], x[144], x[143], x[142], x[129], x[128], x[127], x[170], x[169], x[168], x[179], x[178], x[177], x[6], x[5], x[4], x[33], x[32], x[31], x[146], x[145], x[176], x[175], x[174], x[138], x[137], x[136], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[157], x[156], x[155], x[173], x[172], x[171], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[126], x[125], x[124], x[159], x[158], x[141], x[140], x[139], x[199], x[3]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[148], x[147], x[146], x[145], x[152], x[151], x[154], x[153], x[184], x[183], x[129], x[128], x[127], x[190], x[189], x[159], x[158], x[27], x[26], x[25], x[126], x[125], x[124], x[194], x[193], x[192], x[191], x[135], x[134], x[133], x[150], x[149], x[167], x[166], x[138], x[137], x[136], x[198], x[197], x[196], x[195], x[30], x[29], x[28], x[123], x[122], x[157], x[156], x[155], x[170], x[169], x[168], x[141], x[140], x[139], x[186], x[185], x[6], x[5], x[4], x[33], x[32], x[31], x[176], x[175], x[174], x[173], x[172], x[171], x[132], x[131], x[130], x[144], x[143], x[142], x[182], x[181], x[180], x[179], x[178], x[177], x[15], x[14], x[13], x[24], x[23], x[22], x[121], x[120], x[119], x[162], x[161], x[160], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[9], x[8], x[7], x[188], x[187], x[165], x[164], x[163], x[200], x[3]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[148], x[147], x[146], x[145], x[152], x[151], x[154], x[153], x[184], x[183], x[129], x[128], x[127], x[190], x[189], x[159], x[158], x[27], x[26], x[25], x[126], x[125], x[124], x[194], x[193], x[192], x[191], x[135], x[134], x[133], x[150], x[149], x[167], x[166], x[138], x[137], x[136], x[198], x[197], x[196], x[195], x[30], x[29], x[28], x[123], x[122], x[157], x[156], x[155], x[170], x[169], x[168], x[141], x[140], x[139], x[186], x[185], x[6], x[5], x[4], x[33], x[32], x[31], x[176], x[175], x[174], x[173], x[172], x[171], x[132], x[131], x[130], x[144], x[143], x[142], x[182], x[181], x[180], x[179], x[178], x[177], x[15], x[14], x[13], x[24], x[23], x[22], x[121], x[120], x[119], x[162], x[161], x[160], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[9], x[8], x[7], x[188], x[187], x[165], x[164], x[163], x[200], x[3]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[167], x[166], x[148], x[147], x[192], x[191], x[196], x[195], x[123], x[122], x[152], x[151], x[184], x[183], x[190], x[189], x[188], x[187], x[144], x[143], x[142], x[129], x[128], x[127], x[173], x[172], x[171], x[27], x[26], x[25], x[179], x[178], x[177], x[121], x[120], x[119], x[159], x[158], x[135], x[134], x[133], x[157], x[156], x[155], x[146], x[145], x[194], x[193], x[30], x[29], x[28], x[170], x[169], x[168], x[154], x[153], x[198], x[197], x[165], x[164], x[163], x[150], x[149], x[6], x[5], x[4], x[33], x[32], x[31], x[141], x[140], x[139], x[126], x[125], x[124], x[176], x[175], x[174], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[138], x[137], x[136], x[182], x[181], x[180], x[132], x[131], x[130], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[186], x[185], x[162], x[161], x[160], x[201], x[3]}), .y(y[38]));
  R2ind39 R2ind39_inst(.x({x[167], x[166], x[148], x[147], x[192], x[191], x[196], x[195], x[123], x[122], x[152], x[151], x[184], x[183], x[190], x[189], x[188], x[187], x[144], x[143], x[142], x[129], x[128], x[127], x[173], x[172], x[171], x[27], x[26], x[25], x[179], x[178], x[177], x[121], x[120], x[119], x[159], x[158], x[135], x[134], x[133], x[157], x[156], x[155], x[146], x[145], x[194], x[193], x[30], x[29], x[28], x[170], x[169], x[168], x[154], x[153], x[198], x[197], x[165], x[164], x[163], x[150], x[149], x[6], x[5], x[4], x[33], x[32], x[31], x[141], x[140], x[139], x[126], x[125], x[124], x[176], x[175], x[174], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[138], x[137], x[136], x[182], x[181], x[180], x[132], x[131], x[130], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[186], x[185], x[162], x[161], x[160], x[201], x[3]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[27], x[26], x[25], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[30], x[29], x[28], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[6], x[5], x[4], x[33], x[32], x[31], x[228], x[227], x[226], x[9], x[8], x[7], x[24], x[23], x[22], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[15], x[14], x[13], x[207], x[206], x[205], x[204], x[203], x[202], x[3]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[27], x[26], x[25], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[30], x[29], x[28], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[6], x[5], x[4], x[33], x[32], x[31], x[228], x[227], x[226], x[9], x[8], x[7], x[24], x[23], x[22], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[15], x[14], x[13], x[207], x[206], x[205], x[204], x[203], x[202], x[3]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[270], x[269], x[237], x[236], x[259], x[258], x[239], x[238], x[278], x[277], x[282], x[281], x[246], x[245], x[244], x[216], x[215], x[214], x[248], x[247], x[235], x[234], x[274], x[273], x[27], x[26], x[25], x[276], x[275], x[280], x[279], x[233], x[232], x[231], x[207], x[206], x[219], x[218], x[217], x[262], x[261], x[260], x[272], x[271], x[241], x[240], x[30], x[29], x[28], x[243], x[242], x[268], x[267], x[266], x[228], x[227], x[226], x[213], x[212], x[211], x[254], x[253], x[252], x[33], x[32], x[31], x[257], x[256], x[255], x[265], x[264], x[263], x[205], x[204], x[203], x[6], x[5], x[4], x[251], x[250], x[249], x[222], x[221], x[220], x[9], x[8], x[7], x[24], x[23], x[22], x[225], x[224], x[223], x[15], x[14], x[13], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[230], x[229], x[210], x[209], x[208], x[283], x[3]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[270], x[269], x[237], x[236], x[259], x[258], x[239], x[238], x[278], x[277], x[282], x[281], x[246], x[245], x[244], x[216], x[215], x[214], x[248], x[247], x[235], x[234], x[274], x[273], x[27], x[26], x[25], x[276], x[275], x[280], x[279], x[233], x[232], x[231], x[207], x[206], x[219], x[218], x[217], x[262], x[261], x[260], x[272], x[271], x[241], x[240], x[30], x[29], x[28], x[243], x[242], x[268], x[267], x[266], x[228], x[227], x[226], x[213], x[212], x[211], x[254], x[253], x[252], x[33], x[32], x[31], x[257], x[256], x[255], x[265], x[264], x[263], x[205], x[204], x[203], x[6], x[5], x[4], x[251], x[250], x[249], x[222], x[221], x[220], x[9], x[8], x[7], x[24], x[23], x[22], x[225], x[224], x[223], x[15], x[14], x[13], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[230], x[229], x[210], x[209], x[208], x[283], x[3]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[243], x[242], x[235], x[234], x[276], x[275], x[239], x[238], x[241], x[240], x[225], x[224], x[223], x[282], x[281], x[280], x[279], x[213], x[212], x[211], x[274], x[273], x[27], x[26], x[25], x[257], x[256], x[255], x[219], x[218], x[217], x[237], x[236], x[248], x[247], x[222], x[221], x[220], x[278], x[277], x[230], x[229], x[30], x[29], x[28], x[268], x[267], x[266], x[265], x[264], x[263], x[254], x[253], x[252], x[272], x[271], x[270], x[269], x[33], x[32], x[31], x[207], x[206], x[216], x[215], x[214], x[228], x[227], x[226], x[6], x[5], x[4], x[262], x[261], x[260], x[210], x[209], x[208], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[251], x[250], x[249], x[246], x[245], x[244], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[205], x[204], x[203], x[259], x[258], x[233], x[232], x[231], x[284], x[3]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[243], x[242], x[235], x[234], x[276], x[275], x[239], x[238], x[241], x[240], x[225], x[224], x[223], x[282], x[281], x[280], x[279], x[213], x[212], x[211], x[274], x[273], x[27], x[26], x[25], x[257], x[256], x[255], x[219], x[218], x[217], x[237], x[236], x[248], x[247], x[222], x[221], x[220], x[278], x[277], x[230], x[229], x[30], x[29], x[28], x[268], x[267], x[266], x[265], x[264], x[263], x[254], x[253], x[252], x[272], x[271], x[270], x[269], x[33], x[32], x[31], x[207], x[206], x[216], x[215], x[214], x[228], x[227], x[226], x[6], x[5], x[4], x[262], x[261], x[260], x[210], x[209], x[208], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[251], x[250], x[249], x[246], x[245], x[244], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[205], x[204], x[203], x[259], x[258], x[233], x[232], x[231], x[284], x[3]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[280], x[279], x[248], x[247], x[235], x[234], x[276], x[275], x[239], x[238], x[265], x[264], x[263], x[274], x[273], x[272], x[271], x[207], x[206], x[228], x[227], x[226], x[213], x[212], x[211], x[257], x[256], x[255], x[243], x[242], x[282], x[281], x[27], x[26], x[25], x[259], x[258], x[219], x[218], x[217], x[30], x[29], x[28], x[254], x[253], x[252], x[251], x[250], x[249], x[241], x[240], x[278], x[277], x[205], x[204], x[203], x[230], x[229], x[237], x[236], x[225], x[224], x[223], x[268], x[267], x[266], x[33], x[32], x[31], x[6], x[5], x[4], x[233], x[232], x[231], x[9], x[8], x[7], x[24], x[23], x[22], x[222], x[221], x[220], x[262], x[261], x[260], x[210], x[209], x[208], x[216], x[215], x[214], x[12], x[11], x[10], x[18], x[17], x[16], x[15], x[14], x[13], x[21], x[20], x[19], x[270], x[269], x[246], x[245], x[244], x[285], x[3]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[280], x[279], x[248], x[247], x[235], x[234], x[276], x[275], x[239], x[238], x[265], x[264], x[263], x[274], x[273], x[272], x[271], x[207], x[206], x[228], x[227], x[226], x[213], x[212], x[211], x[257], x[256], x[255], x[243], x[242], x[282], x[281], x[27], x[26], x[25], x[259], x[258], x[219], x[218], x[217], x[30], x[29], x[28], x[254], x[253], x[252], x[251], x[250], x[249], x[241], x[240], x[278], x[277], x[205], x[204], x[203], x[230], x[229], x[237], x[236], x[225], x[224], x[223], x[268], x[267], x[266], x[33], x[32], x[31], x[6], x[5], x[4], x[233], x[232], x[231], x[9], x[8], x[7], x[24], x[23], x[22], x[222], x[221], x[220], x[262], x[261], x[260], x[210], x[209], x[208], x[216], x[215], x[214], x[12], x[11], x[10], x[18], x[17], x[16], x[15], x[14], x[13], x[21], x[20], x[19], x[270], x[269], x[246], x[245], x[244], x[285], x[3]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[366], x[365], x[364], x[363], x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[352], x[351], x[350], x[349], x[348], x[347], x[346], x[27], x[26], x[25], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[336], x[335], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[30], x[29], x[28], x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[6], x[5], x[4], x[33], x[32], x[31], x[311], x[310], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[15], x[14], x[13], x[24], x[23], x[22], x[300], x[299], x[298], x[297], x[296], x[295], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[9], x[8], x[7], x[294], x[293], x[292], x[291], x[290], x[289], x[288], x[287], x[286], x[3]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[366], x[365], x[364], x[363], x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[352], x[351], x[350], x[349], x[348], x[347], x[346], x[27], x[26], x[25], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[336], x[335], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[30], x[29], x[28], x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[6], x[5], x[4], x[33], x[32], x[31], x[311], x[310], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[15], x[14], x[13], x[24], x[23], x[22], x[300], x[299], x[298], x[297], x[296], x[295], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[9], x[8], x[7], x[294], x[293], x[292], x[291], x[290], x[289], x[288], x[287], x[286], x[3]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[331], x[330], x[356], x[355], x[333], x[332], x[347], x[346], x[306], x[305], x[304], x[349], x[348], x[329], x[328], x[366], x[365], x[327], x[326], x[325], x[309], x[308], x[307], x[360], x[359], x[27], x[26], x[25], x[364], x[363], x[316], x[315], x[314], x[291], x[290], x[319], x[318], x[317], x[303], x[302], x[301], x[351], x[350], x[358], x[357], x[30], x[29], x[28], x[324], x[323], x[354], x[353], x[352], x[362], x[361], x[339], x[338], x[337], x[311], x[310], x[6], x[5], x[4], x[33], x[32], x[31], x[345], x[344], x[343], x[289], x[288], x[287], x[322], x[321], x[320], x[336], x[335], x[334], x[15], x[14], x[13], x[24], x[23], x[22], x[300], x[299], x[298], x[342], x[341], x[340], x[294], x[293], x[292], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[9], x[8], x[7], x[313], x[312], x[297], x[296], x[295], x[367], x[3]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[331], x[330], x[356], x[355], x[333], x[332], x[347], x[346], x[306], x[305], x[304], x[349], x[348], x[329], x[328], x[366], x[365], x[327], x[326], x[325], x[309], x[308], x[307], x[360], x[359], x[27], x[26], x[25], x[364], x[363], x[316], x[315], x[314], x[291], x[290], x[319], x[318], x[317], x[303], x[302], x[301], x[351], x[350], x[358], x[357], x[30], x[29], x[28], x[324], x[323], x[354], x[353], x[352], x[362], x[361], x[339], x[338], x[337], x[311], x[310], x[6], x[5], x[4], x[33], x[32], x[31], x[345], x[344], x[343], x[289], x[288], x[287], x[322], x[321], x[320], x[336], x[335], x[334], x[15], x[14], x[13], x[24], x[23], x[22], x[300], x[299], x[298], x[342], x[341], x[340], x[294], x[293], x[292], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[9], x[8], x[7], x[313], x[312], x[297], x[296], x[295], x[367], x[3]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[329], x[328], x[324], x[323], x[333], x[332], x[364], x[363], x[303], x[302], x[301], x[300], x[299], x[298], x[366], x[365], x[309], x[308], x[307], x[331], x[330], x[349], x[348], x[311], x[310], x[27], x[26], x[25], x[345], x[344], x[343], x[362], x[361], x[351], x[350], x[313], x[312], x[30], x[29], x[28], x[354], x[353], x[352], x[306], x[305], x[304], x[319], x[318], x[317], x[294], x[293], x[292], x[360], x[359], x[358], x[357], x[356], x[355], x[6], x[5], x[4], x[33], x[32], x[31], x[291], x[290], x[342], x[341], x[340], x[322], x[321], x[320], x[297], x[296], x[295], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[339], x[338], x[337], x[336], x[335], x[334], x[327], x[326], x[325], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[289], x[288], x[287], x[347], x[346], x[316], x[315], x[314], x[368], x[3]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[329], x[328], x[324], x[323], x[333], x[332], x[364], x[363], x[303], x[302], x[301], x[300], x[299], x[298], x[366], x[365], x[309], x[308], x[307], x[331], x[330], x[349], x[348], x[311], x[310], x[27], x[26], x[25], x[345], x[344], x[343], x[362], x[361], x[351], x[350], x[313], x[312], x[30], x[29], x[28], x[354], x[353], x[352], x[306], x[305], x[304], x[319], x[318], x[317], x[294], x[293], x[292], x[360], x[359], x[358], x[357], x[356], x[355], x[6], x[5], x[4], x[33], x[32], x[31], x[291], x[290], x[342], x[341], x[340], x[322], x[321], x[320], x[297], x[296], x[295], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[339], x[338], x[337], x[336], x[335], x[334], x[327], x[326], x[325], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[289], x[288], x[287], x[347], x[346], x[316], x[315], x[314], x[368], x[3]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[349], x[348], x[329], x[328], x[333], x[332], x[364], x[363], x[362], x[361], x[319], x[318], x[317], x[303], x[302], x[301], x[358], x[357], x[291], x[290], x[309], x[308], x[307], x[345], x[344], x[343], x[342], x[341], x[340], x[324], x[323], x[366], x[365], x[27], x[26], x[25], x[351], x[350], x[347], x[346], x[331], x[330], x[30], x[29], x[28], x[336], x[335], x[334], x[289], x[288], x[287], x[313], x[312], x[300], x[299], x[298], x[354], x[353], x[352], x[6], x[5], x[4], x[33], x[32], x[31], x[322], x[321], x[320], x[311], x[310], x[360], x[359], x[316], x[315], x[314], x[306], x[305], x[304], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[297], x[296], x[295], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[294], x[293], x[292], x[339], x[338], x[337], x[356], x[355], x[327], x[326], x[325], x[369], x[3]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[349], x[348], x[329], x[328], x[333], x[332], x[364], x[363], x[362], x[361], x[319], x[318], x[317], x[303], x[302], x[301], x[358], x[357], x[291], x[290], x[309], x[308], x[307], x[345], x[344], x[343], x[342], x[341], x[340], x[324], x[323], x[366], x[365], x[27], x[26], x[25], x[351], x[350], x[347], x[346], x[331], x[330], x[30], x[29], x[28], x[336], x[335], x[334], x[289], x[288], x[287], x[313], x[312], x[300], x[299], x[298], x[354], x[353], x[352], x[6], x[5], x[4], x[33], x[32], x[31], x[322], x[321], x[320], x[311], x[310], x[360], x[359], x[316], x[315], x[314], x[306], x[305], x[304], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[297], x[296], x[295], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[294], x[293], x[292], x[339], x[338], x[337], x[356], x[355], x[327], x[326], x[325], x[369], x[3]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[39], x[38], x[104], x[103], x[106], x[105], x[37], x[36], x[35], x[74], x[73], x[114], x[113], x[81], x[80], x[63], x[62], x[100], x[99], x[77], x[76], x[75], x[84], x[83], x[82], x[108], x[107], x[51], x[50], x[49], x[96], x[95], x[94], x[57], x[56], x[55], x[48], x[47], x[46], x[79], x[78], x[98], x[97], x[112], x[111], x[69], x[68], x[67], x[102], x[101], x[61], x[60], x[110], x[109], x[6], x[5], x[4], x[27], x[26], x[25], x[59], x[58], x[87], x[86], x[85], x[54], x[53], x[52], x[66], x[65], x[64], x[93], x[92], x[91], x[9], x[8], x[7], x[30], x[29], x[28], x[15], x[14], x[13], x[72], x[71], x[70], x[45], x[44], x[43], x[90], x[89], x[88], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[42], x[41], x[40], x[331], x[330], x[24], x[23], x[22], x[306], x[305], x[304], x[370], x[3]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[39], x[38], x[104], x[103], x[106], x[105], x[37], x[36], x[35], x[74], x[73], x[114], x[113], x[81], x[80], x[63], x[62], x[100], x[99], x[77], x[76], x[75], x[84], x[83], x[82], x[108], x[107], x[51], x[50], x[49], x[96], x[95], x[94], x[57], x[56], x[55], x[48], x[47], x[46], x[79], x[78], x[98], x[97], x[112], x[111], x[69], x[68], x[67], x[102], x[101], x[61], x[60], x[110], x[109], x[6], x[5], x[4], x[27], x[26], x[25], x[59], x[58], x[87], x[86], x[85], x[54], x[53], x[52], x[66], x[65], x[64], x[93], x[92], x[91], x[9], x[8], x[7], x[30], x[29], x[28], x[15], x[14], x[13], x[72], x[71], x[70], x[45], x[44], x[43], x[90], x[89], x[88], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[42], x[41], x[40], x[331], x[330], x[24], x[23], x[22], x[306], x[305], x[304], x[370], x[3]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[104], x[103], x[39], x[38], x[74], x[73], x[114], x[113], x[81], x[80], x[63], x[62], x[77], x[76], x[75], x[102], x[101], x[98], x[97], x[61], x[60], x[37], x[36], x[35], x[51], x[50], x[49], x[96], x[95], x[94], x[112], x[111], x[110], x[109], x[57], x[56], x[55], x[48], x[47], x[46], x[72], x[71], x[70], x[66], x[65], x[64], x[79], x[78], x[108], x[107], x[45], x[44], x[43], x[93], x[92], x[91], x[90], x[89], x[88], x[100], x[99], x[106], x[105], x[6], x[5], x[4], x[27], x[26], x[25], x[54], x[53], x[52], x[87], x[86], x[85], x[59], x[58], x[9], x[8], x[7], x[30], x[29], x[28], x[15], x[14], x[13], x[69], x[68], x[67], x[84], x[83], x[82], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[42], x[41], x[40], x[349], x[348], x[24], x[23], x[22], x[319], x[318], x[317], x[371], x[3]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[104], x[103], x[39], x[38], x[74], x[73], x[114], x[113], x[81], x[80], x[63], x[62], x[77], x[76], x[75], x[102], x[101], x[98], x[97], x[61], x[60], x[37], x[36], x[35], x[51], x[50], x[49], x[96], x[95], x[94], x[112], x[111], x[110], x[109], x[57], x[56], x[55], x[48], x[47], x[46], x[72], x[71], x[70], x[66], x[65], x[64], x[79], x[78], x[108], x[107], x[45], x[44], x[43], x[93], x[92], x[91], x[90], x[89], x[88], x[100], x[99], x[106], x[105], x[6], x[5], x[4], x[27], x[26], x[25], x[54], x[53], x[52], x[87], x[86], x[85], x[59], x[58], x[9], x[8], x[7], x[30], x[29], x[28], x[15], x[14], x[13], x[69], x[68], x[67], x[84], x[83], x[82], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[42], x[41], x[40], x[349], x[348], x[24], x[23], x[22], x[319], x[318], x[317], x[371], x[3]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[114], x[113], x[104], x[103], x[96], x[95], x[94], x[77], x[76], x[75], x[74], x[73], x[39], x[38], x[98], x[97], x[102], x[101], x[110], x[109], x[51], x[50], x[49], x[37], x[36], x[35], x[59], x[58], x[100], x[99], x[112], x[111], x[81], x[80], x[79], x[78], x[61], x[60], x[108], x[107], x[106], x[105], x[66], x[65], x[64], x[63], x[62], x[72], x[71], x[70], x[90], x[89], x[88], x[42], x[41], x[40], x[27], x[26], x[25], x[69], x[68], x[67], x[93], x[92], x[91], x[57], x[56], x[55], x[54], x[53], x[52], x[45], x[44], x[43], x[9], x[8], x[7], x[30], x[29], x[28], x[87], x[86], x[85], x[84], x[83], x[82], x[6], x[5], x[4], x[15], x[14], x[13], x[48], x[47], x[46], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[333], x[332], x[24], x[23], x[22], x[309], x[308], x[307], x[372], x[3]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[114], x[113], x[104], x[103], x[96], x[95], x[94], x[77], x[76], x[75], x[74], x[73], x[39], x[38], x[98], x[97], x[102], x[101], x[110], x[109], x[51], x[50], x[49], x[37], x[36], x[35], x[59], x[58], x[100], x[99], x[112], x[111], x[81], x[80], x[79], x[78], x[61], x[60], x[108], x[107], x[106], x[105], x[66], x[65], x[64], x[63], x[62], x[72], x[71], x[70], x[90], x[89], x[88], x[42], x[41], x[40], x[27], x[26], x[25], x[69], x[68], x[67], x[93], x[92], x[91], x[57], x[56], x[55], x[54], x[53], x[52], x[45], x[44], x[43], x[9], x[8], x[7], x[30], x[29], x[28], x[87], x[86], x[85], x[84], x[83], x[82], x[6], x[5], x[4], x[15], x[14], x[13], x[48], x[47], x[46], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[333], x[332], x[24], x[23], x[22], x[309], x[308], x[307], x[372], x[3]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[74], x[73], x[79], x[78], x[112], x[111], x[110], x[109], x[104], x[103], x[114], x[113], x[102], x[101], x[100], x[99], x[81], x[80], x[39], x[38], x[106], x[105], x[51], x[50], x[49], x[54], x[53], x[52], x[98], x[97], x[93], x[92], x[91], x[90], x[89], x[88], x[77], x[76], x[75], x[96], x[95], x[94], x[72], x[71], x[70], x[69], x[68], x[67], x[59], x[58], x[108], x[107], x[57], x[56], x[55], x[63], x[62], x[37], x[36], x[35], x[84], x[83], x[82], x[27], x[26], x[25], x[61], x[60], x[6], x[5], x[4], x[66], x[65], x[64], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[42], x[41], x[40], x[87], x[86], x[85], x[48], x[47], x[46], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[45], x[44], x[43], x[329], x[328], x[24], x[23], x[22], x[303], x[302], x[301], x[373], x[3]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[74], x[73], x[79], x[78], x[112], x[111], x[110], x[109], x[104], x[103], x[114], x[113], x[102], x[101], x[100], x[99], x[81], x[80], x[39], x[38], x[106], x[105], x[51], x[50], x[49], x[54], x[53], x[52], x[98], x[97], x[93], x[92], x[91], x[90], x[89], x[88], x[77], x[76], x[75], x[96], x[95], x[94], x[72], x[71], x[70], x[69], x[68], x[67], x[59], x[58], x[108], x[107], x[57], x[56], x[55], x[63], x[62], x[37], x[36], x[35], x[84], x[83], x[82], x[27], x[26], x[25], x[61], x[60], x[6], x[5], x[4], x[66], x[65], x[64], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[42], x[41], x[40], x[87], x[86], x[85], x[48], x[47], x[46], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[45], x[44], x[43], x[329], x[328], x[24], x[23], x[22], x[303], x[302], x[301], x[373], x[3]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[123], x[122], x[196], x[195], x[188], x[187], x[190], x[189], x[121], x[120], x[119], x[159], x[158], x[148], x[147], x[179], x[178], x[177], x[198], x[197], x[165], x[164], x[163], x[186], x[185], x[152], x[151], x[27], x[26], x[25], x[170], x[169], x[168], x[141], x[140], x[139], x[129], x[128], x[127], x[194], x[193], x[30], x[29], x[28], x[154], x[153], x[182], x[181], x[180], x[162], x[161], x[160], x[135], x[134], x[133], x[150], x[149], x[167], x[166], x[184], x[183], x[146], x[145], x[192], x[191], x[6], x[5], x[4], x[33], x[32], x[31], x[176], x[175], x[174], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[138], x[137], x[136], x[132], x[131], x[130], x[144], x[143], x[142], x[157], x[156], x[155], x[126], x[125], x[124], x[173], x[172], x[171], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[79], x[78], x[54], x[53], x[52], x[374], x[3]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[123], x[122], x[196], x[195], x[188], x[187], x[190], x[189], x[121], x[120], x[119], x[159], x[158], x[148], x[147], x[179], x[178], x[177], x[198], x[197], x[165], x[164], x[163], x[186], x[185], x[152], x[151], x[27], x[26], x[25], x[170], x[169], x[168], x[141], x[140], x[139], x[129], x[128], x[127], x[194], x[193], x[30], x[29], x[28], x[154], x[153], x[182], x[181], x[180], x[162], x[161], x[160], x[135], x[134], x[133], x[150], x[149], x[167], x[166], x[184], x[183], x[146], x[145], x[192], x[191], x[6], x[5], x[4], x[33], x[32], x[31], x[176], x[175], x[174], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[138], x[137], x[136], x[132], x[131], x[130], x[144], x[143], x[142], x[157], x[156], x[155], x[126], x[125], x[124], x[173], x[172], x[171], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[79], x[78], x[54], x[53], x[52], x[374], x[3]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[188], x[187], x[123], x[122], x[159], x[158], x[148], x[147], x[165], x[164], x[163], x[186], x[185], x[184], x[183], x[152], x[151], x[146], x[145], x[121], x[120], x[119], x[141], x[140], x[139], x[194], x[193], x[192], x[191], x[167], x[166], x[198], x[197], x[129], x[128], x[127], x[162], x[161], x[160], x[157], x[156], x[155], x[135], x[134], x[133], x[190], x[189], x[196], x[195], x[126], x[125], x[124], x[176], x[175], x[174], x[173], x[172], x[171], x[144], x[143], x[142], x[150], x[149], x[182], x[181], x[180], x[154], x[153], x[6], x[5], x[4], x[27], x[26], x[25], x[170], x[169], x[168], x[179], x[178], x[177], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[132], x[131], x[130], x[138], x[137], x[136], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[98], x[97], x[24], x[23], x[22], x[66], x[65], x[64], x[375], x[3]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[188], x[187], x[123], x[122], x[159], x[158], x[148], x[147], x[165], x[164], x[163], x[186], x[185], x[184], x[183], x[152], x[151], x[146], x[145], x[121], x[120], x[119], x[141], x[140], x[139], x[194], x[193], x[192], x[191], x[167], x[166], x[198], x[197], x[129], x[128], x[127], x[162], x[161], x[160], x[157], x[156], x[155], x[135], x[134], x[133], x[190], x[189], x[196], x[195], x[126], x[125], x[124], x[176], x[175], x[174], x[173], x[172], x[171], x[144], x[143], x[142], x[150], x[149], x[182], x[181], x[180], x[154], x[153], x[6], x[5], x[4], x[27], x[26], x[25], x[170], x[169], x[168], x[179], x[178], x[177], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[132], x[131], x[130], x[138], x[137], x[136], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[98], x[97], x[24], x[23], x[22], x[66], x[65], x[64], x[375], x[3]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[188], x[187], x[186], x[185], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[123], x[122], x[154], x[153], x[190], x[189], x[184], x[183], x[192], x[191], x[141], x[140], x[139], x[121], x[120], x[119], x[198], x[197], x[196], x[195], x[194], x[193], x[167], x[166], x[146], x[145], x[138], x[137], x[136], x[170], x[169], x[168], x[152], x[151], x[150], x[149], x[148], x[147], x[157], x[156], x[155], x[173], x[172], x[171], x[6], x[5], x[4], x[27], x[26], x[25], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[144], x[143], x[142], x[126], x[125], x[124], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[81], x[80], x[24], x[23], x[22], x[57], x[56], x[55], x[376], x[3]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[188], x[187], x[186], x[185], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[123], x[122], x[154], x[153], x[190], x[189], x[184], x[183], x[192], x[191], x[141], x[140], x[139], x[121], x[120], x[119], x[198], x[197], x[196], x[195], x[194], x[193], x[167], x[166], x[146], x[145], x[138], x[137], x[136], x[170], x[169], x[168], x[152], x[151], x[150], x[149], x[148], x[147], x[157], x[156], x[155], x[173], x[172], x[171], x[6], x[5], x[4], x[27], x[26], x[25], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[144], x[143], x[142], x[126], x[125], x[124], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[81], x[80], x[24], x[23], x[22], x[57], x[56], x[55], x[376], x[3]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[159], x[158], x[190], x[189], x[194], x[193], x[192], x[191], x[196], x[195], x[188], x[187], x[184], x[183], x[150], x[149], x[123], x[122], x[141], x[140], x[139], x[186], x[185], x[170], x[169], x[168], x[154], x[153], x[198], x[197], x[152], x[151], x[176], x[175], x[174], x[173], x[172], x[171], x[179], x[178], x[177], x[165], x[164], x[163], x[157], x[156], x[155], x[132], x[131], x[130], x[167], x[166], x[148], x[147], x[121], x[120], x[119], x[162], x[161], x[160], x[6], x[5], x[4], x[27], x[26], x[25], x[146], x[145], x[138], x[137], x[136], x[182], x[181], x[180], x[135], x[134], x[133], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[144], x[143], x[142], x[129], x[128], x[127], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[126], x[125], x[124], x[63], x[62], x[24], x[23], x[22], x[48], x[47], x[46], x[377], x[3]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[159], x[158], x[190], x[189], x[194], x[193], x[192], x[191], x[196], x[195], x[188], x[187], x[184], x[183], x[150], x[149], x[123], x[122], x[141], x[140], x[139], x[186], x[185], x[170], x[169], x[168], x[154], x[153], x[198], x[197], x[152], x[151], x[176], x[175], x[174], x[173], x[172], x[171], x[179], x[178], x[177], x[165], x[164], x[163], x[157], x[156], x[155], x[132], x[131], x[130], x[167], x[166], x[148], x[147], x[121], x[120], x[119], x[162], x[161], x[160], x[6], x[5], x[4], x[27], x[26], x[25], x[146], x[145], x[138], x[137], x[136], x[182], x[181], x[180], x[135], x[134], x[133], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[144], x[143], x[142], x[129], x[128], x[127], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[126], x[125], x[124], x[63], x[62], x[24], x[23], x[22], x[48], x[47], x[46], x[377], x[3]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[207], x[206], x[274], x[273], x[272], x[271], x[259], x[258], x[235], x[234], x[278], x[277], x[205], x[204], x[203], x[230], x[229], x[270], x[269], x[239], x[238], x[282], x[281], x[254], x[253], x[252], x[251], x[250], x[249], x[233], x[232], x[231], x[213], x[212], x[211], x[276], x[275], x[243], x[242], x[280], x[279], x[241], x[240], x[262], x[261], x[260], x[210], x[209], x[208], x[246], x[245], x[244], x[219], x[218], x[217], x[237], x[236], x[248], x[247], x[268], x[267], x[266], x[6], x[5], x[4], x[27], x[26], x[25], x[257], x[256], x[255], x[225], x[224], x[223], x[265], x[264], x[263], x[9], x[8], x[7], x[30], x[29], x[28], x[222], x[221], x[220], x[216], x[215], x[214], x[228], x[227], x[226], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[15], x[14], x[13], x[150], x[149], x[24], x[23], x[22], x[132], x[131], x[130], x[378], x[3]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[207], x[206], x[274], x[273], x[272], x[271], x[259], x[258], x[235], x[234], x[278], x[277], x[205], x[204], x[203], x[230], x[229], x[270], x[269], x[239], x[238], x[282], x[281], x[254], x[253], x[252], x[251], x[250], x[249], x[233], x[232], x[231], x[213], x[212], x[211], x[276], x[275], x[243], x[242], x[280], x[279], x[241], x[240], x[262], x[261], x[260], x[210], x[209], x[208], x[246], x[245], x[244], x[219], x[218], x[217], x[237], x[236], x[248], x[247], x[268], x[267], x[266], x[6], x[5], x[4], x[27], x[26], x[25], x[257], x[256], x[255], x[225], x[224], x[223], x[265], x[264], x[263], x[9], x[8], x[7], x[30], x[29], x[28], x[222], x[221], x[220], x[216], x[215], x[214], x[228], x[227], x[226], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[15], x[14], x[13], x[150], x[149], x[24], x[23], x[22], x[132], x[131], x[130], x[378], x[3]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[259], x[258], x[276], x[275], x[243], x[242], x[235], x[234], x[207], x[206], x[230], x[229], x[270], x[269], x[282], x[281], x[280], x[279], x[239], x[238], x[233], x[232], x[231], x[257], x[256], x[255], x[248], x[247], x[278], x[277], x[225], x[224], x[223], x[213], x[212], x[211], x[205], x[204], x[203], x[210], x[209], x[208], x[246], x[245], x[244], x[268], x[267], x[266], x[265], x[264], x[263], x[219], x[218], x[217], x[274], x[273], x[228], x[227], x[226], x[237], x[236], x[262], x[261], x[260], x[272], x[271], x[241], x[240], x[27], x[26], x[25], x[254], x[253], x[252], x[9], x[8], x[7], x[30], x[29], x[28], x[216], x[215], x[214], x[6], x[5], x[4], x[251], x[250], x[249], x[222], x[221], x[220], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[15], x[14], x[13], x[167], x[166], x[24], x[23], x[22], x[144], x[143], x[142], x[379], x[3]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[259], x[258], x[276], x[275], x[243], x[242], x[235], x[234], x[207], x[206], x[230], x[229], x[270], x[269], x[282], x[281], x[280], x[279], x[239], x[238], x[233], x[232], x[231], x[257], x[256], x[255], x[248], x[247], x[278], x[277], x[225], x[224], x[223], x[213], x[212], x[211], x[205], x[204], x[203], x[210], x[209], x[208], x[246], x[245], x[244], x[268], x[267], x[266], x[265], x[264], x[263], x[219], x[218], x[217], x[274], x[273], x[228], x[227], x[226], x[237], x[236], x[262], x[261], x[260], x[272], x[271], x[241], x[240], x[27], x[26], x[25], x[254], x[253], x[252], x[9], x[8], x[7], x[30], x[29], x[28], x[216], x[215], x[214], x[6], x[5], x[4], x[251], x[250], x[249], x[222], x[221], x[220], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[15], x[14], x[13], x[167], x[166], x[24], x[23], x[22], x[144], x[143], x[142], x[379], x[3]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[270], x[269], x[259], x[258], x[246], x[245], x[244], x[276], x[275], x[280], x[279], x[233], x[232], x[231], x[230], x[229], x[207], x[206], x[241], x[240], x[274], x[273], x[282], x[281], x[243], x[242], x[278], x[277], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[210], x[209], x[208], x[205], x[204], x[203], x[222], x[221], x[220], x[254], x[253], x[252], x[272], x[271], x[268], x[267], x[266], x[239], x[238], x[237], x[236], x[235], x[234], x[225], x[224], x[223], x[27], x[26], x[25], x[6], x[5], x[4], x[262], x[261], x[260], x[228], x[227], x[226], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[251], x[250], x[249], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[152], x[151], x[24], x[23], x[22], x[135], x[134], x[133], x[380], x[3]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[270], x[269], x[259], x[258], x[246], x[245], x[244], x[276], x[275], x[280], x[279], x[233], x[232], x[231], x[230], x[229], x[207], x[206], x[241], x[240], x[274], x[273], x[282], x[281], x[243], x[242], x[278], x[277], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[210], x[209], x[208], x[205], x[204], x[203], x[222], x[221], x[220], x[254], x[253], x[252], x[272], x[271], x[268], x[267], x[266], x[239], x[238], x[237], x[236], x[235], x[234], x[225], x[224], x[223], x[27], x[26], x[25], x[6], x[5], x[4], x[262], x[261], x[260], x[228], x[227], x[226], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[251], x[250], x[249], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[152], x[151], x[24], x[23], x[22], x[135], x[134], x[133], x[380], x[3]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[282], x[281], x[280], x[279], x[276], x[275], x[274], x[273], x[230], x[229], x[237], x[236], x[268], x[267], x[266], x[265], x[264], x[263], x[272], x[271], x[259], x[258], x[270], x[269], x[257], x[256], x[255], x[254], x[253], x[252], x[241], x[240], x[278], x[277], x[239], x[238], x[207], x[206], x[210], x[209], x[208], x[243], x[242], x[216], x[215], x[214], x[248], x[247], x[235], x[234], x[251], x[250], x[249], x[233], x[232], x[231], x[246], x[245], x[244], x[6], x[5], x[4], x[27], x[26], x[25], x[222], x[221], x[220], x[262], x[261], x[260], x[219], x[218], x[217], x[205], x[204], x[203], x[9], x[8], x[7], x[30], x[29], x[28], x[225], x[224], x[223], x[15], x[14], x[13], x[228], x[227], x[226], x[213], x[212], x[211], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[148], x[147], x[24], x[23], x[22], x[129], x[128], x[127], x[381], x[3]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[282], x[281], x[280], x[279], x[276], x[275], x[274], x[273], x[230], x[229], x[237], x[236], x[268], x[267], x[266], x[265], x[264], x[263], x[272], x[271], x[259], x[258], x[270], x[269], x[257], x[256], x[255], x[254], x[253], x[252], x[241], x[240], x[278], x[277], x[239], x[238], x[207], x[206], x[210], x[209], x[208], x[243], x[242], x[216], x[215], x[214], x[248], x[247], x[235], x[234], x[251], x[250], x[249], x[233], x[232], x[231], x[246], x[245], x[244], x[6], x[5], x[4], x[27], x[26], x[25], x[222], x[221], x[220], x[262], x[261], x[260], x[219], x[218], x[217], x[205], x[204], x[203], x[9], x[8], x[7], x[30], x[29], x[28], x[225], x[224], x[223], x[15], x[14], x[13], x[228], x[227], x[226], x[213], x[212], x[211], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[148], x[147], x[24], x[23], x[22], x[129], x[128], x[127], x[381], x[3]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[291], x[290], x[329], x[328], x[358], x[357], x[347], x[346], x[333], x[332], x[351], x[350], x[289], x[288], x[287], x[313], x[312], x[356], x[355], x[303], x[302], x[301], x[366], x[365], x[27], x[26], x[25], x[336], x[335], x[334], x[360], x[359], x[316], x[315], x[314], x[309], x[308], x[307], x[331], x[330], x[349], x[348], x[364], x[363], x[324], x[323], x[30], x[29], x[28], x[322], x[321], x[320], x[297], x[296], x[295], x[327], x[326], x[325], x[354], x[353], x[352], x[362], x[361], x[6], x[5], x[4], x[33], x[32], x[31], x[311], x[310], x[339], x[338], x[337], x[306], x[305], x[304], x[319], x[318], x[317], x[345], x[344], x[343], x[300], x[299], x[298], x[15], x[14], x[13], x[24], x[23], x[22], x[9], x[8], x[7], x[342], x[341], x[340], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[294], x[293], x[292], x[237], x[236], x[216], x[215], x[214], x[382], x[3]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[291], x[290], x[329], x[328], x[358], x[357], x[347], x[346], x[333], x[332], x[351], x[350], x[289], x[288], x[287], x[313], x[312], x[356], x[355], x[303], x[302], x[301], x[366], x[365], x[27], x[26], x[25], x[336], x[335], x[334], x[360], x[359], x[316], x[315], x[314], x[309], x[308], x[307], x[331], x[330], x[349], x[348], x[364], x[363], x[324], x[323], x[30], x[29], x[28], x[322], x[321], x[320], x[297], x[296], x[295], x[327], x[326], x[325], x[354], x[353], x[352], x[362], x[361], x[6], x[5], x[4], x[33], x[32], x[31], x[311], x[310], x[339], x[338], x[337], x[306], x[305], x[304], x[319], x[318], x[317], x[345], x[344], x[343], x[300], x[299], x[298], x[15], x[14], x[13], x[24], x[23], x[22], x[9], x[8], x[7], x[342], x[341], x[340], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[294], x[293], x[292], x[237], x[236], x[216], x[215], x[214], x[382], x[3]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[329], x[328], x[347], x[346], x[364], x[363], x[333], x[332], x[324], x[323], x[291], x[290], x[313], x[312], x[356], x[355], x[366], x[365], x[349], x[348], x[303], x[302], x[301], x[316], x[315], x[314], x[345], x[344], x[343], x[362], x[361], x[309], x[308], x[307], x[27], x[26], x[25], x[300], x[299], x[298], x[289], x[288], x[287], x[297], x[296], x[295], x[327], x[326], x[325], x[354], x[353], x[352], x[319], x[318], x[317], x[331], x[330], x[360], x[359], x[30], x[29], x[28], x[342], x[341], x[340], x[351], x[350], x[358], x[357], x[6], x[5], x[4], x[33], x[32], x[31], x[306], x[305], x[304], x[339], x[338], x[337], x[311], x[310], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[322], x[321], x[320], x[336], x[335], x[334], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[294], x[293], x[292], x[248], x[247], x[228], x[227], x[226], x[383], x[3]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[329], x[328], x[347], x[346], x[364], x[363], x[333], x[332], x[324], x[323], x[291], x[290], x[313], x[312], x[356], x[355], x[366], x[365], x[349], x[348], x[303], x[302], x[301], x[316], x[315], x[314], x[345], x[344], x[343], x[362], x[361], x[309], x[308], x[307], x[27], x[26], x[25], x[300], x[299], x[298], x[289], x[288], x[287], x[297], x[296], x[295], x[327], x[326], x[325], x[354], x[353], x[352], x[319], x[318], x[317], x[331], x[330], x[360], x[359], x[30], x[29], x[28], x[342], x[341], x[340], x[351], x[350], x[358], x[357], x[6], x[5], x[4], x[33], x[32], x[31], x[306], x[305], x[304], x[339], x[338], x[337], x[311], x[310], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[322], x[321], x[320], x[336], x[335], x[334], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[294], x[293], x[292], x[248], x[247], x[228], x[227], x[226], x[383], x[3]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[356], x[355], x[347], x[346], x[327], x[326], x[325], x[364], x[363], x[316], x[315], x[314], x[313], x[312], x[291], x[290], x[366], x[365], x[349], x[348], x[324], x[323], x[362], x[361], x[311], x[310], x[27], x[26], x[25], x[351], x[350], x[333], x[332], x[331], x[330], x[329], x[328], x[345], x[344], x[343], x[297], x[296], x[295], x[289], x[288], x[287], x[30], x[29], x[28], x[360], x[359], x[358], x[357], x[354], x[353], x[352], x[319], x[318], x[317], x[300], x[299], x[298], x[342], x[341], x[340], x[294], x[293], x[292], x[6], x[5], x[4], x[33], x[32], x[31], x[322], x[321], x[320], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[339], x[338], x[337], x[336], x[335], x[334], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[239], x[238], x[219], x[218], x[217], x[384], x[3]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[356], x[355], x[347], x[346], x[327], x[326], x[325], x[364], x[363], x[316], x[315], x[314], x[313], x[312], x[291], x[290], x[366], x[365], x[349], x[348], x[324], x[323], x[362], x[361], x[311], x[310], x[27], x[26], x[25], x[351], x[350], x[333], x[332], x[331], x[330], x[329], x[328], x[345], x[344], x[343], x[297], x[296], x[295], x[289], x[288], x[287], x[30], x[29], x[28], x[360], x[359], x[358], x[357], x[354], x[353], x[352], x[319], x[318], x[317], x[300], x[299], x[298], x[342], x[341], x[340], x[294], x[293], x[292], x[6], x[5], x[4], x[33], x[32], x[31], x[322], x[321], x[320], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[339], x[338], x[337], x[336], x[335], x[334], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[239], x[238], x[219], x[218], x[217], x[384], x[3]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[366], x[365], x[364], x[363], x[331], x[330], x[362], x[361], x[313], x[312], x[351], x[350], x[333], x[332], x[354], x[353], x[352], x[358], x[357], x[347], x[346], x[356], x[355], x[27], x[26], x[25], x[345], x[344], x[343], x[306], x[305], x[304], x[349], x[348], x[329], x[328], x[291], x[290], x[342], x[341], x[340], x[297], x[296], x[295], x[30], x[29], x[28], x[324], x[323], x[322], x[321], x[320], x[311], x[310], x[360], x[359], x[309], x[308], x[307], x[336], x[335], x[334], x[316], x[315], x[314], x[327], x[326], x[325], x[6], x[5], x[4], x[33], x[32], x[31], x[319], x[318], x[317], x[303], x[302], x[301], x[289], x[288], x[287], x[15], x[14], x[13], x[24], x[23], x[22], x[300], x[299], x[298], x[294], x[293], x[292], x[339], x[338], x[337], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[9], x[8], x[7], x[235], x[234], x[213], x[212], x[211], x[385], x[3]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[366], x[365], x[364], x[363], x[331], x[330], x[362], x[361], x[313], x[312], x[351], x[350], x[333], x[332], x[354], x[353], x[352], x[358], x[357], x[347], x[346], x[356], x[355], x[27], x[26], x[25], x[345], x[344], x[343], x[306], x[305], x[304], x[349], x[348], x[329], x[328], x[291], x[290], x[342], x[341], x[340], x[297], x[296], x[295], x[30], x[29], x[28], x[324], x[323], x[322], x[321], x[320], x[311], x[310], x[360], x[359], x[309], x[308], x[307], x[336], x[335], x[334], x[316], x[315], x[314], x[327], x[326], x[325], x[6], x[5], x[4], x[33], x[32], x[31], x[319], x[318], x[317], x[303], x[302], x[301], x[289], x[288], x[287], x[15], x[14], x[13], x[24], x[23], x[22], x[300], x[299], x[298], x[294], x[293], x[292], x[339], x[338], x[337], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[9], x[8], x[7], x[235], x[234], x[213], x[212], x[211], x[385], x[3]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[104], x[103], x[81], x[80], x[39], x[38], x[74], x[73], x[114], x[113], x[79], x[78], x[110], x[109], x[98], x[97], x[77], x[76], x[75], x[102], x[101], x[57], x[56], x[55], x[63], x[62], x[37], x[36], x[35], x[27], x[26], x[25], x[51], x[50], x[49], x[96], x[95], x[94], x[54], x[53], x[52], x[90], x[89], x[88], x[66], x[65], x[64], x[108], x[107], x[30], x[29], x[28], x[72], x[71], x[70], x[61], x[60], x[112], x[111], x[48], x[47], x[46], x[100], x[99], x[59], x[58], x[106], x[105], x[6], x[5], x[4], x[33], x[32], x[31], x[87], x[86], x[85], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[45], x[44], x[43], x[93], x[92], x[91], x[69], x[68], x[67], x[42], x[41], x[40], x[84], x[83], x[82], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[243], x[242], x[225], x[224], x[223], x[386], x[3]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[104], x[103], x[81], x[80], x[39], x[38], x[74], x[73], x[114], x[113], x[79], x[78], x[110], x[109], x[98], x[97], x[77], x[76], x[75], x[102], x[101], x[57], x[56], x[55], x[63], x[62], x[37], x[36], x[35], x[27], x[26], x[25], x[51], x[50], x[49], x[96], x[95], x[94], x[54], x[53], x[52], x[90], x[89], x[88], x[66], x[65], x[64], x[108], x[107], x[30], x[29], x[28], x[72], x[71], x[70], x[61], x[60], x[112], x[111], x[48], x[47], x[46], x[100], x[99], x[59], x[58], x[106], x[105], x[6], x[5], x[4], x[33], x[32], x[31], x[87], x[86], x[85], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[45], x[44], x[43], x[93], x[92], x[91], x[69], x[68], x[67], x[42], x[41], x[40], x[84], x[83], x[82], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[243], x[242], x[225], x[224], x[223], x[386], x[3]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[104], x[103], x[74], x[73], x[114], x[113], x[81], x[80], x[39], x[38], x[77], x[76], x[75], x[79], x[78], x[98], x[97], x[51], x[50], x[49], x[96], x[95], x[94], x[57], x[56], x[55], x[63], x[62], x[37], x[36], x[35], x[102], x[101], x[110], x[109], x[100], x[99], x[27], x[26], x[25], x[59], x[58], x[54], x[53], x[52], x[66], x[65], x[64], x[112], x[111], x[108], x[107], x[106], x[105], x[30], x[29], x[28], x[48], x[47], x[46], x[72], x[71], x[70], x[90], x[89], x[88], x[61], x[60], x[69], x[68], x[67], x[6], x[5], x[4], x[33], x[32], x[31], x[42], x[41], x[40], x[93], x[92], x[91], x[87], x[86], x[85], x[84], x[83], x[82], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[45], x[44], x[43], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[282], x[281], x[268], x[267], x[266], x[387], x[3]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[104], x[103], x[74], x[73], x[114], x[113], x[81], x[80], x[39], x[38], x[77], x[76], x[75], x[79], x[78], x[98], x[97], x[51], x[50], x[49], x[96], x[95], x[94], x[57], x[56], x[55], x[63], x[62], x[37], x[36], x[35], x[102], x[101], x[110], x[109], x[100], x[99], x[27], x[26], x[25], x[59], x[58], x[54], x[53], x[52], x[66], x[65], x[64], x[112], x[111], x[108], x[107], x[106], x[105], x[30], x[29], x[28], x[48], x[47], x[46], x[72], x[71], x[70], x[90], x[89], x[88], x[61], x[60], x[69], x[68], x[67], x[6], x[5], x[4], x[33], x[32], x[31], x[42], x[41], x[40], x[93], x[92], x[91], x[87], x[86], x[85], x[84], x[83], x[82], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[45], x[44], x[43], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[282], x[281], x[268], x[267], x[266], x[387], x[3]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[114], x[113], x[104], x[103], x[81], x[80], x[102], x[101], x[98], x[97], x[106], x[105], x[61], x[60], x[96], x[95], x[94], x[112], x[111], x[110], x[109], x[77], x[76], x[75], x[74], x[73], x[39], x[38], x[57], x[56], x[55], x[63], x[62], x[100], x[99], x[27], x[26], x[25], x[72], x[71], x[70], x[79], x[78], x[66], x[65], x[64], x[84], x[83], x[82], x[30], x[29], x[28], x[45], x[44], x[43], x[93], x[92], x[91], x[90], x[89], x[88], x[51], x[50], x[49], x[37], x[36], x[35], x[48], x[47], x[46], x[69], x[68], x[67], x[59], x[58], x[108], x[107], x[6], x[5], x[4], x[33], x[32], x[31], x[54], x[53], x[52], x[9], x[8], x[7], x[24], x[23], x[22], x[15], x[14], x[13], x[42], x[41], x[40], x[87], x[86], x[85], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[276], x[275], x[257], x[256], x[255], x[388], x[3]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[114], x[113], x[104], x[103], x[81], x[80], x[102], x[101], x[98], x[97], x[106], x[105], x[61], x[60], x[96], x[95], x[94], x[112], x[111], x[110], x[109], x[77], x[76], x[75], x[74], x[73], x[39], x[38], x[57], x[56], x[55], x[63], x[62], x[100], x[99], x[27], x[26], x[25], x[72], x[71], x[70], x[79], x[78], x[66], x[65], x[64], x[84], x[83], x[82], x[30], x[29], x[28], x[45], x[44], x[43], x[93], x[92], x[91], x[90], x[89], x[88], x[51], x[50], x[49], x[37], x[36], x[35], x[48], x[47], x[46], x[69], x[68], x[67], x[59], x[58], x[108], x[107], x[6], x[5], x[4], x[33], x[32], x[31], x[54], x[53], x[52], x[9], x[8], x[7], x[24], x[23], x[22], x[15], x[14], x[13], x[42], x[41], x[40], x[87], x[86], x[85], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[276], x[275], x[257], x[256], x[255], x[388], x[3]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[74], x[73], x[98], x[97], x[104], x[103], x[114], x[113], x[81], x[80], x[79], x[78], x[61], x[60], x[100], x[99], x[39], x[38], x[51], x[50], x[49], x[108], x[107], x[106], x[105], x[66], x[65], x[64], x[63], x[62], x[27], x[26], x[25], x[102], x[101], x[77], x[76], x[75], x[96], x[95], x[94], x[57], x[56], x[55], x[54], x[53], x[52], x[30], x[29], x[28], x[45], x[44], x[43], x[112], x[111], x[110], x[109], x[69], x[68], x[67], x[37], x[36], x[35], x[87], x[86], x[85], x[84], x[83], x[82], x[48], x[47], x[46], x[6], x[5], x[4], x[33], x[32], x[31], x[72], x[71], x[70], x[59], x[58], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[93], x[92], x[91], x[90], x[89], x[88], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[42], x[41], x[40], x[280], x[279], x[265], x[264], x[263], x[389], x[3]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[74], x[73], x[98], x[97], x[104], x[103], x[114], x[113], x[81], x[80], x[79], x[78], x[61], x[60], x[100], x[99], x[39], x[38], x[51], x[50], x[49], x[108], x[107], x[106], x[105], x[66], x[65], x[64], x[63], x[62], x[27], x[26], x[25], x[102], x[101], x[77], x[76], x[75], x[96], x[95], x[94], x[57], x[56], x[55], x[54], x[53], x[52], x[30], x[29], x[28], x[45], x[44], x[43], x[112], x[111], x[110], x[109], x[69], x[68], x[67], x[37], x[36], x[35], x[87], x[86], x[85], x[84], x[83], x[82], x[48], x[47], x[46], x[6], x[5], x[4], x[33], x[32], x[31], x[72], x[71], x[70], x[59], x[58], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[93], x[92], x[91], x[90], x[89], x[88], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[42], x[41], x[40], x[280], x[279], x[265], x[264], x[263], x[389], x[3]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[188], x[187], x[123], x[122], x[159], x[158], x[192], x[191], x[152], x[151], x[165], x[164], x[163], x[186], x[185], x[150], x[149], x[184], x[183], x[167], x[166], x[148], x[147], x[121], x[120], x[119], x[198], x[197], x[27], x[26], x[25], x[141], x[140], x[139], x[173], x[172], x[171], x[135], x[134], x[133], x[190], x[189], x[154], x[153], x[196], x[195], x[30], x[29], x[28], x[162], x[161], x[160], x[132], x[131], x[130], x[157], x[156], x[155], x[146], x[145], x[194], x[193], x[144], x[143], x[142], x[129], x[128], x[127], x[182], x[181], x[180], x[6], x[5], x[4], x[33], x[32], x[31], x[170], x[169], x[168], x[138], x[137], x[136], x[179], x[178], x[177], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[126], x[125], x[124], x[176], x[175], x[174], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[324], x[323], x[300], x[299], x[298], x[390], x[3]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[188], x[187], x[123], x[122], x[159], x[158], x[192], x[191], x[152], x[151], x[165], x[164], x[163], x[186], x[185], x[150], x[149], x[184], x[183], x[167], x[166], x[148], x[147], x[121], x[120], x[119], x[198], x[197], x[27], x[26], x[25], x[141], x[140], x[139], x[173], x[172], x[171], x[135], x[134], x[133], x[190], x[189], x[154], x[153], x[196], x[195], x[30], x[29], x[28], x[162], x[161], x[160], x[132], x[131], x[130], x[157], x[156], x[155], x[146], x[145], x[194], x[193], x[144], x[143], x[142], x[129], x[128], x[127], x[182], x[181], x[180], x[6], x[5], x[4], x[33], x[32], x[31], x[170], x[169], x[168], x[138], x[137], x[136], x[179], x[178], x[177], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[126], x[125], x[124], x[176], x[175], x[174], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[324], x[323], x[300], x[299], x[298], x[390], x[3]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[188], x[187], x[159], x[158], x[123], x[122], x[186], x[185], x[152], x[151], x[165], x[164], x[163], x[190], x[189], x[141], x[140], x[139], x[148], x[147], x[121], x[120], x[119], x[154], x[153], x[150], x[149], x[167], x[166], x[184], x[183], x[192], x[191], x[198], x[197], x[196], x[195], x[162], x[161], x[160], x[135], x[134], x[133], x[194], x[193], x[170], x[169], x[168], x[129], x[128], x[127], x[138], x[137], x[136], x[132], x[131], x[130], x[144], x[143], x[142], x[157], x[156], x[155], x[173], x[172], x[171], x[146], x[145], x[182], x[181], x[180], x[179], x[178], x[177], x[6], x[5], x[4], x[27], x[26], x[25], x[176], x[175], x[174], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[126], x[125], x[124], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[366], x[365], x[24], x[23], x[22], x[354], x[353], x[352], x[391], x[3]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[188], x[187], x[159], x[158], x[123], x[122], x[186], x[185], x[152], x[151], x[165], x[164], x[163], x[190], x[189], x[141], x[140], x[139], x[148], x[147], x[121], x[120], x[119], x[154], x[153], x[150], x[149], x[167], x[166], x[184], x[183], x[192], x[191], x[198], x[197], x[196], x[195], x[162], x[161], x[160], x[135], x[134], x[133], x[194], x[193], x[170], x[169], x[168], x[129], x[128], x[127], x[138], x[137], x[136], x[132], x[131], x[130], x[144], x[143], x[142], x[157], x[156], x[155], x[173], x[172], x[171], x[146], x[145], x[182], x[181], x[180], x[179], x[178], x[177], x[6], x[5], x[4], x[27], x[26], x[25], x[176], x[175], x[174], x[9], x[8], x[7], x[15], x[14], x[13], x[30], x[29], x[28], x[126], x[125], x[124], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[33], x[32], x[31], x[366], x[365], x[24], x[23], x[22], x[354], x[353], x[352], x[391], x[3]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[188], x[187], x[196], x[195], x[186], x[185], x[184], x[183], x[152], x[151], x[190], x[189], x[146], x[145], x[194], x[193], x[192], x[191], x[165], x[164], x[163], x[159], x[158], x[123], x[122], x[167], x[166], x[148], x[147], x[179], x[178], x[177], x[27], x[26], x[25], x[162], x[161], x[160], x[157], x[156], x[155], x[135], x[134], x[133], x[170], x[169], x[168], x[154], x[153], x[198], x[197], x[30], x[29], x[28], x[126], x[125], x[124], x[176], x[175], x[174], x[173], x[172], x[171], x[150], x[149], x[141], x[140], x[139], x[121], x[120], x[119], x[144], x[143], x[142], x[129], x[128], x[127], x[6], x[5], x[4], x[33], x[32], x[31], x[138], x[137], x[136], x[182], x[181], x[180], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[132], x[131], x[130], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[364], x[363], x[345], x[344], x[343], x[392], x[3]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[188], x[187], x[196], x[195], x[186], x[185], x[184], x[183], x[152], x[151], x[190], x[189], x[146], x[145], x[194], x[193], x[192], x[191], x[165], x[164], x[163], x[159], x[158], x[123], x[122], x[167], x[166], x[148], x[147], x[179], x[178], x[177], x[27], x[26], x[25], x[162], x[161], x[160], x[157], x[156], x[155], x[135], x[134], x[133], x[170], x[169], x[168], x[154], x[153], x[198], x[197], x[30], x[29], x[28], x[126], x[125], x[124], x[176], x[175], x[174], x[173], x[172], x[171], x[150], x[149], x[141], x[140], x[139], x[121], x[120], x[119], x[144], x[143], x[142], x[129], x[128], x[127], x[6], x[5], x[4], x[33], x[32], x[31], x[138], x[137], x[136], x[182], x[181], x[180], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[132], x[131], x[130], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[364], x[363], x[345], x[344], x[343], x[392], x[3]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[159], x[158], x[190], x[189], x[188], x[187], x[198], x[197], x[196], x[195], x[167], x[166], x[146], x[145], x[123], x[122], x[141], x[140], x[139], x[186], x[185], x[152], x[151], x[150], x[149], x[148], x[147], x[27], x[26], x[25], x[184], x[183], x[170], x[169], x[168], x[165], x[164], x[163], x[182], x[181], x[180], x[179], x[178], x[177], x[144], x[143], x[142], x[30], x[29], x[28], x[126], x[125], x[124], x[194], x[193], x[192], x[191], x[154], x[153], x[121], x[120], x[119], x[162], x[161], x[160], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[6], x[5], x[4], x[33], x[32], x[31], x[157], x[156], x[155], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[176], x[175], x[174], x[173], x[172], x[171], x[138], x[137], x[136], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[362], x[361], x[342], x[341], x[340], x[393], x[3]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[159], x[158], x[190], x[189], x[188], x[187], x[198], x[197], x[196], x[195], x[167], x[166], x[146], x[145], x[123], x[122], x[141], x[140], x[139], x[186], x[185], x[152], x[151], x[150], x[149], x[148], x[147], x[27], x[26], x[25], x[184], x[183], x[170], x[169], x[168], x[165], x[164], x[163], x[182], x[181], x[180], x[179], x[178], x[177], x[144], x[143], x[142], x[30], x[29], x[28], x[126], x[125], x[124], x[194], x[193], x[192], x[191], x[154], x[153], x[121], x[120], x[119], x[162], x[161], x[160], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[6], x[5], x[4], x[33], x[32], x[31], x[157], x[156], x[155], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[176], x[175], x[174], x[173], x[172], x[171], x[138], x[137], x[136], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[362], x[361], x[342], x[341], x[340], x[393], x[3]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[280], x[279], x[259], x[258], x[276], x[275], x[239], x[238], x[207], x[206], x[230], x[229], x[270], x[269], x[237], x[236], x[265], x[264], x[263], x[248], x[247], x[235], x[234], x[278], x[277], x[27], x[26], x[25], x[233], x[232], x[231], x[257], x[256], x[255], x[243], x[242], x[282], x[281], x[219], x[218], x[217], x[205], x[204], x[203], x[274], x[273], x[241], x[240], x[30], x[29], x[28], x[210], x[209], x[208], x[246], x[245], x[244], x[216], x[215], x[214], x[228], x[227], x[226], x[213], x[212], x[211], x[262], x[261], x[260], x[272], x[271], x[33], x[32], x[31], x[225], x[224], x[223], x[268], x[267], x[266], x[254], x[253], x[252], x[222], x[221], x[220], x[9], x[8], x[7], x[24], x[23], x[22], x[6], x[5], x[4], x[15], x[14], x[13], x[251], x[250], x[249], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[61], x[60], x[45], x[44], x[43], x[394], x[3]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[280], x[279], x[259], x[258], x[276], x[275], x[239], x[238], x[207], x[206], x[230], x[229], x[270], x[269], x[237], x[236], x[265], x[264], x[263], x[248], x[247], x[235], x[234], x[278], x[277], x[27], x[26], x[25], x[233], x[232], x[231], x[257], x[256], x[255], x[243], x[242], x[282], x[281], x[219], x[218], x[217], x[205], x[204], x[203], x[274], x[273], x[241], x[240], x[30], x[29], x[28], x[210], x[209], x[208], x[246], x[245], x[244], x[216], x[215], x[214], x[228], x[227], x[226], x[213], x[212], x[211], x[262], x[261], x[260], x[272], x[271], x[33], x[32], x[31], x[225], x[224], x[223], x[268], x[267], x[266], x[254], x[253], x[252], x[222], x[221], x[220], x[9], x[8], x[7], x[24], x[23], x[22], x[6], x[5], x[4], x[15], x[14], x[13], x[251], x[250], x[249], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[61], x[60], x[45], x[44], x[43], x[394], x[3]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[259], x[258], x[230], x[229], x[270], x[269], x[239], x[238], x[207], x[206], x[276], x[275], x[280], x[279], x[274], x[273], x[235], x[234], x[233], x[232], x[231], x[241], x[240], x[237], x[236], x[248], x[247], x[282], x[281], x[278], x[277], x[210], x[209], x[208], x[246], x[245], x[244], x[27], x[26], x[25], x[219], x[218], x[217], x[205], x[204], x[203], x[257], x[256], x[255], x[265], x[264], x[263], x[243], x[242], x[254], x[253], x[252], x[272], x[271], x[30], x[29], x[28], x[213], x[212], x[211], x[222], x[221], x[220], x[216], x[215], x[214], x[228], x[227], x[226], x[268], x[267], x[266], x[262], x[261], x[260], x[6], x[5], x[4], x[33], x[32], x[31], x[225], x[224], x[223], x[251], x[250], x[249], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[112], x[111], x[93], x[92], x[91], x[395], x[3]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[259], x[258], x[230], x[229], x[270], x[269], x[239], x[238], x[207], x[206], x[276], x[275], x[280], x[279], x[274], x[273], x[235], x[234], x[233], x[232], x[231], x[241], x[240], x[237], x[236], x[248], x[247], x[282], x[281], x[278], x[277], x[210], x[209], x[208], x[246], x[245], x[244], x[27], x[26], x[25], x[219], x[218], x[217], x[205], x[204], x[203], x[257], x[256], x[255], x[265], x[264], x[263], x[243], x[242], x[254], x[253], x[252], x[272], x[271], x[30], x[29], x[28], x[213], x[212], x[211], x[222], x[221], x[220], x[216], x[215], x[214], x[228], x[227], x[226], x[268], x[267], x[266], x[262], x[261], x[260], x[6], x[5], x[4], x[33], x[32], x[31], x[225], x[224], x[223], x[251], x[250], x[249], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[112], x[111], x[93], x[92], x[91], x[395], x[3]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[276], x[275], x[243], x[242], x[270], x[269], x[282], x[281], x[280], x[279], x[259], x[258], x[239], x[238], x[274], x[273], x[272], x[271], x[257], x[256], x[255], x[248], x[247], x[235], x[234], x[27], x[26], x[25], x[225], x[224], x[223], x[246], x[245], x[244], x[268], x[267], x[266], x[265], x[264], x[263], x[233], x[232], x[231], x[230], x[229], x[207], x[206], x[219], x[218], x[217], x[254], x[253], x[252], x[251], x[250], x[249], x[241], x[240], x[278], x[277], x[30], x[29], x[28], x[237], x[236], x[228], x[227], x[226], x[213], x[212], x[211], x[6], x[5], x[4], x[33], x[32], x[31], x[210], x[209], x[208], x[205], x[204], x[203], x[222], x[221], x[220], x[262], x[261], x[260], x[9], x[8], x[7], x[24], x[23], x[22], x[216], x[215], x[214], x[15], x[14], x[13], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[102], x[101], x[72], x[71], x[70], x[396], x[3]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[276], x[275], x[243], x[242], x[270], x[269], x[282], x[281], x[280], x[279], x[259], x[258], x[239], x[238], x[274], x[273], x[272], x[271], x[257], x[256], x[255], x[248], x[247], x[235], x[234], x[27], x[26], x[25], x[225], x[224], x[223], x[246], x[245], x[244], x[268], x[267], x[266], x[265], x[264], x[263], x[233], x[232], x[231], x[230], x[229], x[207], x[206], x[219], x[218], x[217], x[254], x[253], x[252], x[251], x[250], x[249], x[241], x[240], x[278], x[277], x[30], x[29], x[28], x[237], x[236], x[228], x[227], x[226], x[213], x[212], x[211], x[6], x[5], x[4], x[33], x[32], x[31], x[210], x[209], x[208], x[205], x[204], x[203], x[222], x[221], x[220], x[262], x[261], x[260], x[9], x[8], x[7], x[24], x[23], x[22], x[216], x[215], x[214], x[15], x[14], x[13], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[102], x[101], x[72], x[71], x[70], x[396], x[3]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[243], x[242], x[274], x[273], x[230], x[229], x[278], x[277], x[248], x[247], x[276], x[275], x[259], x[258], x[270], x[269], x[272], x[271], x[239], x[238], x[237], x[236], x[235], x[234], x[27], x[26], x[25], x[225], x[224], x[223], x[282], x[281], x[280], x[279], x[254], x[253], x[252], x[207], x[206], x[210], x[209], x[208], x[262], x[261], x[260], x[228], x[227], x[226], x[30], x[29], x[28], x[257], x[256], x[255], x[241], x[240], x[233], x[232], x[231], x[246], x[245], x[244], x[251], x[250], x[249], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[33], x[32], x[31], x[268], x[267], x[266], x[265], x[264], x[263], x[205], x[204], x[203], x[24], x[23], x[22], x[222], x[221], x[220], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[110], x[109], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[90], x[89], x[88], x[397], x[3]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[243], x[242], x[274], x[273], x[230], x[229], x[278], x[277], x[248], x[247], x[276], x[275], x[259], x[258], x[270], x[269], x[272], x[271], x[239], x[238], x[237], x[236], x[235], x[234], x[27], x[26], x[25], x[225], x[224], x[223], x[282], x[281], x[280], x[279], x[254], x[253], x[252], x[207], x[206], x[210], x[209], x[208], x[262], x[261], x[260], x[228], x[227], x[226], x[30], x[29], x[28], x[257], x[256], x[255], x[241], x[240], x[233], x[232], x[231], x[246], x[245], x[244], x[251], x[250], x[249], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[33], x[32], x[31], x[268], x[267], x[266], x[265], x[264], x[263], x[205], x[204], x[203], x[24], x[23], x[22], x[222], x[221], x[220], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[110], x[109], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[90], x[89], x[88], x[397], x[3]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[333], x[332], x[347], x[346], x[331], x[330], x[364], x[363], x[362], x[361], x[349], x[348], x[329], x[328], x[291], x[290], x[313], x[312], x[356], x[355], x[309], x[308], x[307], x[27], x[26], x[25], x[316], x[315], x[314], x[306], x[305], x[304], x[345], x[344], x[343], x[342], x[341], x[340], x[324], x[323], x[366], x[365], x[319], x[318], x[317], x[303], x[302], x[301], x[289], x[288], x[287], x[360], x[359], x[30], x[29], x[28], x[297], x[296], x[295], x[327], x[326], x[325], x[351], x[350], x[311], x[310], x[358], x[357], x[6], x[5], x[4], x[33], x[32], x[31], x[300], x[299], x[298], x[354], x[353], x[352], x[339], x[338], x[337], x[15], x[14], x[13], x[24], x[23], x[22], x[9], x[8], x[7], x[322], x[321], x[320], x[294], x[293], x[292], x[336], x[335], x[334], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[146], x[145], x[126], x[125], x[124], x[398], x[3]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[333], x[332], x[347], x[346], x[331], x[330], x[364], x[363], x[362], x[361], x[349], x[348], x[329], x[328], x[291], x[290], x[313], x[312], x[356], x[355], x[309], x[308], x[307], x[27], x[26], x[25], x[316], x[315], x[314], x[306], x[305], x[304], x[345], x[344], x[343], x[342], x[341], x[340], x[324], x[323], x[366], x[365], x[319], x[318], x[317], x[303], x[302], x[301], x[289], x[288], x[287], x[360], x[359], x[30], x[29], x[28], x[297], x[296], x[295], x[327], x[326], x[325], x[351], x[350], x[311], x[310], x[358], x[357], x[6], x[5], x[4], x[33], x[32], x[31], x[300], x[299], x[298], x[354], x[353], x[352], x[339], x[338], x[337], x[15], x[14], x[13], x[24], x[23], x[22], x[9], x[8], x[7], x[322], x[321], x[320], x[294], x[293], x[292], x[336], x[335], x[334], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[146], x[145], x[126], x[125], x[124], x[398], x[3]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[333], x[332], x[347], x[346], x[313], x[312], x[356], x[355], x[329], x[328], x[291], x[290], x[331], x[330], x[349], x[348], x[364], x[363], x[309], x[308], x[307], x[316], x[315], x[314], x[362], x[361], x[366], x[365], x[351], x[350], x[297], x[296], x[295], x[327], x[326], x[325], x[27], x[26], x[25], x[303], x[302], x[301], x[289], x[288], x[287], x[311], x[310], x[306], x[305], x[304], x[319], x[318], x[317], x[345], x[344], x[343], x[324], x[323], x[360], x[359], x[358], x[357], x[30], x[29], x[28], x[342], x[341], x[340], x[354], x[353], x[352], x[322], x[321], x[320], x[6], x[5], x[4], x[33], x[32], x[31], x[294], x[293], x[292], x[300], x[299], x[298], x[339], x[338], x[337], x[336], x[335], x[334], x[15], x[14], x[13], x[24], x[23], x[22], x[9], x[8], x[7], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[194], x[193], x[176], x[175], x[174], x[399], x[3]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[333], x[332], x[347], x[346], x[313], x[312], x[356], x[355], x[329], x[328], x[291], x[290], x[331], x[330], x[349], x[348], x[364], x[363], x[309], x[308], x[307], x[316], x[315], x[314], x[362], x[361], x[366], x[365], x[351], x[350], x[297], x[296], x[295], x[327], x[326], x[325], x[27], x[26], x[25], x[303], x[302], x[301], x[289], x[288], x[287], x[311], x[310], x[306], x[305], x[304], x[319], x[318], x[317], x[345], x[344], x[343], x[324], x[323], x[360], x[359], x[358], x[357], x[30], x[29], x[28], x[342], x[341], x[340], x[354], x[353], x[352], x[322], x[321], x[320], x[6], x[5], x[4], x[33], x[32], x[31], x[294], x[293], x[292], x[300], x[299], x[298], x[339], x[338], x[337], x[336], x[335], x[334], x[15], x[14], x[13], x[24], x[23], x[22], x[9], x[8], x[7], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[194], x[193], x[176], x[175], x[174], x[399], x[3]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[364], x[363], x[333], x[332], x[324], x[323], x[356], x[355], x[366], x[365], x[347], x[346], x[349], x[348], x[329], x[328], x[358], x[357], x[345], x[344], x[343], x[362], x[361], x[309], x[308], x[307], x[351], x[350], x[27], x[26], x[25], x[300], x[299], x[298], x[327], x[326], x[325], x[354], x[353], x[352], x[331], x[330], x[316], x[315], x[314], x[313], x[312], x[291], x[290], x[319], x[318], x[317], x[303], x[302], x[301], x[336], x[335], x[334], x[30], x[29], x[28], x[342], x[341], x[340], x[322], x[321], x[320], x[311], x[310], x[360], x[359], x[6], x[5], x[4], x[33], x[32], x[31], x[306], x[305], x[304], x[297], x[296], x[295], x[289], x[288], x[287], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[294], x[293], x[292], x[339], x[338], x[337], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[184], x[183], x[157], x[156], x[155], x[400], x[3]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[364], x[363], x[333], x[332], x[324], x[323], x[356], x[355], x[366], x[365], x[347], x[346], x[349], x[348], x[329], x[328], x[358], x[357], x[345], x[344], x[343], x[362], x[361], x[309], x[308], x[307], x[351], x[350], x[27], x[26], x[25], x[300], x[299], x[298], x[327], x[326], x[325], x[354], x[353], x[352], x[331], x[330], x[316], x[315], x[314], x[313], x[312], x[291], x[290], x[319], x[318], x[317], x[303], x[302], x[301], x[336], x[335], x[334], x[30], x[29], x[28], x[342], x[341], x[340], x[322], x[321], x[320], x[311], x[310], x[360], x[359], x[6], x[5], x[4], x[33], x[32], x[31], x[306], x[305], x[304], x[297], x[296], x[295], x[289], x[288], x[287], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[294], x[293], x[292], x[339], x[338], x[337], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[184], x[183], x[157], x[156], x[155], x[400], x[3]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[349], x[348], x[324], x[323], x[313], x[312], x[333], x[332], x[331], x[330], x[329], x[328], x[364], x[363], x[351], x[350], x[347], x[346], x[356], x[355], x[360], x[359], x[358], x[357], x[319], x[318], x[317], x[27], x[26], x[25], x[300], x[299], x[298], x[366], x[365], x[291], x[290], x[297], x[296], x[295], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[30], x[29], x[28], x[345], x[344], x[343], x[362], x[361], x[322], x[321], x[320], x[316], x[315], x[314], x[327], x[326], x[325], x[339], x[338], x[337], x[336], x[335], x[334], x[33], x[32], x[31], x[354], x[353], x[352], x[311], x[310], x[289], x[288], x[287], x[24], x[23], x[22], x[342], x[341], x[340], x[6], x[5], x[4], x[294], x[293], x[292], x[9], x[8], x[7], x[15], x[14], x[13], x[192], x[191], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[173], x[172], x[171], x[401], x[3]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[349], x[348], x[324], x[323], x[313], x[312], x[333], x[332], x[331], x[330], x[329], x[328], x[364], x[363], x[351], x[350], x[347], x[346], x[356], x[355], x[360], x[359], x[358], x[357], x[319], x[318], x[317], x[27], x[26], x[25], x[300], x[299], x[298], x[366], x[365], x[291], x[290], x[297], x[296], x[295], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[30], x[29], x[28], x[345], x[344], x[343], x[362], x[361], x[322], x[321], x[320], x[316], x[315], x[314], x[327], x[326], x[325], x[339], x[338], x[337], x[336], x[335], x[334], x[33], x[32], x[31], x[354], x[353], x[352], x[311], x[310], x[289], x[288], x[287], x[24], x[23], x[22], x[342], x[341], x[340], x[6], x[5], x[4], x[294], x[293], x[292], x[9], x[8], x[7], x[15], x[14], x[13], x[192], x[191], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[173], x[172], x[171], x[401], x[3]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[114], x[113], x[104], x[103], x[106], x[105], x[102], x[101], x[112], x[111], x[110], x[109], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[39], x[38], x[74], x[73], x[84], x[83], x[82], x[27], x[26], x[25], x[72], x[71], x[70], x[63], x[62], x[93], x[92], x[91], x[90], x[89], x[88], x[69], x[68], x[67], x[108], x[107], x[66], x[65], x[64], x[30], x[29], x[28], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[37], x[36], x[35], x[51], x[50], x[49], x[33], x[32], x[31], x[48], x[47], x[46], x[87], x[86], x[85], x[24], x[23], x[22], x[45], x[44], x[43], x[42], x[41], x[40], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[154], x[153], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[138], x[137], x[136], x[402], x[3]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[114], x[113], x[104], x[103], x[106], x[105], x[102], x[101], x[112], x[111], x[110], x[109], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[39], x[38], x[74], x[73], x[84], x[83], x[82], x[27], x[26], x[25], x[72], x[71], x[70], x[63], x[62], x[93], x[92], x[91], x[90], x[89], x[88], x[69], x[68], x[67], x[108], x[107], x[66], x[65], x[64], x[30], x[29], x[28], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[37], x[36], x[35], x[51], x[50], x[49], x[33], x[32], x[31], x[48], x[47], x[46], x[87], x[86], x[85], x[24], x[23], x[22], x[45], x[44], x[43], x[42], x[41], x[40], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[154], x[153], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[138], x[137], x[136], x[402], x[3]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[104], x[103], x[114], x[113], x[74], x[73], x[81], x[80], x[39], x[38], x[77], x[76], x[75], x[96], x[95], x[94], x[79], x[78], x[98], x[97], x[51], x[50], x[49], x[112], x[111], x[100], x[99], x[106], x[105], x[57], x[56], x[55], x[63], x[62], x[37], x[36], x[35], x[102], x[101], x[110], x[109], x[108], x[107], x[27], x[26], x[25], x[61], x[60], x[54], x[53], x[52], x[66], x[65], x[64], x[93], x[92], x[91], x[69], x[68], x[67], x[84], x[83], x[82], x[30], x[29], x[28], x[48], x[47], x[46], x[72], x[71], x[70], x[90], x[89], x[88], x[59], x[58], x[87], x[86], x[85], x[33], x[32], x[31], x[45], x[44], x[43], x[24], x[23], x[22], x[42], x[41], x[40], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[198], x[197], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[182], x[181], x[180], x[403], x[3]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[104], x[103], x[114], x[113], x[74], x[73], x[81], x[80], x[39], x[38], x[77], x[76], x[75], x[96], x[95], x[94], x[79], x[78], x[98], x[97], x[51], x[50], x[49], x[112], x[111], x[100], x[99], x[106], x[105], x[57], x[56], x[55], x[63], x[62], x[37], x[36], x[35], x[102], x[101], x[110], x[109], x[108], x[107], x[27], x[26], x[25], x[61], x[60], x[54], x[53], x[52], x[66], x[65], x[64], x[93], x[92], x[91], x[69], x[68], x[67], x[84], x[83], x[82], x[30], x[29], x[28], x[48], x[47], x[46], x[72], x[71], x[70], x[90], x[89], x[88], x[59], x[58], x[87], x[86], x[85], x[33], x[32], x[31], x[45], x[44], x[43], x[24], x[23], x[22], x[42], x[41], x[40], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[198], x[197], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[182], x[181], x[180], x[403], x[3]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[81], x[80], x[98], x[97], x[74], x[73], x[63], x[62], x[102], x[101], x[57], x[56], x[55], x[110], x[109], x[100], x[99], x[104], x[103], x[114], x[113], x[59], x[58], x[112], x[111], x[79], x[78], x[39], x[38], x[66], x[65], x[64], x[108], x[107], x[106], x[105], x[51], x[50], x[49], x[48], x[47], x[46], x[72], x[71], x[70], x[61], x[60], x[90], x[89], x[88], x[69], x[68], x[67], x[77], x[76], x[75], x[96], x[95], x[94], x[42], x[41], x[40], x[93], x[92], x[91], x[54], x[53], x[52], x[37], x[36], x[35], x[87], x[86], x[85], x[84], x[83], x[82], x[27], x[26], x[25], x[45], x[44], x[43], x[30], x[29], x[28], x[6], x[5], x[4], x[33], x[32], x[31], x[9], x[8], x[7], x[15], x[14], x[13], x[190], x[189], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[170], x[169], x[168], x[404], x[3]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[81], x[80], x[98], x[97], x[74], x[73], x[63], x[62], x[102], x[101], x[57], x[56], x[55], x[110], x[109], x[100], x[99], x[104], x[103], x[114], x[113], x[59], x[58], x[112], x[111], x[79], x[78], x[39], x[38], x[66], x[65], x[64], x[108], x[107], x[106], x[105], x[51], x[50], x[49], x[48], x[47], x[46], x[72], x[71], x[70], x[61], x[60], x[90], x[89], x[88], x[69], x[68], x[67], x[77], x[76], x[75], x[96], x[95], x[94], x[42], x[41], x[40], x[93], x[92], x[91], x[54], x[53], x[52], x[37], x[36], x[35], x[87], x[86], x[85], x[84], x[83], x[82], x[27], x[26], x[25], x[45], x[44], x[43], x[30], x[29], x[28], x[6], x[5], x[4], x[33], x[32], x[31], x[9], x[8], x[7], x[15], x[14], x[13], x[190], x[189], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[170], x[169], x[168], x[404], x[3]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[104], x[103], x[98], x[97], x[102], x[101], x[110], x[109], x[39], x[38], x[74], x[73], x[114], x[113], x[112], x[111], x[81], x[80], x[61], x[60], x[79], x[78], x[77], x[76], x[75], x[66], x[65], x[64], x[63], x[62], x[72], x[71], x[70], x[90], x[89], x[88], x[37], x[36], x[35], x[27], x[26], x[25], x[100], x[99], x[59], x[58], x[51], x[50], x[49], x[96], x[95], x[94], x[93], x[92], x[91], x[57], x[56], x[55], x[45], x[44], x[43], x[54], x[53], x[52], x[30], x[29], x[28], x[108], x[107], x[106], x[105], x[48], x[47], x[46], x[33], x[32], x[31], x[69], x[68], x[67], x[42], x[41], x[40], x[24], x[23], x[22], x[87], x[86], x[85], x[84], x[83], x[82], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[196], x[195], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[179], x[178], x[177], x[405], x[3]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[104], x[103], x[98], x[97], x[102], x[101], x[110], x[109], x[39], x[38], x[74], x[73], x[114], x[113], x[112], x[111], x[81], x[80], x[61], x[60], x[79], x[78], x[77], x[76], x[75], x[66], x[65], x[64], x[63], x[62], x[72], x[71], x[70], x[90], x[89], x[88], x[37], x[36], x[35], x[27], x[26], x[25], x[100], x[99], x[59], x[58], x[51], x[50], x[49], x[96], x[95], x[94], x[93], x[92], x[91], x[57], x[56], x[55], x[45], x[44], x[43], x[54], x[53], x[52], x[30], x[29], x[28], x[108], x[107], x[106], x[105], x[48], x[47], x[46], x[33], x[32], x[31], x[69], x[68], x[67], x[42], x[41], x[40], x[24], x[23], x[22], x[87], x[86], x[85], x[84], x[83], x[82], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[196], x[195], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[179], x[178], x[177], x[405], x[3]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[196], x[195], x[188], x[187], x[190], x[189], x[186], x[185], x[184], x[183], x[194], x[193], x[192], x[191], x[179], x[178], x[177], x[165], x[164], x[163], x[123], x[122], x[159], x[158], x[170], x[169], x[168], x[198], x[197], x[167], x[166], x[162], x[161], x[160], x[27], x[26], x[25], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[176], x[175], x[174], x[173], x[172], x[171], x[30], x[29], x[28], x[146], x[145], x[121], x[120], x[119], x[141], x[140], x[139], x[182], x[181], x[180], x[144], x[143], x[142], x[33], x[32], x[31], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[24], x[23], x[22], x[126], x[125], x[124], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[241], x[240], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[222], x[221], x[220], x[406], x[3]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[196], x[195], x[188], x[187], x[190], x[189], x[186], x[185], x[184], x[183], x[194], x[193], x[192], x[191], x[179], x[178], x[177], x[165], x[164], x[163], x[123], x[122], x[159], x[158], x[170], x[169], x[168], x[198], x[197], x[167], x[166], x[162], x[161], x[160], x[27], x[26], x[25], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[176], x[175], x[174], x[173], x[172], x[171], x[30], x[29], x[28], x[146], x[145], x[121], x[120], x[119], x[141], x[140], x[139], x[182], x[181], x[180], x[144], x[143], x[142], x[33], x[32], x[31], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[24], x[23], x[22], x[126], x[125], x[124], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[241], x[240], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[222], x[221], x[220], x[406], x[3]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[188], x[187], x[159], x[158], x[123], x[122], x[186], x[185], x[190], x[189], x[196], x[195], x[152], x[151], x[165], x[164], x[163], x[141], x[140], x[139], x[198], x[197], x[194], x[193], x[148], x[147], x[121], x[120], x[119], x[162], x[161], x[160], x[150], x[149], x[167], x[166], x[184], x[183], x[192], x[191], x[170], x[169], x[168], x[179], x[178], x[177], x[27], x[26], x[25], x[146], x[145], x[135], x[134], x[133], x[154], x[153], x[182], x[181], x[180], x[176], x[175], x[174], x[30], x[29], x[28], x[129], x[128], x[127], x[132], x[131], x[130], x[144], x[143], x[142], x[157], x[156], x[155], x[173], x[172], x[171], x[33], x[32], x[31], x[126], x[125], x[124], x[138], x[137], x[136], x[24], x[23], x[22], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[278], x[277], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[262], x[261], x[260], x[407], x[3]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[188], x[187], x[159], x[158], x[123], x[122], x[186], x[185], x[190], x[189], x[196], x[195], x[152], x[151], x[165], x[164], x[163], x[141], x[140], x[139], x[198], x[197], x[194], x[193], x[148], x[147], x[121], x[120], x[119], x[162], x[161], x[160], x[150], x[149], x[167], x[166], x[184], x[183], x[192], x[191], x[170], x[169], x[168], x[179], x[178], x[177], x[27], x[26], x[25], x[146], x[145], x[135], x[134], x[133], x[154], x[153], x[182], x[181], x[180], x[176], x[175], x[174], x[30], x[29], x[28], x[129], x[128], x[127], x[132], x[131], x[130], x[144], x[143], x[142], x[157], x[156], x[155], x[173], x[172], x[171], x[33], x[32], x[31], x[126], x[125], x[124], x[138], x[137], x[136], x[24], x[23], x[22], x[6], x[5], x[4], x[9], x[8], x[7], x[15], x[14], x[13], x[278], x[277], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[262], x[261], x[260], x[407], x[3]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[152], x[151], x[190], x[189], x[159], x[158], x[148], x[147], x[154], x[153], x[184], x[183], x[192], x[191], x[167], x[166], x[198], x[197], x[196], x[195], x[188], x[187], x[194], x[193], x[135], x[134], x[133], x[123], x[122], x[170], x[169], x[168], x[141], x[140], x[139], x[186], x[185], x[27], x[26], x[25], x[129], x[128], x[127], x[138], x[137], x[136], x[157], x[156], x[155], x[146], x[145], x[150], x[149], x[173], x[172], x[171], x[144], x[143], x[142], x[182], x[181], x[180], x[179], x[178], x[177], x[165], x[164], x[163], x[30], x[29], x[28], x[176], x[175], x[174], x[121], x[120], x[119], x[162], x[161], x[160], x[6], x[5], x[4], x[33], x[32], x[31], x[126], x[125], x[124], x[132], x[131], x[130], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[274], x[273], x[254], x[253], x[252], x[408], x[3]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[152], x[151], x[190], x[189], x[159], x[158], x[148], x[147], x[154], x[153], x[184], x[183], x[192], x[191], x[167], x[166], x[198], x[197], x[196], x[195], x[188], x[187], x[194], x[193], x[135], x[134], x[133], x[123], x[122], x[170], x[169], x[168], x[141], x[140], x[139], x[186], x[185], x[27], x[26], x[25], x[129], x[128], x[127], x[138], x[137], x[136], x[157], x[156], x[155], x[146], x[145], x[150], x[149], x[173], x[172], x[171], x[144], x[143], x[142], x[182], x[181], x[180], x[179], x[178], x[177], x[165], x[164], x[163], x[30], x[29], x[28], x[176], x[175], x[174], x[121], x[120], x[119], x[162], x[161], x[160], x[6], x[5], x[4], x[33], x[32], x[31], x[126], x[125], x[124], x[132], x[131], x[130], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[274], x[273], x[254], x[253], x[252], x[408], x[3]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[188], x[187], x[184], x[183], x[192], x[191], x[123], x[122], x[159], x[158], x[194], x[193], x[167], x[166], x[146], x[145], x[190], x[189], x[154], x[153], x[165], x[164], x[163], x[186], x[185], x[152], x[151], x[148], x[147], x[157], x[156], x[155], x[173], x[172], x[171], x[150], x[149], x[121], x[120], x[119], x[27], x[26], x[25], x[198], x[197], x[196], x[195], x[141], x[140], x[139], x[176], x[175], x[174], x[144], x[143], x[142], x[126], x[125], x[124], x[30], x[29], x[28], x[170], x[169], x[168], x[138], x[137], x[136], x[162], x[161], x[160], x[135], x[134], x[133], x[129], x[128], x[127], x[132], x[131], x[130], x[6], x[5], x[4], x[33], x[32], x[31], x[182], x[181], x[180], x[179], x[178], x[177], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[272], x[271], x[251], x[250], x[249], x[409], x[3]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[188], x[187], x[184], x[183], x[192], x[191], x[123], x[122], x[159], x[158], x[194], x[193], x[167], x[166], x[146], x[145], x[190], x[189], x[154], x[153], x[165], x[164], x[163], x[186], x[185], x[152], x[151], x[148], x[147], x[157], x[156], x[155], x[173], x[172], x[171], x[150], x[149], x[121], x[120], x[119], x[27], x[26], x[25], x[198], x[197], x[196], x[195], x[141], x[140], x[139], x[176], x[175], x[174], x[144], x[143], x[142], x[126], x[125], x[124], x[30], x[29], x[28], x[170], x[169], x[168], x[138], x[137], x[136], x[162], x[161], x[160], x[135], x[134], x[133], x[129], x[128], x[127], x[132], x[131], x[130], x[6], x[5], x[4], x[33], x[32], x[31], x[182], x[181], x[180], x[179], x[178], x[177], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[272], x[271], x[251], x[250], x[249], x[409], x[3]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[276], x[275], x[282], x[281], x[280], x[279], x[274], x[273], x[272], x[271], x[270], x[269], x[259], x[258], x[257], x[256], x[255], x[268], x[267], x[266], x[265], x[264], x[263], x[254], x[253], x[252], x[278], x[277], x[248], x[247], x[251], x[250], x[249], x[246], x[245], x[244], x[27], x[26], x[25], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[207], x[206], x[230], x[229], x[30], x[29], x[28], x[262], x[261], x[260], x[228], x[227], x[226], x[6], x[5], x[4], x[33], x[32], x[31], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[205], x[204], x[203], x[210], x[209], x[208], x[9], x[8], x[7], x[24], x[23], x[22], x[15], x[14], x[13], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[311], x[310], x[294], x[293], x[292], x[410], x[3]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[276], x[275], x[282], x[281], x[280], x[279], x[274], x[273], x[272], x[271], x[270], x[269], x[259], x[258], x[257], x[256], x[255], x[268], x[267], x[266], x[265], x[264], x[263], x[254], x[253], x[252], x[278], x[277], x[248], x[247], x[251], x[250], x[249], x[246], x[245], x[244], x[27], x[26], x[25], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[207], x[206], x[230], x[229], x[30], x[29], x[28], x[262], x[261], x[260], x[228], x[227], x[226], x[6], x[5], x[4], x[33], x[32], x[31], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[205], x[204], x[203], x[210], x[209], x[208], x[9], x[8], x[7], x[24], x[23], x[22], x[15], x[14], x[13], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[311], x[310], x[294], x[293], x[292], x[410], x[3]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[259], x[258], x[270], x[269], x[230], x[229], x[282], x[281], x[274], x[273], x[239], x[238], x[207], x[206], x[276], x[275], x[280], x[279], x[278], x[277], x[272], x[271], x[243], x[242], x[235], x[234], x[233], x[232], x[231], x[246], x[245], x[244], x[237], x[236], x[248], x[247], x[210], x[209], x[208], x[268], x[267], x[266], x[254], x[253], x[252], x[27], x[26], x[25], x[219], x[218], x[217], x[205], x[204], x[203], x[257], x[256], x[255], x[265], x[264], x[263], x[241], x[240], x[262], x[261], x[260], x[251], x[250], x[249], x[30], x[29], x[28], x[225], x[224], x[223], x[213], x[212], x[211], x[216], x[215], x[214], x[228], x[227], x[226], x[6], x[5], x[4], x[33], x[32], x[31], x[222], x[221], x[220], x[9], x[8], x[7], x[24], x[23], x[22], x[15], x[14], x[13], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[360], x[359], x[339], x[338], x[337], x[411], x[3]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[259], x[258], x[270], x[269], x[230], x[229], x[282], x[281], x[274], x[273], x[239], x[238], x[207], x[206], x[276], x[275], x[280], x[279], x[278], x[277], x[272], x[271], x[243], x[242], x[235], x[234], x[233], x[232], x[231], x[246], x[245], x[244], x[237], x[236], x[248], x[247], x[210], x[209], x[208], x[268], x[267], x[266], x[254], x[253], x[252], x[27], x[26], x[25], x[219], x[218], x[217], x[205], x[204], x[203], x[257], x[256], x[255], x[265], x[264], x[263], x[241], x[240], x[262], x[261], x[260], x[251], x[250], x[249], x[30], x[29], x[28], x[225], x[224], x[223], x[213], x[212], x[211], x[216], x[215], x[214], x[228], x[227], x[226], x[6], x[5], x[4], x[33], x[32], x[31], x[222], x[221], x[220], x[9], x[8], x[7], x[24], x[23], x[22], x[15], x[14], x[13], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[360], x[359], x[339], x[338], x[337], x[411], x[3]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[276], x[275], x[239], x[238], x[280], x[279], x[274], x[273], x[235], x[234], x[241], x[240], x[282], x[281], x[248], x[247], x[278], x[277], x[230], x[229], x[257], x[256], x[255], x[243], x[242], x[219], x[218], x[217], x[265], x[264], x[263], x[254], x[253], x[252], x[272], x[271], x[259], x[258], x[270], x[269], x[27], x[26], x[25], x[213], x[212], x[211], x[222], x[221], x[220], x[268], x[267], x[266], x[237], x[236], x[207], x[206], x[228], x[227], x[226], x[262], x[261], x[260], x[210], x[209], x[208], x[30], x[29], x[28], x[225], x[224], x[223], x[251], x[250], x[249], x[233], x[232], x[231], x[246], x[245], x[244], x[6], x[5], x[4], x[33], x[32], x[31], x[216], x[215], x[214], x[205], x[204], x[203], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[351], x[350], x[322], x[321], x[320], x[412], x[3]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[276], x[275], x[239], x[238], x[280], x[279], x[274], x[273], x[235], x[234], x[241], x[240], x[282], x[281], x[248], x[247], x[278], x[277], x[230], x[229], x[257], x[256], x[255], x[243], x[242], x[219], x[218], x[217], x[265], x[264], x[263], x[254], x[253], x[252], x[272], x[271], x[259], x[258], x[270], x[269], x[27], x[26], x[25], x[213], x[212], x[211], x[222], x[221], x[220], x[268], x[267], x[266], x[237], x[236], x[207], x[206], x[228], x[227], x[226], x[262], x[261], x[260], x[210], x[209], x[208], x[30], x[29], x[28], x[225], x[224], x[223], x[251], x[250], x[249], x[233], x[232], x[231], x[246], x[245], x[244], x[6], x[5], x[4], x[33], x[32], x[31], x[216], x[215], x[214], x[205], x[204], x[203], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[351], x[350], x[322], x[321], x[320], x[412], x[3]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[276], x[275], x[280], x[279], x[282], x[281], x[243], x[242], x[259], x[258], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[207], x[206], x[274], x[273], x[241], x[240], x[230], x[229], x[270], x[269], x[268], x[267], x[266], x[239], x[238], x[235], x[234], x[225], x[224], x[223], x[237], x[236], x[27], x[26], x[25], x[278], x[277], x[233], x[232], x[231], x[228], x[227], x[226], x[205], x[204], x[203], x[30], x[29], x[28], x[254], x[253], x[252], x[272], x[271], x[222], x[221], x[220], x[210], x[209], x[208], x[246], x[245], x[244], x[219], x[218], x[217], x[213], x[212], x[211], x[216], x[215], x[214], x[33], x[32], x[31], x[6], x[5], x[4], x[262], x[261], x[260], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[251], x[250], x[249], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[358], x[357], x[336], x[335], x[334], x[413], x[3]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[276], x[275], x[280], x[279], x[282], x[281], x[243], x[242], x[259], x[258], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[207], x[206], x[274], x[273], x[241], x[240], x[230], x[229], x[270], x[269], x[268], x[267], x[266], x[239], x[238], x[235], x[234], x[225], x[224], x[223], x[237], x[236], x[27], x[26], x[25], x[278], x[277], x[233], x[232], x[231], x[228], x[227], x[226], x[205], x[204], x[203], x[30], x[29], x[28], x[254], x[253], x[252], x[272], x[271], x[222], x[221], x[220], x[210], x[209], x[208], x[246], x[245], x[244], x[219], x[218], x[217], x[213], x[212], x[211], x[216], x[215], x[214], x[33], x[32], x[31], x[6], x[5], x[4], x[262], x[261], x[260], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[251], x[250], x[249], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[358], x[357], x[336], x[335], x[334], x[413], x[3]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[364], x[363], x[366], x[365], x[358], x[357], x[356], x[355], x[347], x[346], x[362], x[361], x[351], x[350], x[349], x[348], x[345], x[344], x[343], x[333], x[332], x[331], x[330], x[329], x[328], x[354], x[353], x[352], x[336], x[335], x[334], x[327], x[326], x[325], x[27], x[26], x[25], x[324], x[323], x[316], x[315], x[314], x[291], x[290], x[313], x[312], x[342], x[341], x[340], x[322], x[321], x[320], x[360], x[359], x[319], x[318], x[317], x[30], x[29], x[28], x[311], x[310], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[6], x[5], x[4], x[33], x[32], x[31], x[300], x[299], x[298], x[289], x[288], x[287], x[297], x[296], x[295], x[339], x[338], x[337], x[15], x[14], x[13], x[24], x[23], x[22], x[9], x[8], x[7], x[294], x[293], x[292], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[59], x[58], x[42], x[41], x[40], x[414], x[3]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[364], x[363], x[366], x[365], x[358], x[357], x[356], x[355], x[347], x[346], x[362], x[361], x[351], x[350], x[349], x[348], x[345], x[344], x[343], x[333], x[332], x[331], x[330], x[329], x[328], x[354], x[353], x[352], x[336], x[335], x[334], x[327], x[326], x[325], x[27], x[26], x[25], x[324], x[323], x[316], x[315], x[314], x[291], x[290], x[313], x[312], x[342], x[341], x[340], x[322], x[321], x[320], x[360], x[359], x[319], x[318], x[317], x[30], x[29], x[28], x[311], x[310], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[6], x[5], x[4], x[33], x[32], x[31], x[300], x[299], x[298], x[289], x[288], x[287], x[297], x[296], x[295], x[339], x[338], x[337], x[15], x[14], x[13], x[24], x[23], x[22], x[9], x[8], x[7], x[294], x[293], x[292], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[59], x[58], x[42], x[41], x[40], x[414], x[3]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[333], x[332], x[347], x[346], x[356], x[355], x[313], x[312], x[366], x[365], x[329], x[328], x[291], x[290], x[331], x[330], x[349], x[348], x[364], x[363], x[351], x[350], x[358], x[357], x[324], x[323], x[309], x[308], x[307], x[316], x[315], x[314], x[327], x[326], x[325], x[362], x[361], x[297], x[296], x[295], x[360], x[359], x[354], x[353], x[352], x[27], x[26], x[25], x[303], x[302], x[301], x[289], x[288], x[287], x[306], x[305], x[304], x[319], x[318], x[317], x[345], x[344], x[343], x[322], x[321], x[320], x[336], x[335], x[334], x[30], x[29], x[28], x[300], x[299], x[298], x[342], x[341], x[340], x[311], x[310], x[339], x[338], x[337], x[6], x[5], x[4], x[33], x[32], x[31], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[294], x[293], x[292], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[108], x[107], x[87], x[86], x[85], x[415], x[3]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[333], x[332], x[347], x[346], x[356], x[355], x[313], x[312], x[366], x[365], x[329], x[328], x[291], x[290], x[331], x[330], x[349], x[348], x[364], x[363], x[351], x[350], x[358], x[357], x[324], x[323], x[309], x[308], x[307], x[316], x[315], x[314], x[327], x[326], x[325], x[362], x[361], x[297], x[296], x[295], x[360], x[359], x[354], x[353], x[352], x[27], x[26], x[25], x[303], x[302], x[301], x[289], x[288], x[287], x[306], x[305], x[304], x[319], x[318], x[317], x[345], x[344], x[343], x[322], x[321], x[320], x[336], x[335], x[334], x[30], x[29], x[28], x[300], x[299], x[298], x[342], x[341], x[340], x[311], x[310], x[339], x[338], x[337], x[6], x[5], x[4], x[33], x[32], x[31], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[294], x[293], x[292], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[108], x[107], x[87], x[86], x[85], x[415], x[3]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[333], x[332], x[329], x[328], x[364], x[363], x[349], x[348], x[366], x[365], x[309], x[308], x[307], x[362], x[361], x[351], x[350], x[313], x[312], x[303], x[302], x[301], x[311], x[310], x[345], x[344], x[343], x[324], x[323], x[331], x[330], x[319], x[318], x[317], x[360], x[359], x[358], x[357], x[347], x[346], x[356], x[355], x[27], x[26], x[25], x[354], x[353], x[352], x[291], x[290], x[342], x[341], x[340], x[322], x[321], x[320], x[297], x[296], x[295], x[30], x[29], x[28], x[294], x[293], x[292], x[300], x[299], x[298], x[306], x[305], x[304], x[339], x[338], x[337], x[336], x[335], x[334], x[316], x[315], x[314], x[327], x[326], x[325], x[6], x[5], x[4], x[33], x[32], x[31], x[289], x[288], x[287], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[100], x[99], x[69], x[68], x[67], x[416], x[3]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[333], x[332], x[329], x[328], x[364], x[363], x[349], x[348], x[366], x[365], x[309], x[308], x[307], x[362], x[361], x[351], x[350], x[313], x[312], x[303], x[302], x[301], x[311], x[310], x[345], x[344], x[343], x[324], x[323], x[331], x[330], x[319], x[318], x[317], x[360], x[359], x[358], x[357], x[347], x[346], x[356], x[355], x[27], x[26], x[25], x[354], x[353], x[352], x[291], x[290], x[342], x[341], x[340], x[322], x[321], x[320], x[297], x[296], x[295], x[30], x[29], x[28], x[294], x[293], x[292], x[300], x[299], x[298], x[306], x[305], x[304], x[339], x[338], x[337], x[336], x[335], x[334], x[316], x[315], x[314], x[327], x[326], x[325], x[6], x[5], x[4], x[33], x[32], x[31], x[289], x[288], x[287], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[100], x[99], x[69], x[68], x[67], x[416], x[3]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[364], x[363], x[366], x[365], x[349], x[348], x[324], x[323], x[362], x[361], x[347], x[346], x[333], x[332], x[329], x[328], x[345], x[344], x[343], x[331], x[330], x[291], x[290], x[313], x[312], x[356], x[355], x[354], x[353], x[352], x[319], x[318], x[317], x[300], x[299], x[298], x[342], x[341], x[340], x[27], x[26], x[25], x[351], x[350], x[311], x[310], x[316], x[315], x[314], x[309], x[308], x[307], x[303], x[302], x[301], x[306], x[305], x[304], x[289], x[288], x[287], x[30], x[29], x[28], x[360], x[359], x[358], x[357], x[297], x[296], x[295], x[327], x[326], x[325], x[6], x[5], x[4], x[33], x[32], x[31], x[322], x[321], x[320], x[294], x[293], x[292], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[339], x[338], x[337], x[336], x[335], x[334], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[106], x[105], x[84], x[83], x[82], x[417], x[3]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[364], x[363], x[366], x[365], x[349], x[348], x[324], x[323], x[362], x[361], x[347], x[346], x[333], x[332], x[329], x[328], x[345], x[344], x[343], x[331], x[330], x[291], x[290], x[313], x[312], x[356], x[355], x[354], x[353], x[352], x[319], x[318], x[317], x[300], x[299], x[298], x[342], x[341], x[340], x[27], x[26], x[25], x[351], x[350], x[311], x[310], x[316], x[315], x[314], x[309], x[308], x[307], x[303], x[302], x[301], x[306], x[305], x[304], x[289], x[288], x[287], x[30], x[29], x[28], x[360], x[359], x[358], x[357], x[297], x[296], x[295], x[327], x[326], x[325], x[6], x[5], x[4], x[33], x[32], x[31], x[322], x[321], x[320], x[294], x[293], x[292], x[9], x[8], x[7], x[15], x[14], x[13], x[24], x[23], x[22], x[339], x[338], x[337], x[336], x[335], x[334], x[21], x[20], x[19], x[12], x[11], x[10], x[18], x[17], x[16], x[106], x[105], x[84], x[83], x[82], x[417], x[3]}), .y(y[151]));
endmodule

