/* modified netlist. Source: module LED in file ../CaseStudies/11_LED_round_based_encryption/FPGA_based/LED_synthesis.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module LED_GHPC_ClockGating_d1 (CLK, IN_reset, IN_plaintext_s0, IN_key_s0, IN_key_s1, IN_plaintext_s1, Fresh, OUT_done, OUT_ciphertext_s0, OUT_ciphertext_s1, Synch);
    input CLK ;
    input IN_reset ;
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input [127:0] IN_key_s1 ;
    input [63:0] IN_plaintext_s1 ;
    input [63:0] Fresh ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s0 ;
    output [63:0] OUT_ciphertext_s1 ;
    output Synch ;
    wire \LED_128_Instance/addkey1_265 ;
    wire \LED_128_Instance/roundconstant[5]_roundconstant[4]_XOR_7_o ;
    wire \LED_128_Instance/addkey ;
    wire \LED_128_Instance/roundconstant_001001 ;
    wire \LED_128_Instance/ks[3]_INV_6_o ;
    wire [54:3] \LED_128_Instance/addconst_out ;
    wire N2 ;
    wire N4 ;
    wire N6 ;
    wire N8 ;
    wire N12 ;
    wire N14 ;
    wire N16 ;
    wire N18 ;
    wire N20 ;
    wire N22 ;
    wire N24 ;
    wire N26 ;
    wire N28 ;
    wire N32 ;
    wire N34 ;
    wire N36 ;
    wire N38 ;
    wire N40 ;
    wire N42 ;
    wire N44 ;
    wire N46 ;
    wire N48 ;
    wire N52 ;
    wire N54 ;
    wire N56 ;
    wire N58 ;
    wire N60 ;
    wire N62 ;
    wire N64 ;
    wire N66 ;
    wire N68 ;
    wire N72 ;
    wire N74 ;
    wire N76 ;
    wire N78 ;
    wire N80 ;
    wire internal_done_glue_set_843 ;
    wire N82 ;
    wire N84 ;
    wire N86 ;
    wire N88 ;
    wire N90 ;
    wire N92 ;
    wire N94 ;
    wire N96 ;
    wire N98 ;
    wire N100 ;
    wire N102 ;
    wire N104 ;
    wire [5:0] \LED_128_Instance/roundconstant ;
    wire [63:0] \LED_128_Instance/mixcolumns_out ;
    wire [63:0] \LED_128_Instance/subcells_out ;
    wire [63:0] \LED_128_Instance/addroundkey_out ;
    wire [3:0] \LED_128_Instance/ks ;
    wire [63:0] \LED_128_Instance/state ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_869 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_901 ;
    wire new_AGEMA_signal_905 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_913 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_921 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1439 ;
    wire clk_gated ;

    /* cells in depth 0 */
    LUT6 #( .INIT ( 64'h0000001000000000 ) ) \GND_3_o_roundconstant[5]_equal_1_o<5>1 ( .I0 (\LED_128_Instance/roundconstant [5]), .I1 (\LED_128_Instance/roundconstant [4]), .I2 (\LED_128_Instance/roundconstant [3]), .I3 (\LED_128_Instance/roundconstant [2]), .I4 (\LED_128_Instance/roundconstant [1]), .I5 (\LED_128_Instance/roundconstant [0]), .O (\LED_128_Instance/roundconstant_001001 ) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[9].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[73], IN_key_s0[73]}), .I1 ({IN_key_s1[9], IN_key_s0[9]}), .I2 ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[8].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[72], IN_key_s0[72]}), .I1 ({IN_key_s1[8], IN_key_s0[8]}), .I2 ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[7].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[71], IN_key_s0[71]}), .I1 ({IN_key_s1[7], IN_key_s0[7]}), .I2 ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[63].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[127], IN_key_s0[127]}), .I1 ({IN_key_s1[63], IN_key_s0[63]}), .I2 ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[62].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[126], IN_key_s0[126]}), .I1 ({IN_key_s1[62], IN_key_s0[62]}), .I2 ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[61].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[125], IN_key_s0[125]}), .I1 ({IN_key_s1[61], IN_key_s0[61]}), .I2 ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[60].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[124], IN_key_s0[124]}), .I1 ({IN_key_s1[60], IN_key_s0[60]}), .I2 ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[59].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[123], IN_key_s0[123]}), .I1 ({IN_key_s1[59], IN_key_s0[59]}), .I2 ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[58].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[122], IN_key_s0[122]}), .I1 ({IN_key_s1[58], IN_key_s0[58]}), .I2 ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[57].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[121], IN_key_s0[121]}), .I1 ({IN_key_s1[57], IN_key_s0[57]}), .I2 ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[56].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[120], IN_key_s0[120]}), .I1 ({IN_key_s1[56], IN_key_s0[56]}), .I2 ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[55].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[119], IN_key_s0[119]}), .I1 ({IN_key_s1[55], IN_key_s0[55]}), .I2 ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[51].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[115], IN_key_s0[115]}), .I1 ({IN_key_s1[51], IN_key_s0[51]}), .I2 ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[50].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[114], IN_key_s0[114]}), .I1 ({IN_key_s1[50], IN_key_s0[50]}), .I2 ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[47].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[111], IN_key_s0[111]}), .I1 ({IN_key_s1[47], IN_key_s0[47]}), .I2 ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[46].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[110], IN_key_s0[110]}), .I1 ({IN_key_s1[46], IN_key_s0[46]}), .I2 ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[45].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[109], IN_key_s0[109]}), .I1 ({IN_key_s1[45], IN_key_s0[45]}), .I2 ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[44].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[108], IN_key_s0[108]}), .I1 ({IN_key_s1[44], IN_key_s0[44]}), .I2 ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[43].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[107], IN_key_s0[107]}), .I1 ({IN_key_s1[43], IN_key_s0[43]}), .I2 ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[42].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[106], IN_key_s0[106]}), .I1 ({IN_key_s1[42], IN_key_s0[42]}), .I2 ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[41].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[105], IN_key_s0[105]}), .I1 ({IN_key_s1[41], IN_key_s0[41]}), .I2 ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[40].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[104], IN_key_s0[104]}), .I1 ({IN_key_s1[40], IN_key_s0[40]}), .I2 ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[39].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[103], IN_key_s0[103]}), .I1 ({IN_key_s1[39], IN_key_s0[39]}), .I2 ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[35].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[99], IN_key_s0[99]}), .I1 ({IN_key_s1[35], IN_key_s0[35]}), .I2 ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[34].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[98], IN_key_s0[98]}), .I1 ({IN_key_s1[34], IN_key_s0[34]}), .I2 ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[32].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[96], IN_key_s0[96]}), .I1 ({IN_key_s1[32], IN_key_s0[32]}), .I2 ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[31].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[95], IN_key_s0[95]}), .I1 ({IN_key_s1[31], IN_key_s0[31]}), .I2 ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[30].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[94], IN_key_s0[94]}), .I1 ({IN_key_s1[30], IN_key_s0[30]}), .I2 ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[2].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[66], IN_key_s0[66]}), .I1 ({IN_key_s1[2], IN_key_s0[2]}), .I2 ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[29].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[93], IN_key_s0[93]}), .I1 ({IN_key_s1[29], IN_key_s0[29]}), .I2 ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[28].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[92], IN_key_s0[92]}), .I1 ({IN_key_s1[28], IN_key_s0[28]}), .I2 ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[27].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[91], IN_key_s0[91]}), .I1 ({IN_key_s1[27], IN_key_s0[27]}), .I2 ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[26].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[90], IN_key_s0[90]}), .I1 ({IN_key_s1[26], IN_key_s0[26]}), .I2 ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[25].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[89], IN_key_s0[89]}), .I1 ({IN_key_s1[25], IN_key_s0[25]}), .I2 ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[24].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[88], IN_key_s0[88]}), .I1 ({IN_key_s1[24], IN_key_s0[24]}), .I2 ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[23].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[87], IN_key_s0[87]}), .I1 ({IN_key_s1[23], IN_key_s0[23]}), .I2 ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[1].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[65], IN_key_s0[65]}), .I1 ({IN_key_s1[1], IN_key_s0[1]}), .I2 ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[18].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[82], IN_key_s0[82]}), .I1 ({IN_key_s1[18], IN_key_s0[18]}), .I2 ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[17].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[81], IN_key_s0[81]}), .I1 ({IN_key_s1[17], IN_key_s0[17]}), .I2 ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[15].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[79], IN_key_s0[79]}), .I1 ({IN_key_s1[15], IN_key_s0[15]}), .I2 ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[14].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[78], IN_key_s0[78]}), .I1 ({IN_key_s1[14], IN_key_s0[14]}), .I2 ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[13].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[77], IN_key_s0[77]}), .I1 ({IN_key_s1[13], IN_key_s0[13]}), .I2 ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[12].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[76], IN_key_s0[76]}), .I1 ({IN_key_s1[12], IN_key_s0[12]}), .I2 ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[11].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[75], IN_key_s0[75]}), .I1 ({IN_key_s1[11], IN_key_s0[11]}), .I2 ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[10].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[74], IN_key_s0[74]}), .I1 ({IN_key_s1[10], IN_key_s0[10]}), .I2 ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[0].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[64], IN_key_s0[64]}), .I1 ({IN_key_s1[0], IN_key_s0[0]}), .I2 ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[6].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[6], IN_key_s0[6]}), .I3 ({IN_key_s1[70], IN_key_s0[70]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1049, \LED_128_Instance/addroundkey_out [6]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[5].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[5], IN_key_s0[5]}), .I3 ({IN_key_s1[69], IN_key_s0[69]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1053, \LED_128_Instance/addroundkey_out [5]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[54].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[54], IN_key_s0[54]}), .I3 ({IN_key_s1[118], IN_key_s0[118]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1057, \LED_128_Instance/addroundkey_out [54]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[53].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[53], IN_key_s0[53]}), .I3 ({IN_key_s1[117], IN_key_s0[117]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1061, \LED_128_Instance/addroundkey_out [53]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[52].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[52], IN_key_s0[52]}), .I3 ({IN_key_s1[116], IN_key_s0[116]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1065, \LED_128_Instance/addroundkey_out [52]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[4].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[4], IN_key_s0[4]}), .I3 ({IN_key_s1[68], IN_key_s0[68]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1069, \LED_128_Instance/addroundkey_out [4]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[49].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[49], IN_key_s0[49]}), .I3 ({IN_key_s1[113], IN_key_s0[113]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1073, \LED_128_Instance/addroundkey_out [49]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[48].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[48], IN_key_s0[48]}), .I3 ({IN_key_s1[112], IN_key_s0[112]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1077, \LED_128_Instance/addroundkey_out [48]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[3].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[3], IN_key_s0[3]}), .I3 ({IN_key_s1[67], IN_key_s0[67]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1081, \LED_128_Instance/addroundkey_out [3]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[38].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[38], IN_key_s0[38]}), .I3 ({IN_key_s1[102], IN_key_s0[102]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1085, \LED_128_Instance/addroundkey_out [38]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[37].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[37], IN_key_s0[37]}), .I3 ({IN_key_s1[101], IN_key_s0[101]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1089, \LED_128_Instance/addroundkey_out [37]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[36].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[36], IN_key_s0[36]}), .I3 ({IN_key_s1[100], IN_key_s0[100]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1093, \LED_128_Instance/addroundkey_out [36]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[33].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[33], IN_key_s0[33]}), .I3 ({IN_key_s1[97], IN_key_s0[97]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1097, \LED_128_Instance/addroundkey_out [33]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[22].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[22], IN_key_s0[22]}), .I3 ({IN_key_s1[86], IN_key_s0[86]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1101, \LED_128_Instance/addroundkey_out [22]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[21].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[21], IN_key_s0[21]}), .I3 ({IN_key_s1[85], IN_key_s0[85]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1105, \LED_128_Instance/addroundkey_out [21]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[20].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[20], IN_key_s0[20]}), .I3 ({IN_key_s1[84], IN_key_s0[84]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1109, \LED_128_Instance/addroundkey_out [20]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[19].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[19], IN_key_s0[19]}), .I3 ({IN_key_s1[83], IN_key_s0[83]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1113, \LED_128_Instance/addroundkey_out [19]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[16].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[16], IN_key_s0[16]}), .I3 ({IN_key_s1[80], IN_key_s0[80]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1117, \LED_128_Instance/addroundkey_out [16]}) ) ;
    LUT4 #( .INIT ( 16'h8001 ) ) \LED_128_Instance/addkey1 ( .I0 (\LED_128_Instance/ks [0]), .I1 (\LED_128_Instance/ks [1]), .I2 (\LED_128_Instance/ks [2]), .I3 (\LED_128_Instance/ks [3]), .O (\LED_128_Instance/addkey ) ) ;
    LUT4 #( .INIT ( 16'h0001 ) ) \LED_128_Instance/addkey21 ( .I0 (\LED_128_Instance/ks [3]), .I1 (\LED_128_Instance/ks [2]), .I2 (\LED_128_Instance/ks [1]), .I3 (\LED_128_Instance/ks [0]), .O (\LED_128_Instance/addkey1_265 ) ) ;
    LUT2 #( .INIT ( 4'h9 ) ) \LED_128_Instance/Mxor_roundconstant[5]_roundconstant[4]_XOR_7_o_xo<0>1 ( .I0 (\LED_128_Instance/roundconstant [4]), .I1 (\LED_128_Instance/roundconstant [5]), .O (\LED_128_Instance/roundconstant[5]_roundconstant[4]_XOR_7_o ) ) ;
    LUT2 #( .INIT ( 4'hE ) ) internal_done_glue_set ( .I0 (OUT_done), .I1 (\LED_128_Instance/roundconstant_001001 ), .O (internal_done_glue_set_843) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<3:0>_3_xo<0>1 ( .I0 ({IN_key_s1[3], IN_key_s0[3]}), .I1 ({IN_key_s1[67], IN_key_s0[67]}), .I2 ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1118, \LED_128_Instance/addconst_out [3]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<35:32>_1_xo<0>1 ( .I0 ({IN_key_s1[33], IN_key_s0[33]}), .I1 ({IN_key_s1[97], IN_key_s0[97]}), .I2 ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1119, \LED_128_Instance/addconst_out [33]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<19:16>_3_xo<0>1 ( .I0 ({IN_key_s1[19], IN_key_s0[19]}), .I1 ({IN_key_s1[83], IN_key_s0[83]}), .I2 ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1120, \LED_128_Instance/addconst_out [19]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<19:16>_0_xo<0>1 ( .I0 ({IN_key_s1[16], IN_key_s0[16]}), .I1 ({IN_key_s1[80], IN_key_s0[80]}), .I2 ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1121, \LED_128_Instance/addconst_out [16]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<38:36>_2_xo<0>1 ( .I0 ({IN_key_s1[38], IN_key_s0[38]}), .I1 ({IN_key_s1[102], IN_key_s0[102]}), .I2 ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [5]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1122, \LED_128_Instance/addconst_out [38]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<38:36>_1_xo<0>1 ( .I0 ({IN_key_s1[37], IN_key_s0[37]}), .I1 ({IN_key_s1[101], IN_key_s0[101]}), .I2 ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [4]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1123, \LED_128_Instance/addconst_out [37]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<38:36>_0_xo<0>1 ( .I0 ({IN_key_s1[36], IN_key_s0[36]}), .I1 ({IN_key_s1[100], IN_key_s0[100]}), .I2 ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [3]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1124, \LED_128_Instance/addconst_out [36]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<6:4>_2_xo<0>1 ( .I0 ({IN_key_s1[6], IN_key_s0[6]}), .I1 ({IN_key_s1[70], IN_key_s0[70]}), .I2 ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [5]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1125, \LED_128_Instance/addconst_out [6]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<6:4>_1_xo<0>1 ( .I0 ({IN_key_s1[5], IN_key_s0[5]}), .I1 ({IN_key_s1[69], IN_key_s0[69]}), .I2 ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [4]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1126, \LED_128_Instance/addconst_out [5]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<6:4>_0_xo<0>1 ( .I0 ({IN_key_s1[4], IN_key_s0[4]}), .I1 ({IN_key_s1[68], IN_key_s0[68]}), .I2 ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [3]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1127, \LED_128_Instance/addconst_out [4]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<51:48>_1_xo<0>1 ( .I0 ({IN_key_s1[49], IN_key_s0[49]}), .I1 ({IN_key_s1[113], IN_key_s0[113]}), .I2 ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1128, \LED_128_Instance/addconst_out [49]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<51:48>_0_xo<0>1 ( .I0 ({IN_key_s1[48], IN_key_s0[48]}), .I1 ({IN_key_s1[112], IN_key_s0[112]}), .I2 ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1129, \LED_128_Instance/addconst_out [48]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<54:52>_2_xo<0>1 ( .I0 ({IN_key_s1[54], IN_key_s0[54]}), .I1 ({IN_key_s1[118], IN_key_s0[118]}), .I2 ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [2]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1130, \LED_128_Instance/addconst_out [54]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<54:52>_1_xo<0>1 ( .I0 ({IN_key_s1[53], IN_key_s0[53]}), .I1 ({IN_key_s1[117], IN_key_s0[117]}), .I2 ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [1]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1131, \LED_128_Instance/addconst_out [53]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<54:52>_0_xo<0>1 ( .I0 ({IN_key_s1[52], IN_key_s0[52]}), .I1 ({IN_key_s1[116], IN_key_s0[116]}), .I2 ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [0]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1132, \LED_128_Instance/addconst_out [52]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<22:20>_2_xo<0>1 ( .I0 ({IN_key_s1[22], IN_key_s0[22]}), .I1 ({IN_key_s1[86], IN_key_s0[86]}), .I2 ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [2]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1133, \LED_128_Instance/addconst_out [22]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<22:20>_1_xo<0>1 ( .I0 ({IN_key_s1[21], IN_key_s0[21]}), .I1 ({IN_key_s1[85], IN_key_s0[85]}), .I2 ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [1]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1134, \LED_128_Instance/addconst_out [21]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<22:20>_0_xo<0>1 ( .I0 ({IN_key_s1[20], IN_key_s0[20]}), .I1 ({IN_key_s1[84], IN_key_s0[84]}), .I2 ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [0]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1135, \LED_128_Instance/addconst_out [20]}) ) ;
    INV \LED_128_Instance/ks[3]_INV_6_o1_INV_0 ( .I (\LED_128_Instance/ks [3]), .O (\LED_128_Instance/ks[3]_INV_6_o ) ) ;
    ClockGatingController #(3) ClockGatingInst ( .clk (CLK), .rst (IN_reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[0].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}), .I1 ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}), .I2 ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}), .I3 ({new_AGEMA_signal_1118, \LED_128_Instance/addconst_out [3]}), .clk (CLK), .r (Fresh[0]), .O ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[0].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}), .I1 ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}), .I2 ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}), .I3 ({new_AGEMA_signal_1118, \LED_128_Instance/addconst_out [3]}), .clk (CLK), .r (Fresh[1]), .O ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[0].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}), .I1 ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}), .I2 ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}), .I3 ({new_AGEMA_signal_1118, \LED_128_Instance/addconst_out [3]}), .clk (CLK), .r (Fresh[2]), .O ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[0].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}), .I1 ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}), .I2 ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}), .I3 ({new_AGEMA_signal_1118, \LED_128_Instance/addconst_out [3]}), .clk (CLK), .r (Fresh[3]), .O ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[1].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1127, \LED_128_Instance/addconst_out [4]}), .I1 ({new_AGEMA_signal_1126, \LED_128_Instance/addconst_out [5]}), .I2 ({new_AGEMA_signal_1125, \LED_128_Instance/addconst_out [6]}), .I3 ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}), .clk (CLK), .r (Fresh[4]), .O ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[1].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1127, \LED_128_Instance/addconst_out [4]}), .I1 ({new_AGEMA_signal_1126, \LED_128_Instance/addconst_out [5]}), .I2 ({new_AGEMA_signal_1125, \LED_128_Instance/addconst_out [6]}), .I3 ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}), .clk (CLK), .r (Fresh[5]), .O ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[1].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1127, \LED_128_Instance/addconst_out [4]}), .I1 ({new_AGEMA_signal_1126, \LED_128_Instance/addconst_out [5]}), .I2 ({new_AGEMA_signal_1125, \LED_128_Instance/addconst_out [6]}), .I3 ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}), .clk (CLK), .r (Fresh[6]), .O ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[1].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1127, \LED_128_Instance/addconst_out [4]}), .I1 ({new_AGEMA_signal_1126, \LED_128_Instance/addconst_out [5]}), .I2 ({new_AGEMA_signal_1125, \LED_128_Instance/addconst_out [6]}), .I3 ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}), .clk (CLK), .r (Fresh[7]), .O ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[2].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}), .I1 ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}), .I2 ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}), .I3 ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}), .clk (CLK), .r (Fresh[8]), .O ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[2].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}), .I1 ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}), .I2 ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}), .I3 ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}), .clk (CLK), .r (Fresh[9]), .O ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[2].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}), .I1 ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}), .I2 ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}), .I3 ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}), .clk (CLK), .r (Fresh[10]), .O ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[2].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}), .I1 ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}), .I2 ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}), .I3 ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}), .clk (CLK), .r (Fresh[11]), .O ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[3].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}), .I1 ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}), .I2 ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}), .I3 ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}), .clk (CLK), .r (Fresh[12]), .O ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[3].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}), .I1 ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}), .I2 ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}), .I3 ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}), .clk (CLK), .r (Fresh[13]), .O ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[3].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}), .I1 ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}), .I2 ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}), .I3 ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}), .clk (CLK), .r (Fresh[14]), .O ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[3].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}), .I1 ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}), .I2 ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}), .I3 ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}), .clk (CLK), .r (Fresh[15]), .O ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[4].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1121, \LED_128_Instance/addconst_out [16]}), .I1 ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}), .I2 ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}), .I3 ({new_AGEMA_signal_1120, \LED_128_Instance/addconst_out [19]}), .clk (CLK), .r (Fresh[16]), .O ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[4].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1121, \LED_128_Instance/addconst_out [16]}), .I1 ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}), .I2 ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}), .I3 ({new_AGEMA_signal_1120, \LED_128_Instance/addconst_out [19]}), .clk (CLK), .r (Fresh[17]), .O ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[4].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1121, \LED_128_Instance/addconst_out [16]}), .I1 ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}), .I2 ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}), .I3 ({new_AGEMA_signal_1120, \LED_128_Instance/addconst_out [19]}), .clk (CLK), .r (Fresh[18]), .O ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[4].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1121, \LED_128_Instance/addconst_out [16]}), .I1 ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}), .I2 ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}), .I3 ({new_AGEMA_signal_1120, \LED_128_Instance/addconst_out [19]}), .clk (CLK), .r (Fresh[19]), .O ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[5].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1135, \LED_128_Instance/addconst_out [20]}), .I1 ({new_AGEMA_signal_1134, \LED_128_Instance/addconst_out [21]}), .I2 ({new_AGEMA_signal_1133, \LED_128_Instance/addconst_out [22]}), .I3 ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}), .clk (CLK), .r (Fresh[20]), .O ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[5].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1135, \LED_128_Instance/addconst_out [20]}), .I1 ({new_AGEMA_signal_1134, \LED_128_Instance/addconst_out [21]}), .I2 ({new_AGEMA_signal_1133, \LED_128_Instance/addconst_out [22]}), .I3 ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}), .clk (CLK), .r (Fresh[21]), .O ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[5].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1135, \LED_128_Instance/addconst_out [20]}), .I1 ({new_AGEMA_signal_1134, \LED_128_Instance/addconst_out [21]}), .I2 ({new_AGEMA_signal_1133, \LED_128_Instance/addconst_out [22]}), .I3 ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}), .clk (CLK), .r (Fresh[22]), .O ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[5].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1135, \LED_128_Instance/addconst_out [20]}), .I1 ({new_AGEMA_signal_1134, \LED_128_Instance/addconst_out [21]}), .I2 ({new_AGEMA_signal_1133, \LED_128_Instance/addconst_out [22]}), .I3 ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}), .clk (CLK), .r (Fresh[23]), .O ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[6].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}), .I1 ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}), .I2 ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}), .I3 ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}), .clk (CLK), .r (Fresh[24]), .O ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[6].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}), .I1 ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}), .I2 ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}), .I3 ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}), .clk (CLK), .r (Fresh[25]), .O ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[6].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}), .I1 ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}), .I2 ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}), .I3 ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}), .clk (CLK), .r (Fresh[26]), .O ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[6].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}), .I1 ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}), .I2 ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}), .I3 ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}), .clk (CLK), .r (Fresh[27]), .O ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[7].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}), .I1 ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}), .I2 ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}), .I3 ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}), .clk (CLK), .r (Fresh[28]), .O ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[7].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}), .I1 ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}), .I2 ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}), .I3 ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}), .clk (CLK), .r (Fresh[29]), .O ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[7].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}), .I1 ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}), .I2 ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}), .I3 ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}), .clk (CLK), .r (Fresh[30]), .O ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[7].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}), .I1 ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}), .I2 ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}), .I3 ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}), .clk (CLK), .r (Fresh[31]), .O ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[8].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}), .I1 ({new_AGEMA_signal_1119, \LED_128_Instance/addconst_out [33]}), .I2 ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}), .I3 ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}), .clk (CLK), .r (Fresh[32]), .O ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[8].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}), .I1 ({new_AGEMA_signal_1119, \LED_128_Instance/addconst_out [33]}), .I2 ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}), .I3 ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}), .clk (CLK), .r (Fresh[33]), .O ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[8].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}), .I1 ({new_AGEMA_signal_1119, \LED_128_Instance/addconst_out [33]}), .I2 ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}), .I3 ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}), .clk (CLK), .r (Fresh[34]), .O ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[8].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}), .I1 ({new_AGEMA_signal_1119, \LED_128_Instance/addconst_out [33]}), .I2 ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}), .I3 ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}), .clk (CLK), .r (Fresh[35]), .O ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[9].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1124, \LED_128_Instance/addconst_out [36]}), .I1 ({new_AGEMA_signal_1123, \LED_128_Instance/addconst_out [37]}), .I2 ({new_AGEMA_signal_1122, \LED_128_Instance/addconst_out [38]}), .I3 ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}), .clk (CLK), .r (Fresh[36]), .O ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[9].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1124, \LED_128_Instance/addconst_out [36]}), .I1 ({new_AGEMA_signal_1123, \LED_128_Instance/addconst_out [37]}), .I2 ({new_AGEMA_signal_1122, \LED_128_Instance/addconst_out [38]}), .I3 ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}), .clk (CLK), .r (Fresh[37]), .O ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[9].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1124, \LED_128_Instance/addconst_out [36]}), .I1 ({new_AGEMA_signal_1123, \LED_128_Instance/addconst_out [37]}), .I2 ({new_AGEMA_signal_1122, \LED_128_Instance/addconst_out [38]}), .I3 ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}), .clk (CLK), .r (Fresh[38]), .O ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[9].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1124, \LED_128_Instance/addconst_out [36]}), .I1 ({new_AGEMA_signal_1123, \LED_128_Instance/addconst_out [37]}), .I2 ({new_AGEMA_signal_1122, \LED_128_Instance/addconst_out [38]}), .I3 ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}), .clk (CLK), .r (Fresh[39]), .O ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[10].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}), .I1 ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}), .I2 ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}), .I3 ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}), .clk (CLK), .r (Fresh[40]), .O ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[10].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}), .I1 ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}), .I2 ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}), .I3 ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}), .clk (CLK), .r (Fresh[41]), .O ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[10].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}), .I1 ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}), .I2 ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}), .I3 ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}), .clk (CLK), .r (Fresh[42]), .O ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[10].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}), .I1 ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}), .I2 ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}), .I3 ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}), .clk (CLK), .r (Fresh[43]), .O ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[11].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}), .I1 ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}), .I2 ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}), .I3 ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}), .clk (CLK), .r (Fresh[44]), .O ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[11].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}), .I1 ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}), .I2 ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}), .I3 ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}), .clk (CLK), .r (Fresh[45]), .O ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[11].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}), .I1 ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}), .I2 ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}), .I3 ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}), .clk (CLK), .r (Fresh[46]), .O ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[11].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}), .I1 ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}), .I2 ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}), .I3 ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}), .clk (CLK), .r (Fresh[47]), .O ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[12].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1129, \LED_128_Instance/addconst_out [48]}), .I1 ({new_AGEMA_signal_1128, \LED_128_Instance/addconst_out [49]}), .I2 ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}), .I3 ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}), .clk (CLK), .r (Fresh[48]), .O ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[12].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1129, \LED_128_Instance/addconst_out [48]}), .I1 ({new_AGEMA_signal_1128, \LED_128_Instance/addconst_out [49]}), .I2 ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}), .I3 ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}), .clk (CLK), .r (Fresh[49]), .O ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[12].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1129, \LED_128_Instance/addconst_out [48]}), .I1 ({new_AGEMA_signal_1128, \LED_128_Instance/addconst_out [49]}), .I2 ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}), .I3 ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}), .clk (CLK), .r (Fresh[50]), .O ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[12].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1129, \LED_128_Instance/addconst_out [48]}), .I1 ({new_AGEMA_signal_1128, \LED_128_Instance/addconst_out [49]}), .I2 ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}), .I3 ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}), .clk (CLK), .r (Fresh[51]), .O ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[13].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1132, \LED_128_Instance/addconst_out [52]}), .I1 ({new_AGEMA_signal_1131, \LED_128_Instance/addconst_out [53]}), .I2 ({new_AGEMA_signal_1130, \LED_128_Instance/addconst_out [54]}), .I3 ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}), .clk (CLK), .r (Fresh[52]), .O ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[13].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1132, \LED_128_Instance/addconst_out [52]}), .I1 ({new_AGEMA_signal_1131, \LED_128_Instance/addconst_out [53]}), .I2 ({new_AGEMA_signal_1130, \LED_128_Instance/addconst_out [54]}), .I3 ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}), .clk (CLK), .r (Fresh[53]), .O ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[13].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1132, \LED_128_Instance/addconst_out [52]}), .I1 ({new_AGEMA_signal_1131, \LED_128_Instance/addconst_out [53]}), .I2 ({new_AGEMA_signal_1130, \LED_128_Instance/addconst_out [54]}), .I3 ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}), .clk (CLK), .r (Fresh[54]), .O ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[13].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1132, \LED_128_Instance/addconst_out [52]}), .I1 ({new_AGEMA_signal_1131, \LED_128_Instance/addconst_out [53]}), .I2 ({new_AGEMA_signal_1130, \LED_128_Instance/addconst_out [54]}), .I3 ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}), .clk (CLK), .r (Fresh[55]), .O ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[14].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}), .I1 ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}), .I2 ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}), .I3 ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}), .clk (CLK), .r (Fresh[56]), .O ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[14].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}), .I1 ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}), .I2 ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}), .I3 ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}), .clk (CLK), .r (Fresh[57]), .O ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[14].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}), .I1 ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}), .I2 ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}), .I3 ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}), .clk (CLK), .r (Fresh[58]), .O ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[14].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}), .I1 ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}), .I2 ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}), .I3 ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}), .clk (CLK), .r (Fresh[59]), .O ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[15].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}), .I1 ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}), .I2 ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}), .I3 ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}), .clk (CLK), .r (Fresh[60]), .O ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[15].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}), .I1 ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}), .I2 ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}), .I3 ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}), .clk (CLK), .r (Fresh[61]), .O ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[15].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}), .I1 ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}), .I2 ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}), .I3 ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}), .clk (CLK), .r (Fresh[62]), .O ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[15].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}), .I1 ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}), .I2 ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}), .I3 ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}), .clk (CLK), .r (Fresh[63]), .O ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[0].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1203, \LED_128_Instance/mixcolumns_out [0]}), .I1 ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}), .I2 ({IN_plaintext_s1[0], IN_plaintext_s0[0]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1265, \LED_128_Instance/state [0]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[1].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1334, \LED_128_Instance/mixcolumns_out [1]}), .I1 ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}), .I2 ({IN_plaintext_s1[1], IN_plaintext_s0[1]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1345, \LED_128_Instance/state [1]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[2].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1200, \LED_128_Instance/mixcolumns_out [2]}), .I1 ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}), .I2 ({IN_plaintext_s1[2], IN_plaintext_s0[2]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1267, \LED_128_Instance/state [2]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[3].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1202, \LED_128_Instance/mixcolumns_out [3]}), .I1 ({new_AGEMA_signal_1081, \LED_128_Instance/addroundkey_out [3]}), .I2 ({IN_plaintext_s1[3], IN_plaintext_s0[3]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1269, \LED_128_Instance/state [3]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[4].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1207, \LED_128_Instance/mixcolumns_out [4]}), .I1 ({new_AGEMA_signal_1069, \LED_128_Instance/addroundkey_out [4]}), .I2 ({IN_plaintext_s1[4], IN_plaintext_s0[4]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1271, \LED_128_Instance/state [4]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[5].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1336, \LED_128_Instance/mixcolumns_out [5]}), .I1 ({new_AGEMA_signal_1053, \LED_128_Instance/addroundkey_out [5]}), .I2 ({IN_plaintext_s1[5], IN_plaintext_s0[5]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1347, \LED_128_Instance/state [5]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[6].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1204, \LED_128_Instance/mixcolumns_out [6]}), .I1 ({new_AGEMA_signal_1049, \LED_128_Instance/addroundkey_out [6]}), .I2 ({IN_plaintext_s1[6], IN_plaintext_s0[6]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1273, \LED_128_Instance/state [6]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[7].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1206, \LED_128_Instance/mixcolumns_out [7]}), .I1 ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}), .I2 ({IN_plaintext_s1[7], IN_plaintext_s0[7]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1275, \LED_128_Instance/state [7]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[8].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1210, \LED_128_Instance/mixcolumns_out [8]}), .I1 ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}), .I2 ({IN_plaintext_s1[8], IN_plaintext_s0[8]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1277, \LED_128_Instance/state [8]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[9].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1338, \LED_128_Instance/mixcolumns_out [9]}), .I1 ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}), .I2 ({IN_plaintext_s1[9], IN_plaintext_s0[9]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1349, \LED_128_Instance/state [9]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[10].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1209, \LED_128_Instance/mixcolumns_out [10]}), .I1 ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}), .I2 ({IN_plaintext_s1[10], IN_plaintext_s0[10]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1279, \LED_128_Instance/state [10]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[11].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1211, \LED_128_Instance/mixcolumns_out [11]}), .I1 ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}), .I2 ({IN_plaintext_s1[11], IN_plaintext_s0[11]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1281, \LED_128_Instance/state [11]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[12].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1215, \LED_128_Instance/mixcolumns_out [12]}), .I1 ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}), .I2 ({IN_plaintext_s1[12], IN_plaintext_s0[12]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1283, \LED_128_Instance/state [12]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[13].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1332, \LED_128_Instance/mixcolumns_out [13]}), .I1 ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}), .I2 ({IN_plaintext_s1[13], IN_plaintext_s0[13]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1351, \LED_128_Instance/state [13]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[14].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1213, \LED_128_Instance/mixcolumns_out [14]}), .I1 ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}), .I2 ({IN_plaintext_s1[14], IN_plaintext_s0[14]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1285, \LED_128_Instance/state [14]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[15].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1214, \LED_128_Instance/mixcolumns_out [15]}), .I1 ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}), .I2 ({IN_plaintext_s1[15], IN_plaintext_s0[15]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1287, \LED_128_Instance/state [15]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[16].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1297, \LED_128_Instance/mixcolumns_out [16]}), .I1 ({new_AGEMA_signal_1117, \LED_128_Instance/addroundkey_out [16]}), .I2 ({IN_plaintext_s1[16], IN_plaintext_s0[16]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1353, \LED_128_Instance/state [16]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[17].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1304, \LED_128_Instance/mixcolumns_out [17]}), .I1 ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}), .I2 ({IN_plaintext_s1[17], IN_plaintext_s0[17]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1355, \LED_128_Instance/state [17]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[18].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1340, \LED_128_Instance/mixcolumns_out [18]}), .I1 ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}), .I2 ({IN_plaintext_s1[18], IN_plaintext_s0[18]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1357, \LED_128_Instance/state [18]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[19].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1296, \LED_128_Instance/mixcolumns_out [19]}), .I1 ({new_AGEMA_signal_1113, \LED_128_Instance/addroundkey_out [19]}), .I2 ({IN_plaintext_s1[19], IN_plaintext_s0[19]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1359, \LED_128_Instance/state [19]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[20].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1306, \LED_128_Instance/mixcolumns_out [20]}), .I1 ({new_AGEMA_signal_1109, \LED_128_Instance/addroundkey_out [20]}), .I2 ({IN_plaintext_s1[20], IN_plaintext_s0[20]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1361, \LED_128_Instance/state [20]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[21].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1313, \LED_128_Instance/mixcolumns_out [21]}), .I1 ({new_AGEMA_signal_1105, \LED_128_Instance/addroundkey_out [21]}), .I2 ({IN_plaintext_s1[21], IN_plaintext_s0[21]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1363, \LED_128_Instance/state [21]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[22].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1341, \LED_128_Instance/mixcolumns_out [22]}), .I1 ({new_AGEMA_signal_1101, \LED_128_Instance/addroundkey_out [22]}), .I2 ({IN_plaintext_s1[22], IN_plaintext_s0[22]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1365, \LED_128_Instance/state [22]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[23].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1305, \LED_128_Instance/mixcolumns_out [23]}), .I1 ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}), .I2 ({IN_plaintext_s1[23], IN_plaintext_s0[23]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1367, \LED_128_Instance/state [23]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[24].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1314, \LED_128_Instance/mixcolumns_out [24]}), .I1 ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}), .I2 ({IN_plaintext_s1[24], IN_plaintext_s0[24]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1369, \LED_128_Instance/state [24]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[25].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1322, \LED_128_Instance/mixcolumns_out [25]}), .I1 ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}), .I2 ({IN_plaintext_s1[25], IN_plaintext_s0[25]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1371, \LED_128_Instance/state [25]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[26].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1342, \LED_128_Instance/mixcolumns_out [26]}), .I1 ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}), .I2 ({IN_plaintext_s1[26], IN_plaintext_s0[26]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1373, \LED_128_Instance/state [26]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[27].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1315, \LED_128_Instance/mixcolumns_out [27]}), .I1 ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}), .I2 ({IN_plaintext_s1[27], IN_plaintext_s0[27]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1375, \LED_128_Instance/state [27]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[28].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1323, \LED_128_Instance/mixcolumns_out [28]}), .I1 ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}), .I2 ({IN_plaintext_s1[28], IN_plaintext_s0[28]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1377, \LED_128_Instance/state [28]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[29].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1331, \LED_128_Instance/mixcolumns_out [29]}), .I1 ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}), .I2 ({IN_plaintext_s1[29], IN_plaintext_s0[29]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1379, \LED_128_Instance/state [29]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[30].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1343, \LED_128_Instance/mixcolumns_out [30]}), .I1 ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}), .I2 ({IN_plaintext_s1[30], IN_plaintext_s0[30]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1381, \LED_128_Instance/state [30]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[31].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1324, \LED_128_Instance/mixcolumns_out [31]}), .I1 ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}), .I2 ({IN_plaintext_s1[31], IN_plaintext_s0[31]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1383, \LED_128_Instance/state [31]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[32].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1303, \LED_128_Instance/mixcolumns_out [32]}), .I1 ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}), .I2 ({IN_plaintext_s1[32], IN_plaintext_s0[32]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1385, \LED_128_Instance/state [32]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[33].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1299, \LED_128_Instance/mixcolumns_out [33]}), .I1 ({new_AGEMA_signal_1097, \LED_128_Instance/addroundkey_out [33]}), .I2 ({IN_plaintext_s1[33], IN_plaintext_s0[33]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1387, \LED_128_Instance/state [33]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[34].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1302, \LED_128_Instance/mixcolumns_out [34]}), .I1 ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}), .I2 ({IN_plaintext_s1[34], IN_plaintext_s0[34]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1389, \LED_128_Instance/state [34]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[35].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1298, \LED_128_Instance/mixcolumns_out [35]}), .I1 ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}), .I2 ({IN_plaintext_s1[35], IN_plaintext_s0[35]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1391, \LED_128_Instance/state [35]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[36].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1312, \LED_128_Instance/mixcolumns_out [36]}), .I1 ({new_AGEMA_signal_1093, \LED_128_Instance/addroundkey_out [36]}), .I2 ({IN_plaintext_s1[36], IN_plaintext_s0[36]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1393, \LED_128_Instance/state [36]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[37].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1308, \LED_128_Instance/mixcolumns_out [37]}), .I1 ({new_AGEMA_signal_1089, \LED_128_Instance/addroundkey_out [37]}), .I2 ({IN_plaintext_s1[37], IN_plaintext_s0[37]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1395, \LED_128_Instance/state [37]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[38].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1311, \LED_128_Instance/mixcolumns_out [38]}), .I1 ({new_AGEMA_signal_1085, \LED_128_Instance/addroundkey_out [38]}), .I2 ({IN_plaintext_s1[38], IN_plaintext_s0[38]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1397, \LED_128_Instance/state [38]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[39].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1307, \LED_128_Instance/mixcolumns_out [39]}), .I1 ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}), .I2 ({IN_plaintext_s1[39], IN_plaintext_s0[39]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1399, \LED_128_Instance/state [39]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[40].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1321, \LED_128_Instance/mixcolumns_out [40]}), .I1 ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}), .I2 ({IN_plaintext_s1[40], IN_plaintext_s0[40]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1401, \LED_128_Instance/state [40]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[41].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1317, \LED_128_Instance/mixcolumns_out [41]}), .I1 ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}), .I2 ({IN_plaintext_s1[41], IN_plaintext_s0[41]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1403, \LED_128_Instance/state [41]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[42].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1320, \LED_128_Instance/mixcolumns_out [42]}), .I1 ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}), .I2 ({IN_plaintext_s1[42], IN_plaintext_s0[42]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1405, \LED_128_Instance/state [42]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[43].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1316, \LED_128_Instance/mixcolumns_out [43]}), .I1 ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}), .I2 ({IN_plaintext_s1[43], IN_plaintext_s0[43]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1407, \LED_128_Instance/state [43]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[44].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1330, \LED_128_Instance/mixcolumns_out [44]}), .I1 ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}), .I2 ({IN_plaintext_s1[44], IN_plaintext_s0[44]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1409, \LED_128_Instance/state [44]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[45].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1326, \LED_128_Instance/mixcolumns_out [45]}), .I1 ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}), .I2 ({IN_plaintext_s1[45], IN_plaintext_s0[45]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1411, \LED_128_Instance/state [45]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[46].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1329, \LED_128_Instance/mixcolumns_out [46]}), .I1 ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}), .I2 ({IN_plaintext_s1[46], IN_plaintext_s0[46]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1413, \LED_128_Instance/state [46]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[47].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1325, \LED_128_Instance/mixcolumns_out [47]}), .I1 ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}), .I2 ({IN_plaintext_s1[47], IN_plaintext_s0[47]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1415, \LED_128_Instance/state [47]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[48].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1301, \LED_128_Instance/mixcolumns_out [48]}), .I1 ({new_AGEMA_signal_1077, \LED_128_Instance/addroundkey_out [48]}), .I2 ({IN_plaintext_s1[48], IN_plaintext_s0[48]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1417, \LED_128_Instance/state [48]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[49].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1300, \LED_128_Instance/mixcolumns_out [49]}), .I1 ({new_AGEMA_signal_1073, \LED_128_Instance/addroundkey_out [49]}), .I2 ({IN_plaintext_s1[49], IN_plaintext_s0[49]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1419, \LED_128_Instance/state [49]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[50].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1201, \LED_128_Instance/mixcolumns_out [50]}), .I1 ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}), .I2 ({IN_plaintext_s1[50], IN_plaintext_s0[50]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1289, \LED_128_Instance/state [50]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[51].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1335, \LED_128_Instance/mixcolumns_out [51]}), .I1 ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}), .I2 ({IN_plaintext_s1[51], IN_plaintext_s0[51]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1421, \LED_128_Instance/state [51]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[52].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1310, \LED_128_Instance/mixcolumns_out [52]}), .I1 ({new_AGEMA_signal_1065, \LED_128_Instance/addroundkey_out [52]}), .I2 ({IN_plaintext_s1[52], IN_plaintext_s0[52]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1423, \LED_128_Instance/state [52]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[53].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1309, \LED_128_Instance/mixcolumns_out [53]}), .I1 ({new_AGEMA_signal_1061, \LED_128_Instance/addroundkey_out [53]}), .I2 ({IN_plaintext_s1[53], IN_plaintext_s0[53]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1425, \LED_128_Instance/state [53]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[54].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1205, \LED_128_Instance/mixcolumns_out [54]}), .I1 ({new_AGEMA_signal_1057, \LED_128_Instance/addroundkey_out [54]}), .I2 ({IN_plaintext_s1[54], IN_plaintext_s0[54]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1291, \LED_128_Instance/state [54]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[55].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1337, \LED_128_Instance/mixcolumns_out [55]}), .I1 ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}), .I2 ({IN_plaintext_s1[55], IN_plaintext_s0[55]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1427, \LED_128_Instance/state [55]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[56].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1319, \LED_128_Instance/mixcolumns_out [56]}), .I1 ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}), .I2 ({IN_plaintext_s1[56], IN_plaintext_s0[56]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1429, \LED_128_Instance/state [56]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[57].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1318, \LED_128_Instance/mixcolumns_out [57]}), .I1 ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}), .I2 ({IN_plaintext_s1[57], IN_plaintext_s0[57]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1431, \LED_128_Instance/state [57]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[58].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1208, \LED_128_Instance/mixcolumns_out [58]}), .I1 ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}), .I2 ({IN_plaintext_s1[58], IN_plaintext_s0[58]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1293, \LED_128_Instance/state [58]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[59].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1339, \LED_128_Instance/mixcolumns_out [59]}), .I1 ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}), .I2 ({IN_plaintext_s1[59], IN_plaintext_s0[59]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1433, \LED_128_Instance/state [59]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[60].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1328, \LED_128_Instance/mixcolumns_out [60]}), .I1 ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}), .I2 ({IN_plaintext_s1[60], IN_plaintext_s0[60]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1435, \LED_128_Instance/state [60]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[61].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1327, \LED_128_Instance/mixcolumns_out [61]}), .I1 ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}), .I2 ({IN_plaintext_s1[61], IN_plaintext_s0[61]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1437, \LED_128_Instance/state [61]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[62].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1212, \LED_128_Instance/mixcolumns_out [62]}), .I1 ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}), .I2 ({IN_plaintext_s1[62], IN_plaintext_s0[62]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1295, \LED_128_Instance/state [62]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[63].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1333, \LED_128_Instance/mixcolumns_out [63]}), .I1 ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}), .I2 ({IN_plaintext_s1[63], IN_plaintext_s0[63]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1439, \LED_128_Instance/state [63]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<2>1 ( .I0 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .I1 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I2 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I3 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I4 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .O ({new_AGEMA_signal_1200, \LED_128_Instance/mixcolumns_out [2]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<50>1 ( .I0 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I1 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .I2 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I3 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I4 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .I5 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .O ({new_AGEMA_signal_1201, \LED_128_Instance/mixcolumns_out [50]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<3>1 ( .I0 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I1 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I2 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I3 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .O ({new_AGEMA_signal_1202, \LED_128_Instance/mixcolumns_out [3]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<0>1 ( .I0 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I1 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I2 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I3 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .O ({new_AGEMA_signal_1203, \LED_128_Instance/mixcolumns_out [0]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<6>1 ( .I0 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I1 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I2 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I3 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I4 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .O ({new_AGEMA_signal_1204, \LED_128_Instance/mixcolumns_out [6]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<54>1 ( .I0 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I1 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I2 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I3 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I4 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I5 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .O ({new_AGEMA_signal_1205, \LED_128_Instance/mixcolumns_out [54]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<7>1 ( .I0 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I1 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I2 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I3 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .O ({new_AGEMA_signal_1206, \LED_128_Instance/mixcolumns_out [7]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<4>1 ( .I0 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I1 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .I2 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I3 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .O ({new_AGEMA_signal_1207, \LED_128_Instance/mixcolumns_out [4]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<58>1 ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I2 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .I3 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I4 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I5 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .O ({new_AGEMA_signal_1208, \LED_128_Instance/mixcolumns_out [58]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<10>1 ( .I0 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I1 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I2 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I3 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I4 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .O ({new_AGEMA_signal_1209, \LED_128_Instance/mixcolumns_out [10]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<8>1 ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I2 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I3 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .O ({new_AGEMA_signal_1210, \LED_128_Instance/mixcolumns_out [8]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<11>1 ( .I0 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I1 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I2 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I3 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .O ({new_AGEMA_signal_1211, \LED_128_Instance/mixcolumns_out [11]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<62>1 ( .I0 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I1 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .I2 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I3 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I4 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I5 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .O ({new_AGEMA_signal_1212, \LED_128_Instance/mixcolumns_out [62]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<14>1 ( .I0 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .I1 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I2 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I3 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I4 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1213, \LED_128_Instance/mixcolumns_out [14]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<15>1 ( .I0 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I1 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I2 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I3 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .O ({new_AGEMA_signal_1214, \LED_128_Instance/mixcolumns_out [15]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<12>1 ( .I0 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I1 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I2 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I3 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .O ({new_AGEMA_signal_1215, \LED_128_Instance/mixcolumns_out [12]}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<19>_SW0 ( .I0 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .I1 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I2 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .O ({new_AGEMA_signal_1216, N2}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<19> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I2 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I3 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .I4 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I5 ({new_AGEMA_signal_1216, N2}), .O ({new_AGEMA_signal_1296, \LED_128_Instance/mixcolumns_out [19]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<16>_SW0 ( .I0 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I1 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1217, N4}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<16> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I2 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .I3 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I4 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I5 ({new_AGEMA_signal_1217, N4}), .O ({new_AGEMA_signal_1297, \LED_128_Instance/mixcolumns_out [16]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<35>_SW0 ( .I0 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .I1 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I2 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I3 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I4 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1218, N6}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<35> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I2 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I3 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I4 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I5 ({new_AGEMA_signal_1218, N6}), .O ({new_AGEMA_signal_1298, \LED_128_Instance/mixcolumns_out [35]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<33>_SW0 ( .I0 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I1 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I2 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I3 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I4 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1219, N8}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<33> ( .I0 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I1 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I2 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I3 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I4 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .I5 ({new_AGEMA_signal_1219, N8}), .O ({new_AGEMA_signal_1299, \LED_128_Instance/mixcolumns_out [33]}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<49>_SW0 ( .I0 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I1 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I2 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1220, N12}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<49> ( .I0 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I1 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I2 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I3 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .I4 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I5 ({new_AGEMA_signal_1220, N12}), .O ({new_AGEMA_signal_1300, \LED_128_Instance/mixcolumns_out [49]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<48>_SW0 ( .I0 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .I1 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .I2 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I3 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .O ({new_AGEMA_signal_1221, N14}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<48> ( .I0 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I1 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I2 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I3 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I4 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I5 ({new_AGEMA_signal_1221, N14}), .O ({new_AGEMA_signal_1301, \LED_128_Instance/mixcolumns_out [48]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<34>_SW0 ( .I0 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I1 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I2 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I3 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .O ({new_AGEMA_signal_1222, N16}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<34> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I2 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I3 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I4 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .I5 ({new_AGEMA_signal_1222, N16}), .O ({new_AGEMA_signal_1302, \LED_128_Instance/mixcolumns_out [34]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<32>_SW0 ( .I0 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .I1 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I2 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I3 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I4 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .O ({new_AGEMA_signal_1223, N18}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<32> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I2 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I3 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I4 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .I5 ({new_AGEMA_signal_1223, N18}), .O ({new_AGEMA_signal_1303, \LED_128_Instance/mixcolumns_out [32]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<17>_SW0 ( .I0 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I1 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I2 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I3 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .O ({new_AGEMA_signal_1224, N20}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<17> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I2 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I3 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .I4 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I5 ({new_AGEMA_signal_1224, N20}), .O ({new_AGEMA_signal_1304, \LED_128_Instance/mixcolumns_out [17]}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<23>_SW0 ( .I0 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I1 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I2 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1225, N22}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<23> ( .I0 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .I1 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I2 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I3 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I4 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I5 ({new_AGEMA_signal_1225, N22}), .O ({new_AGEMA_signal_1305, \LED_128_Instance/mixcolumns_out [23]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<20>_SW0 ( .I0 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I1 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .O ({new_AGEMA_signal_1226, N24}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<20> ( .I0 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .I1 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I2 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I3 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I4 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I5 ({new_AGEMA_signal_1226, N24}), .O ({new_AGEMA_signal_1306, \LED_128_Instance/mixcolumns_out [20]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<39>_SW0 ( .I0 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I1 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I2 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I3 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I4 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1227, N26}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<39> ( .I0 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .I1 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I2 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I3 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I4 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I5 ({new_AGEMA_signal_1227, N26}), .O ({new_AGEMA_signal_1307, \LED_128_Instance/mixcolumns_out [39]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<37>_SW0 ( .I0 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I1 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I2 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I3 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I4 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1228, N28}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<37> ( .I0 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .I1 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I2 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I3 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I4 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I5 ({new_AGEMA_signal_1228, N28}), .O ({new_AGEMA_signal_1308, \LED_128_Instance/mixcolumns_out [37]}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<53>_SW0 ( .I0 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I1 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I2 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .O ({new_AGEMA_signal_1229, N32}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<53> ( .I0 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .I1 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I2 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I3 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I4 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I5 ({new_AGEMA_signal_1229, N32}), .O ({new_AGEMA_signal_1309, \LED_128_Instance/mixcolumns_out [53]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<52>_SW0 ( .I0 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I1 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I2 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I3 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1230, N34}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<52> ( .I0 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I1 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I2 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I3 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I4 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I5 ({new_AGEMA_signal_1230, N34}), .O ({new_AGEMA_signal_1310, \LED_128_Instance/mixcolumns_out [52]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<38>_SW0 ( .I0 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I1 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I2 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I3 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1231, N36}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<38> ( .I0 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .I1 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I2 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I3 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I4 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I5 ({new_AGEMA_signal_1231, N36}), .O ({new_AGEMA_signal_1311, \LED_128_Instance/mixcolumns_out [38]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<36>_SW0 ( .I0 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I1 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I2 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I3 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I4 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1232, N38}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<36> ( .I0 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .I1 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .I2 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I3 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I4 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I5 ({new_AGEMA_signal_1232, N38}), .O ({new_AGEMA_signal_1312, \LED_128_Instance/mixcolumns_out [36]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<21>_SW0 ( .I0 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I1 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I2 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I3 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1233, N40}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<21> ( .I0 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .I1 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I2 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I3 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I4 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I5 ({new_AGEMA_signal_1233, N40}), .O ({new_AGEMA_signal_1313, \LED_128_Instance/mixcolumns_out [21]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<24>_SW0 ( .I0 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I1 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .O ({new_AGEMA_signal_1234, N42}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<24> ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I2 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I3 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I4 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .I5 ({new_AGEMA_signal_1234, N42}), .O ({new_AGEMA_signal_1314, \LED_128_Instance/mixcolumns_out [24]}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<27>_SW0 ( .I0 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I1 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I2 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .O ({new_AGEMA_signal_1235, N44}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<27> ( .I0 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I1 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I2 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I3 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I4 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .I5 ({new_AGEMA_signal_1235, N44}), .O ({new_AGEMA_signal_1315, \LED_128_Instance/mixcolumns_out [27]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<43>_SW0 ( .I0 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I1 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I2 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .I3 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I4 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .O ({new_AGEMA_signal_1236, N46}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<43> ( .I0 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I1 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I2 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I3 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I4 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .I5 ({new_AGEMA_signal_1236, N46}), .O ({new_AGEMA_signal_1316, \LED_128_Instance/mixcolumns_out [43]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<41>_SW0 ( .I0 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .I1 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I2 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I3 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .I4 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .O ({new_AGEMA_signal_1237, N48}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<41> ( .I0 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I1 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I2 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I3 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I4 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I5 ({new_AGEMA_signal_1237, N48}), .O ({new_AGEMA_signal_1317, \LED_128_Instance/mixcolumns_out [41]}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<57>_SW0 ( .I0 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I1 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I2 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .O ({new_AGEMA_signal_1238, N52}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<57> ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I2 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I3 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I4 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .I5 ({new_AGEMA_signal_1238, N52}), .O ({new_AGEMA_signal_1318, \LED_128_Instance/mixcolumns_out [57]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<56>_SW0 ( .I0 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I1 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I2 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I3 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .O ({new_AGEMA_signal_1239, N54}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<56> ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I2 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I3 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I4 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I5 ({new_AGEMA_signal_1239, N54}), .O ({new_AGEMA_signal_1319, \LED_128_Instance/mixcolumns_out [56]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<42>_SW0 ( .I0 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I1 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I2 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I3 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .O ({new_AGEMA_signal_1240, N56}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<42> ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I2 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I3 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I4 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .I5 ({new_AGEMA_signal_1240, N56}), .O ({new_AGEMA_signal_1320, \LED_128_Instance/mixcolumns_out [42]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<40>_SW0 ( .I0 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .I1 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I2 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I3 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I4 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .O ({new_AGEMA_signal_1241, N58}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<40> ( .I0 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I1 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I2 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I3 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I4 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .I5 ({new_AGEMA_signal_1241, N58}), .O ({new_AGEMA_signal_1321, \LED_128_Instance/mixcolumns_out [40]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<25>_SW0 ( .I0 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .I1 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I2 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .I3 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .O ({new_AGEMA_signal_1242, N60}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<25> ( .I0 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I1 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I2 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I3 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I4 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I5 ({new_AGEMA_signal_1242, N60}), .O ({new_AGEMA_signal_1322, \LED_128_Instance/mixcolumns_out [25]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<28>_SW0 ( .I0 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I1 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .O ({new_AGEMA_signal_1243, N62}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<28> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I2 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I3 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I4 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I5 ({new_AGEMA_signal_1243, N62}), .O ({new_AGEMA_signal_1323, \LED_128_Instance/mixcolumns_out [28]}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<31>_SW0 ( .I0 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I1 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .I2 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1244, N64}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<31> ( .I0 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I1 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I2 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I3 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I4 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I5 ({new_AGEMA_signal_1244, N64}), .O ({new_AGEMA_signal_1324, \LED_128_Instance/mixcolumns_out [31]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<47>_SW0 ( .I0 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I1 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I2 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I3 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .I4 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1245, N66}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<47> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I2 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I3 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I4 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I5 ({new_AGEMA_signal_1245, N66}), .O ({new_AGEMA_signal_1325, \LED_128_Instance/mixcolumns_out [47]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<45>_SW0 ( .I0 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I1 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I2 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I3 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .I4 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1246, N68}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<45> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I2 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I3 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I4 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I5 ({new_AGEMA_signal_1246, N68}), .O ({new_AGEMA_signal_1326, \LED_128_Instance/mixcolumns_out [45]}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<61>_SW0 ( .I0 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I1 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I2 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1247, N72}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<61> ( .I0 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I1 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I2 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I3 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I4 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I5 ({new_AGEMA_signal_1247, N72}), .O ({new_AGEMA_signal_1327, \LED_128_Instance/mixcolumns_out [61]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<60>_SW0 ( .I0 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I1 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I2 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I3 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .O ({new_AGEMA_signal_1248, N74}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<60> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I2 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I3 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I4 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I5 ({new_AGEMA_signal_1248, N74}), .O ({new_AGEMA_signal_1328, \LED_128_Instance/mixcolumns_out [60]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<46>_SW0 ( .I0 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I1 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I2 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I3 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .O ({new_AGEMA_signal_1249, N76}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<46> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I2 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I3 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I4 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I5 ({new_AGEMA_signal_1249, N76}), .O ({new_AGEMA_signal_1329, \LED_128_Instance/mixcolumns_out [46]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<44>_SW0 ( .I0 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I1 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I2 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .I3 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .I4 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1250, N78}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<44> ( .I0 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I1 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I2 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I3 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I4 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I5 ({new_AGEMA_signal_1250, N78}), .O ({new_AGEMA_signal_1330, \LED_128_Instance/mixcolumns_out [44]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<29>_SW0 ( .I0 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I1 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I2 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .I3 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .O ({new_AGEMA_signal_1251, N80}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<29> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I2 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I3 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I4 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I5 ({new_AGEMA_signal_1251, N80}), .O ({new_AGEMA_signal_1331, \LED_128_Instance/mixcolumns_out [29]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<13>31_SW0 ( .I0 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I1 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .O ({new_AGEMA_signal_1252, N82}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<13>1 ( .I0 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I1 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I2 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I3 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I4 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I5 ({new_AGEMA_signal_1252, N82}), .O ({new_AGEMA_signal_1332, \LED_128_Instance/mixcolumns_out [13]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<13>31_SW1 ( .I0 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I1 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .O ({new_AGEMA_signal_1253, N84}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<63>1 ( .I0 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I1 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I2 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I3 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I4 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I5 ({new_AGEMA_signal_1253, N84}), .O ({new_AGEMA_signal_1333, \LED_128_Instance/mixcolumns_out [63]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<18>41_SW0 ( .I0 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I1 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1254, N86}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<1>1 ( .I0 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I1 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I2 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I3 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I4 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I5 ({new_AGEMA_signal_1254, N86}), .O ({new_AGEMA_signal_1334, \LED_128_Instance/mixcolumns_out [1]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<18>41_SW1 ( .I0 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I1 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1255, N88}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<51>1 ( .I0 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I1 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I2 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I3 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I4 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I5 ({new_AGEMA_signal_1255, N88}), .O ({new_AGEMA_signal_1335, \LED_128_Instance/mixcolumns_out [51]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<22>41_SW0 ( .I0 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I1 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .O ({new_AGEMA_signal_1256, N90}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<5>1 ( .I0 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I1 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I2 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I3 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I4 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .I5 ({new_AGEMA_signal_1256, N90}), .O ({new_AGEMA_signal_1336, \LED_128_Instance/mixcolumns_out [5]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<22>41_SW1 ( .I0 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I1 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .O ({new_AGEMA_signal_1257, N92}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<55>1 ( .I0 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I1 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I2 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I3 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I4 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I5 ({new_AGEMA_signal_1257, N92}), .O ({new_AGEMA_signal_1337, \LED_128_Instance/mixcolumns_out [55]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<26>41_SW0 ( .I0 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I1 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .O ({new_AGEMA_signal_1258, N94}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<9>1 ( .I0 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I1 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I2 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I3 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I4 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .I5 ({new_AGEMA_signal_1258, N94}), .O ({new_AGEMA_signal_1338, \LED_128_Instance/mixcolumns_out [9]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<26>41_SW1 ( .I0 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I1 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .O ({new_AGEMA_signal_1259, N96}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<59>1 ( .I0 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I1 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I2 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I3 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I4 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I5 ({new_AGEMA_signal_1259, N96}), .O ({new_AGEMA_signal_1339, \LED_128_Instance/mixcolumns_out [59]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<18>_SW1 ( .I0 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I1 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I2 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I3 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .I4 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I5 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .O ({new_AGEMA_signal_1260, N98}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<18> ( .I0 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I1 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I2 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I3 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I4 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .I5 ({new_AGEMA_signal_1260, N98}), .O ({new_AGEMA_signal_1340, \LED_128_Instance/mixcolumns_out [18]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<22>_SW1 ( .I0 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I1 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I2 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I3 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I4 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I5 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .O ({new_AGEMA_signal_1261, N100}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<22> ( .I0 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I1 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I2 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I3 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I4 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .I5 ({new_AGEMA_signal_1261, N100}), .O ({new_AGEMA_signal_1341, \LED_128_Instance/mixcolumns_out [22]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<26>_SW1 ( .I0 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I1 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .I2 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I3 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I4 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .I5 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .O ({new_AGEMA_signal_1262, N102}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<26> ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I2 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I3 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I4 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I5 ({new_AGEMA_signal_1262, N102}), .O ({new_AGEMA_signal_1342, \LED_128_Instance/mixcolumns_out [26]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<30>_SW1 ( .I0 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I1 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .I2 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I3 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I4 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I5 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .O ({new_AGEMA_signal_1263, N104}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<30> ( .I0 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I1 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .I2 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I3 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I4 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I5 ({new_AGEMA_signal_1263, N104}), .O ({new_AGEMA_signal_1343, \LED_128_Instance/mixcolumns_out [30]}) ) ;

    /* register cells */
    FDR \LED_128_Instance/roundconstant_5 ( .D (\LED_128_Instance/roundconstant [4]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/roundconstant [5]) ) ;
    FDR \LED_128_Instance/roundconstant_4 ( .D (\LED_128_Instance/roundconstant [3]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/roundconstant [4]) ) ;
    FDR \LED_128_Instance/roundconstant_3 ( .D (\LED_128_Instance/roundconstant [2]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/roundconstant [3]) ) ;
    FDR \LED_128_Instance/roundconstant_2 ( .D (\LED_128_Instance/roundconstant [1]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/roundconstant [2]) ) ;
    FDR \LED_128_Instance/roundconstant_1 ( .D (\LED_128_Instance/roundconstant [0]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/roundconstant [1]) ) ;
    FDS \LED_128_Instance/roundconstant_0 ( .D (\LED_128_Instance/roundconstant[5]_roundconstant[4]_XOR_7_o ), .C (clk_gated), .S (IN_reset), .Q (\LED_128_Instance/roundconstant [0]) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_63 ( .D ({new_AGEMA_signal_1439, \LED_128_Instance/state [63]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_62 ( .D ({new_AGEMA_signal_1295, \LED_128_Instance/state [62]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_61 ( .D ({new_AGEMA_signal_1437, \LED_128_Instance/state [61]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_60 ( .D ({new_AGEMA_signal_1435, \LED_128_Instance/state [60]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_59 ( .D ({new_AGEMA_signal_1433, \LED_128_Instance/state [59]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_58 ( .D ({new_AGEMA_signal_1293, \LED_128_Instance/state [58]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_57 ( .D ({new_AGEMA_signal_1431, \LED_128_Instance/state [57]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_56 ( .D ({new_AGEMA_signal_1429, \LED_128_Instance/state [56]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_55 ( .D ({new_AGEMA_signal_1427, \LED_128_Instance/state [55]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_54 ( .D ({new_AGEMA_signal_1291, \LED_128_Instance/state [54]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_53 ( .D ({new_AGEMA_signal_1425, \LED_128_Instance/state [53]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_52 ( .D ({new_AGEMA_signal_1423, \LED_128_Instance/state [52]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_51 ( .D ({new_AGEMA_signal_1421, \LED_128_Instance/state [51]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_50 ( .D ({new_AGEMA_signal_1289, \LED_128_Instance/state [50]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_49 ( .D ({new_AGEMA_signal_1419, \LED_128_Instance/state [49]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_48 ( .D ({new_AGEMA_signal_1417, \LED_128_Instance/state [48]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_47 ( .D ({new_AGEMA_signal_1415, \LED_128_Instance/state [47]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_46 ( .D ({new_AGEMA_signal_1413, \LED_128_Instance/state [46]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_45 ( .D ({new_AGEMA_signal_1411, \LED_128_Instance/state [45]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_44 ( .D ({new_AGEMA_signal_1409, \LED_128_Instance/state [44]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_43 ( .D ({new_AGEMA_signal_1407, \LED_128_Instance/state [43]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_42 ( .D ({new_AGEMA_signal_1405, \LED_128_Instance/state [42]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_41 ( .D ({new_AGEMA_signal_1403, \LED_128_Instance/state [41]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_40 ( .D ({new_AGEMA_signal_1401, \LED_128_Instance/state [40]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_39 ( .D ({new_AGEMA_signal_1399, \LED_128_Instance/state [39]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_38 ( .D ({new_AGEMA_signal_1397, \LED_128_Instance/state [38]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_37 ( .D ({new_AGEMA_signal_1395, \LED_128_Instance/state [37]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_36 ( .D ({new_AGEMA_signal_1393, \LED_128_Instance/state [36]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_35 ( .D ({new_AGEMA_signal_1391, \LED_128_Instance/state [35]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_34 ( .D ({new_AGEMA_signal_1389, \LED_128_Instance/state [34]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_33 ( .D ({new_AGEMA_signal_1387, \LED_128_Instance/state [33]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_32 ( .D ({new_AGEMA_signal_1385, \LED_128_Instance/state [32]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_31 ( .D ({new_AGEMA_signal_1383, \LED_128_Instance/state [31]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_30 ( .D ({new_AGEMA_signal_1381, \LED_128_Instance/state [30]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_29 ( .D ({new_AGEMA_signal_1379, \LED_128_Instance/state [29]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_28 ( .D ({new_AGEMA_signal_1377, \LED_128_Instance/state [28]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_27 ( .D ({new_AGEMA_signal_1375, \LED_128_Instance/state [27]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_26 ( .D ({new_AGEMA_signal_1373, \LED_128_Instance/state [26]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_25 ( .D ({new_AGEMA_signal_1371, \LED_128_Instance/state [25]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_24 ( .D ({new_AGEMA_signal_1369, \LED_128_Instance/state [24]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_23 ( .D ({new_AGEMA_signal_1367, \LED_128_Instance/state [23]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_22 ( .D ({new_AGEMA_signal_1365, \LED_128_Instance/state [22]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_21 ( .D ({new_AGEMA_signal_1363, \LED_128_Instance/state [21]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_20 ( .D ({new_AGEMA_signal_1361, \LED_128_Instance/state [20]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_19 ( .D ({new_AGEMA_signal_1359, \LED_128_Instance/state [19]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_18 ( .D ({new_AGEMA_signal_1357, \LED_128_Instance/state [18]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_17 ( .D ({new_AGEMA_signal_1355, \LED_128_Instance/state [17]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_16 ( .D ({new_AGEMA_signal_1353, \LED_128_Instance/state [16]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_15 ( .D ({new_AGEMA_signal_1287, \LED_128_Instance/state [15]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_14 ( .D ({new_AGEMA_signal_1285, \LED_128_Instance/state [14]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_13 ( .D ({new_AGEMA_signal_1351, \LED_128_Instance/state [13]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_12 ( .D ({new_AGEMA_signal_1283, \LED_128_Instance/state [12]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_11 ( .D ({new_AGEMA_signal_1281, \LED_128_Instance/state [11]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_10 ( .D ({new_AGEMA_signal_1279, \LED_128_Instance/state [10]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_9 ( .D ({new_AGEMA_signal_1349, \LED_128_Instance/state [9]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_8 ( .D ({new_AGEMA_signal_1277, \LED_128_Instance/state [8]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_7 ( .D ({new_AGEMA_signal_1275, \LED_128_Instance/state [7]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_6 ( .D ({new_AGEMA_signal_1273, \LED_128_Instance/state [6]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_5 ( .D ({new_AGEMA_signal_1347, \LED_128_Instance/state [5]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_4 ( .D ({new_AGEMA_signal_1271, \LED_128_Instance/state [4]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_3 ( .D ({new_AGEMA_signal_1269, \LED_128_Instance/state [3]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_2 ( .D ({new_AGEMA_signal_1267, \LED_128_Instance/state [2]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_1 ( .D ({new_AGEMA_signal_1345, \LED_128_Instance/state [1]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \LED_128_Instance/cipherstate_0 ( .D ({new_AGEMA_signal_1265, \LED_128_Instance/state [0]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    FDR \LED_128_Instance/ks_3 ( .D (\LED_128_Instance/ks [2]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/ks [3]) ) ;
    FDR \LED_128_Instance/ks_2 ( .D (\LED_128_Instance/ks [1]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/ks [2]) ) ;
    FDR \LED_128_Instance/ks_1 ( .D (\LED_128_Instance/ks [0]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/ks [1]) ) ;
    FDR \LED_128_Instance/ks_0 ( .D (\LED_128_Instance/ks[3]_INV_6_o ), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/ks [0]) ) ;
    FDR internal_done ( .D (internal_done_glue_set_843), .C (clk_gated), .R (IN_reset), .Q (OUT_done) ) ;
endmodule
