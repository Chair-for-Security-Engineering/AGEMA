/* modified netlist. Source: module AES in file /AES_round-based/AGEMA/AES.v */
/* clock gating is added to the circuit, the latency increased 1 time(s)  */

module AES_GHPCLL_ANF_ClockGating_d1 (plaintext_s0, key_s0, clk, reset, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] key_s1 ;
    input [127:0] plaintext_s1 ;
    input [40959:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_423 ;
    wire signal_425 ;
    wire signal_427 ;
    wire signal_429 ;
    wire signal_431 ;
    wire signal_433 ;
    wire signal_435 ;
    wire signal_437 ;
    wire signal_439 ;
    wire signal_441 ;
    wire signal_443 ;
    wire signal_445 ;
    wire signal_447 ;
    wire signal_449 ;
    wire signal_451 ;
    wire signal_453 ;
    wire signal_455 ;
    wire signal_457 ;
    wire signal_459 ;
    wire signal_461 ;
    wire signal_463 ;
    wire signal_465 ;
    wire signal_467 ;
    wire signal_469 ;
    wire signal_471 ;
    wire signal_473 ;
    wire signal_475 ;
    wire signal_477 ;
    wire signal_479 ;
    wire signal_481 ;
    wire signal_483 ;
    wire signal_485 ;
    wire signal_487 ;
    wire signal_489 ;
    wire signal_491 ;
    wire signal_493 ;
    wire signal_495 ;
    wire signal_497 ;
    wire signal_499 ;
    wire signal_501 ;
    wire signal_503 ;
    wire signal_505 ;
    wire signal_507 ;
    wire signal_509 ;
    wire signal_511 ;
    wire signal_513 ;
    wire signal_515 ;
    wire signal_517 ;
    wire signal_519 ;
    wire signal_521 ;
    wire signal_523 ;
    wire signal_525 ;
    wire signal_527 ;
    wire signal_529 ;
    wire signal_531 ;
    wire signal_533 ;
    wire signal_535 ;
    wire signal_537 ;
    wire signal_539 ;
    wire signal_541 ;
    wire signal_543 ;
    wire signal_545 ;
    wire signal_547 ;
    wire signal_549 ;
    wire signal_551 ;
    wire signal_553 ;
    wire signal_555 ;
    wire signal_557 ;
    wire signal_559 ;
    wire signal_561 ;
    wire signal_563 ;
    wire signal_565 ;
    wire signal_567 ;
    wire signal_569 ;
    wire signal_571 ;
    wire signal_573 ;
    wire signal_575 ;
    wire signal_577 ;
    wire signal_579 ;
    wire signal_581 ;
    wire signal_583 ;
    wire signal_585 ;
    wire signal_587 ;
    wire signal_589 ;
    wire signal_591 ;
    wire signal_593 ;
    wire signal_595 ;
    wire signal_597 ;
    wire signal_599 ;
    wire signal_601 ;
    wire signal_603 ;
    wire signal_605 ;
    wire signal_607 ;
    wire signal_609 ;
    wire signal_611 ;
    wire signal_613 ;
    wire signal_615 ;
    wire signal_617 ;
    wire signal_619 ;
    wire signal_621 ;
    wire signal_623 ;
    wire signal_625 ;
    wire signal_627 ;
    wire signal_629 ;
    wire signal_631 ;
    wire signal_633 ;
    wire signal_635 ;
    wire signal_637 ;
    wire signal_639 ;
    wire signal_641 ;
    wire signal_643 ;
    wire signal_645 ;
    wire signal_647 ;
    wire signal_649 ;
    wire signal_651 ;
    wire signal_653 ;
    wire signal_655 ;
    wire signal_657 ;
    wire signal_659 ;
    wire signal_661 ;
    wire signal_663 ;
    wire signal_665 ;
    wire signal_667 ;
    wire signal_669 ;
    wire signal_671 ;
    wire signal_673 ;
    wire signal_675 ;
    wire signal_792 ;
    wire signal_912 ;
    wire signal_1032 ;
    wire signal_1152 ;
    wire signal_1272 ;
    wire signal_1392 ;
    wire signal_1512 ;
    wire signal_1632 ;
    wire signal_1752 ;
    wire signal_1872 ;
    wire signal_1992 ;
    wire signal_2112 ;
    wire signal_2232 ;
    wire signal_2352 ;
    wire signal_2472 ;
    wire signal_2592 ;
    wire signal_2597 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2855 ;
    wire signal_2857 ;
    wire signal_2859 ;
    wire signal_2861 ;
    wire signal_2863 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2877 ;
    wire signal_2879 ;
    wire signal_2881 ;
    wire signal_2883 ;
    wire signal_2885 ;
    wire signal_2887 ;
    wire signal_2889 ;
    wire signal_2891 ;
    wire signal_2893 ;
    wire signal_2895 ;
    wire signal_2897 ;
    wire signal_2899 ;
    wire signal_2901 ;
    wire signal_2903 ;
    wire signal_2905 ;
    wire signal_2907 ;
    wire signal_2909 ;
    wire signal_2911 ;
    wire signal_2913 ;
    wire signal_2915 ;
    wire signal_2917 ;
    wire signal_2919 ;
    wire signal_2921 ;
    wire signal_2923 ;
    wire signal_2925 ;
    wire signal_2927 ;
    wire signal_2929 ;
    wire signal_2931 ;
    wire signal_2933 ;
    wire signal_2935 ;
    wire signal_2937 ;
    wire signal_2939 ;
    wire signal_2941 ;
    wire signal_2943 ;
    wire signal_2945 ;
    wire signal_2947 ;
    wire signal_2949 ;
    wire signal_2951 ;
    wire signal_2953 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2959 ;
    wire signal_2961 ;
    wire signal_2963 ;
    wire signal_2965 ;
    wire signal_2967 ;
    wire signal_2969 ;
    wire signal_2971 ;
    wire signal_2973 ;
    wire signal_2975 ;
    wire signal_2977 ;
    wire signal_2979 ;
    wire signal_2981 ;
    wire signal_2983 ;
    wire signal_2985 ;
    wire signal_2987 ;
    wire signal_2989 ;
    wire signal_2991 ;
    wire signal_2993 ;
    wire signal_2995 ;
    wire signal_2997 ;
    wire signal_2999 ;
    wire signal_3001 ;
    wire signal_3003 ;
    wire signal_3005 ;
    wire signal_3007 ;
    wire signal_3009 ;
    wire signal_3011 ;
    wire signal_3013 ;
    wire signal_3015 ;
    wire signal_3017 ;
    wire signal_3019 ;
    wire signal_3021 ;
    wire signal_3023 ;
    wire signal_3025 ;
    wire signal_3027 ;
    wire signal_3029 ;
    wire signal_3031 ;
    wire signal_3033 ;
    wire signal_3035 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3043 ;
    wire signal_3045 ;
    wire signal_3047 ;
    wire signal_3049 ;
    wire signal_3051 ;
    wire signal_3053 ;
    wire signal_3055 ;
    wire signal_3057 ;
    wire signal_3059 ;
    wire signal_3061 ;
    wire signal_3063 ;
    wire signal_3065 ;
    wire signal_3067 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3079 ;
    wire signal_3081 ;
    wire signal_3083 ;
    wire signal_3085 ;
    wire signal_3087 ;
    wire signal_3089 ;
    wire signal_3091 ;
    wire signal_3093 ;
    wire signal_3095 ;
    wire signal_3097 ;
    wire signal_3099 ;
    wire signal_3101 ;
    wire signal_3103 ;
    wire signal_3105 ;
    wire signal_3107 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3874 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3882 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3890 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3898 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3906 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3914 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3922 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3930 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3938 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3946 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3954 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3962 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3970 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3978 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3986 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4394 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4402 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4410 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4418 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4426 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4434 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4442 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4450 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4458 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4466 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4474 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4482 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4490 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4498 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4506 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4514 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5401 ;
    wire signal_5403 ;
    wire signal_5405 ;
    wire signal_5407 ;
    wire signal_5409 ;
    wire signal_5411 ;
    wire signal_5413 ;
    wire signal_5415 ;
    wire signal_5417 ;
    wire signal_5419 ;
    wire signal_5421 ;
    wire signal_5423 ;
    wire signal_5425 ;
    wire signal_5427 ;
    wire signal_5429 ;
    wire signal_5431 ;
    wire signal_5433 ;
    wire signal_5435 ;
    wire signal_5437 ;
    wire signal_5439 ;
    wire signal_5441 ;
    wire signal_5443 ;
    wire signal_5445 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5478 ;
    wire signal_5480 ;
    wire signal_5482 ;
    wire signal_5484 ;
    wire signal_5486 ;
    wire signal_5488 ;
    wire signal_5490 ;
    wire signal_5492 ;
    wire signal_5494 ;
    wire signal_5496 ;
    wire signal_5498 ;
    wire signal_5500 ;
    wire signal_5502 ;
    wire signal_5504 ;
    wire signal_5506 ;
    wire signal_5508 ;
    wire signal_5510 ;
    wire signal_5512 ;
    wire signal_5514 ;
    wire signal_5516 ;
    wire signal_5518 ;
    wire signal_5520 ;
    wire signal_5522 ;
    wire signal_5524 ;
    wire signal_5526 ;
    wire signal_5528 ;
    wire signal_5530 ;
    wire signal_5532 ;
    wire signal_5534 ;
    wire signal_5536 ;
    wire signal_5538 ;
    wire signal_5540 ;
    wire signal_5542 ;
    wire signal_5544 ;
    wire signal_5546 ;
    wire signal_5548 ;
    wire signal_5550 ;
    wire signal_5552 ;
    wire signal_5554 ;
    wire signal_5556 ;
    wire signal_5558 ;
    wire signal_5560 ;
    wire signal_5562 ;
    wire signal_5564 ;
    wire signal_5566 ;
    wire signal_5568 ;
    wire signal_5570 ;
    wire signal_5572 ;
    wire signal_5574 ;
    wire signal_5576 ;
    wire signal_5578 ;
    wire signal_5580 ;
    wire signal_5582 ;
    wire signal_5584 ;
    wire signal_5586 ;
    wire signal_5588 ;
    wire signal_5590 ;
    wire signal_5592 ;
    wire signal_5594 ;
    wire signal_5596 ;
    wire signal_5598 ;
    wire signal_5600 ;
    wire signal_5602 ;
    wire signal_5604 ;
    wire signal_5606 ;
    wire signal_5608 ;
    wire signal_5610 ;
    wire signal_5612 ;
    wire signal_5614 ;
    wire signal_5616 ;
    wire signal_5618 ;
    wire signal_5620 ;
    wire signal_5622 ;
    wire signal_5624 ;
    wire signal_5626 ;
    wire signal_5628 ;
    wire signal_5630 ;
    wire signal_5632 ;
    wire signal_5634 ;
    wire signal_5636 ;
    wire signal_5638 ;
    wire signal_5640 ;
    wire signal_5642 ;
    wire signal_5644 ;
    wire signal_5646 ;
    wire signal_5648 ;
    wire signal_5650 ;
    wire signal_5652 ;
    wire signal_5654 ;
    wire signal_5656 ;
    wire signal_5658 ;
    wire signal_5660 ;
    wire signal_5662 ;
    wire signal_5664 ;
    wire signal_5666 ;
    wire signal_5668 ;
    wire signal_5670 ;
    wire signal_5672 ;
    wire signal_5674 ;
    wire signal_5676 ;
    wire signal_5678 ;
    wire signal_5680 ;
    wire signal_5682 ;
    wire signal_5684 ;
    wire signal_5686 ;
    wire signal_5688 ;
    wire signal_5690 ;
    wire signal_5692 ;
    wire signal_5694 ;
    wire signal_5696 ;
    wire signal_5698 ;
    wire signal_5700 ;
    wire signal_5702 ;
    wire signal_5704 ;
    wire signal_5706 ;
    wire signal_5708 ;
    wire signal_5710 ;
    wire signal_5712 ;
    wire signal_5714 ;
    wire signal_5716 ;
    wire signal_5718 ;
    wire signal_5720 ;
    wire signal_5722 ;
    wire signal_5724 ;
    wire signal_5726 ;
    wire signal_5728 ;
    wire signal_5730 ;
    wire signal_5732 ;
    wire signal_5734 ;
    wire signal_5736 ;
    wire signal_5738 ;
    wire signal_5740 ;
    wire signal_5742 ;
    wire signal_5744 ;
    wire signal_5746 ;
    wire signal_5748 ;
    wire signal_5750 ;
    wire signal_5752 ;
    wire signal_5754 ;
    wire signal_5756 ;
    wire signal_5758 ;
    wire signal_5760 ;
    wire signal_5762 ;
    wire signal_5764 ;
    wire signal_5766 ;
    wire signal_5768 ;
    wire signal_5770 ;
    wire signal_5772 ;
    wire signal_5774 ;
    wire signal_5776 ;
    wire signal_5778 ;
    wire signal_5780 ;
    wire signal_5782 ;
    wire signal_5784 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5820 ;
    wire signal_5822 ;
    wire signal_5824 ;
    wire signal_5826 ;
    wire signal_5828 ;
    wire signal_5830 ;
    wire signal_5832 ;
    wire signal_5834 ;
    wire signal_5836 ;
    wire signal_5838 ;
    wire signal_5840 ;
    wire signal_5842 ;
    wire signal_5844 ;
    wire signal_5846 ;
    wire signal_5848 ;
    wire signal_5850 ;
    wire signal_5852 ;
    wire signal_5854 ;
    wire signal_5856 ;
    wire signal_5858 ;
    wire signal_5860 ;
    wire signal_5862 ;
    wire signal_5864 ;
    wire signal_5866 ;
    wire signal_5868 ;
    wire signal_5870 ;
    wire signal_5872 ;
    wire signal_5874 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5910 ;
    wire signal_5912 ;
    wire signal_5914 ;
    wire signal_5916 ;
    wire signal_5918 ;
    wire signal_5920 ;
    wire signal_5922 ;
    wire signal_5924 ;
    wire signal_5926 ;
    wire signal_5928 ;
    wire signal_5930 ;
    wire signal_5932 ;
    wire signal_5934 ;
    wire signal_5936 ;
    wire signal_5938 ;
    wire signal_5940 ;
    wire signal_5942 ;
    wire signal_5944 ;
    wire signal_5946 ;
    wire signal_5948 ;
    wire signal_5950 ;
    wire signal_5952 ;
    wire signal_5954 ;
    wire signal_5956 ;
    wire signal_5958 ;
    wire signal_5960 ;
    wire signal_5962 ;
    wire signal_5964 ;
    wire signal_5966 ;
    wire signal_5968 ;
    wire signal_5970 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5982 ;
    wire signal_5984 ;
    wire signal_5986 ;
    wire signal_5988 ;
    wire signal_5990 ;
    wire signal_5992 ;
    wire signal_5994 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6003 ;
    wire signal_6005 ;
    wire signal_6007 ;
    wire signal_6009 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6016 ;
    wire signal_6018 ;
    wire signal_6020 ;
    wire signal_46981 ;

    /* cells in depth 0 */
    INV_X1 cell_0 ( .A (signal_395), .ZN (signal_400) ) ;
    INV_X1 cell_1 ( .A (signal_395), .ZN (signal_401) ) ;
    INV_X1 cell_2 ( .A (signal_395), .ZN (signal_398) ) ;
    INV_X1 cell_3 ( .A (signal_395), .ZN (signal_396) ) ;
    INV_X1 cell_4 ( .A (signal_395), .ZN (signal_397) ) ;
    INV_X1 cell_5 ( .A (signal_395), .ZN (signal_399) ) ;
    NOR2_X1 cell_6 ( .A1 (signal_406), .A2 (signal_411), .ZN (signal_395) ) ;
    INV_X1 cell_7 ( .A (signal_4388), .ZN (signal_406) ) ;
    INV_X1 cell_8 ( .A (signal_395), .ZN (signal_402) ) ;
    NOR2_X1 cell_9 ( .A1 (signal_4386), .A2 (signal_4387), .ZN (signal_404) ) ;
    INV_X1 cell_10 ( .A (signal_404), .ZN (signal_403) ) ;
    NOR2_X1 cell_11 ( .A1 (signal_4388), .A2 (signal_403), .ZN (signal_4384) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_4388), .A2 (signal_4385), .ZN (signal_418) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_418), .A2 (signal_403), .ZN (signal_4383) ) ;
    NAND2_X1 cell_14 ( .A1 (signal_4385), .A2 (signal_404), .ZN (signal_411) ) ;
    INV_X1 cell_15 ( .A (signal_4386), .ZN (signal_409) ) ;
    AND2_X1 cell_16 ( .A1 (signal_409), .A2 (signal_4387), .ZN (signal_414) ) ;
    NAND2_X1 cell_17 ( .A1 (signal_418), .A2 (signal_414), .ZN (signal_405) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_402), .A2 (signal_405), .ZN (signal_4382) ) ;
    NOR2_X1 cell_19 ( .A1 (signal_4385), .A2 (signal_406), .ZN (signal_416) ) ;
    NAND2_X1 cell_20 ( .A1 (signal_414), .A2 (signal_416), .ZN (signal_408) ) ;
    NAND2_X1 cell_21 ( .A1 (signal_4385), .A2 (signal_4384), .ZN (signal_407) ) ;
    NAND2_X1 cell_22 ( .A1 (signal_408), .A2 (signal_407), .ZN (signal_4381) ) ;
    NOR2_X1 cell_23 ( .A1 (signal_4387), .A2 (signal_409), .ZN (signal_412) ) ;
    NAND2_X1 cell_24 ( .A1 (signal_418), .A2 (signal_412), .ZN (signal_410) ) ;
    NAND2_X1 cell_25 ( .A1 (signal_411), .A2 (signal_410), .ZN (signal_4380) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_416), .A2 (signal_412), .ZN (signal_413) ) ;
    NAND2_X1 cell_27 ( .A1 (signal_402), .A2 (signal_413), .ZN (signal_4379) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_156 ( .a ({signal_4549, signal_3870}), .b ({signal_4550, signal_4378}), .c ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_157 ( .a ({signal_4552, signal_3770}), .b ({signal_4553, signal_4278}), .c ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_158 ( .a ({signal_4555, signal_3769}), .b ({signal_4556, signal_4277}), .c ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_159 ( .a ({signal_4558, signal_3768}), .b ({signal_4559, signal_4276}), .c ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_160 ( .a ({signal_4561, signal_3767}), .b ({signal_4562, signal_4275}), .c ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_161 ( .a ({signal_4564, signal_3766}), .b ({signal_4565, signal_4274}), .c ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_162 ( .a ({signal_4567, signal_3765}), .b ({signal_4568, signal_4273}), .c ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_163 ( .a ({signal_4570, signal_3764}), .b ({signal_4571, signal_4272}), .c ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_164 ( .a ({signal_4573, signal_3763}), .b ({signal_4574, signal_4271}), .c ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_165 ( .a ({signal_4576, signal_3762}), .b ({signal_4577, signal_4270}), .c ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_166 ( .a ({signal_4579, signal_3761}), .b ({signal_4580, signal_4269}), .c ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_167 ( .a ({signal_4582, signal_3860}), .b ({signal_4583, signal_4368}), .c ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_168 ( .a ({signal_4585, signal_3760}), .b ({signal_4586, signal_4268}), .c ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_169 ( .a ({signal_4588, signal_3759}), .b ({signal_4589, signal_4267}), .c ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_170 ( .a ({signal_4591, signal_3758}), .b ({signal_4592, signal_4266}), .c ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_171 ( .a ({signal_4594, signal_3757}), .b ({signal_4595, signal_4265}), .c ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_172 ( .a ({signal_4597, signal_3756}), .b ({signal_4598, signal_4264}), .c ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_173 ( .a ({signal_4600, signal_3755}), .b ({signal_4601, signal_4263}), .c ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_174 ( .a ({signal_4603, signal_3754}), .b ({signal_4604, signal_4262}), .c ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_175 ( .a ({signal_4606, signal_3753}), .b ({signal_4607, signal_4261}), .c ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_176 ( .a ({signal_4609, signal_3752}), .b ({signal_4610, signal_4260}), .c ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_177 ( .a ({signal_4612, signal_3751}), .b ({signal_4613, signal_4259}), .c ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_178 ( .a ({signal_4615, signal_3859}), .b ({signal_4616, signal_4367}), .c ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_179 ( .a ({signal_4618, signal_3750}), .b ({signal_4619, signal_4258}), .c ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_180 ( .a ({signal_4621, signal_3749}), .b ({signal_4622, signal_4257}), .c ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_181 ( .a ({signal_4624, signal_3748}), .b ({signal_4625, signal_4256}), .c ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_182 ( .a ({signal_4627, signal_3747}), .b ({signal_4628, signal_4255}), .c ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_183 ( .a ({signal_4630, signal_3746}), .b ({signal_4631, signal_4254}), .c ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_184 ( .a ({signal_4633, signal_3745}), .b ({signal_4634, signal_4253}), .c ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_185 ( .a ({signal_4636, signal_3744}), .b ({signal_4637, signal_4252}), .c ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_186 ( .a ({signal_4639, signal_3743}), .b ({signal_4640, signal_4251}), .c ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_187 ( .a ({signal_4642, signal_3858}), .b ({signal_4643, signal_4366}), .c ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_188 ( .a ({signal_4645, signal_3857}), .b ({signal_4646, signal_4365}), .c ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_189 ( .a ({signal_4648, signal_3856}), .b ({signal_4649, signal_4364}), .c ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_190 ( .a ({signal_4651, signal_3855}), .b ({signal_4652, signal_4363}), .c ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_191 ( .a ({signal_4654, signal_3854}), .b ({signal_4655, signal_4362}), .c ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_192 ( .a ({signal_4657, signal_3853}), .b ({signal_4658, signal_4361}), .c ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_193 ( .a ({signal_4660, signal_3852}), .b ({signal_4661, signal_4360}), .c ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_194 ( .a ({signal_4663, signal_3851}), .b ({signal_4664, signal_4359}), .c ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_195 ( .a ({signal_4666, signal_3869}), .b ({signal_4667, signal_4377}), .c ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_196 ( .a ({signal_4669, signal_3850}), .b ({signal_4670, signal_4358}), .c ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_197 ( .a ({signal_4672, signal_3849}), .b ({signal_4673, signal_4357}), .c ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_198 ( .a ({signal_4675, signal_3848}), .b ({signal_4676, signal_4356}), .c ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_199 ( .a ({signal_4678, signal_3847}), .b ({signal_4679, signal_4355}), .c ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_200 ( .a ({signal_4681, signal_3846}), .b ({signal_4682, signal_4354}), .c ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_201 ( .a ({signal_4684, signal_3845}), .b ({signal_4685, signal_4353}), .c ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_202 ( .a ({signal_4687, signal_3844}), .b ({signal_4688, signal_4352}), .c ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_203 ( .a ({signal_4690, signal_3843}), .b ({signal_4691, signal_4351}), .c ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_204 ( .a ({signal_4693, signal_3842}), .b ({signal_4694, signal_4350}), .c ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_205 ( .a ({signal_4696, signal_3841}), .b ({signal_4697, signal_4349}), .c ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_206 ( .a ({signal_4699, signal_3868}), .b ({signal_4700, signal_4376}), .c ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_207 ( .a ({signal_4702, signal_3840}), .b ({signal_4703, signal_4348}), .c ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_208 ( .a ({signal_4705, signal_3839}), .b ({signal_4706, signal_4347}), .c ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_209 ( .a ({signal_4708, signal_3838}), .b ({signal_4709, signal_4346}), .c ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_210 ( .a ({signal_4711, signal_3837}), .b ({signal_4712, signal_4345}), .c ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_211 ( .a ({signal_4714, signal_3836}), .b ({signal_4715, signal_4344}), .c ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_212 ( .a ({signal_4717, signal_3835}), .b ({signal_4718, signal_4343}), .c ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_213 ( .a ({signal_4720, signal_3834}), .b ({signal_4721, signal_4342}), .c ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_214 ( .a ({signal_4723, signal_3833}), .b ({signal_4724, signal_4341}), .c ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_215 ( .a ({signal_4726, signal_3832}), .b ({signal_4727, signal_4340}), .c ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_216 ( .a ({signal_4729, signal_3831}), .b ({signal_4730, signal_4339}), .c ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_217 ( .a ({signal_4732, signal_3867}), .b ({signal_4733, signal_4375}), .c ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_218 ( .a ({signal_4735, signal_3830}), .b ({signal_4736, signal_4338}), .c ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_219 ( .a ({signal_4738, signal_3829}), .b ({signal_4739, signal_4337}), .c ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_220 ( .a ({signal_4741, signal_3828}), .b ({signal_4742, signal_4336}), .c ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_221 ( .a ({signal_4744, signal_3827}), .b ({signal_4745, signal_4335}), .c ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_222 ( .a ({signal_4747, signal_3826}), .b ({signal_4748, signal_4334}), .c ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_223 ( .a ({signal_4750, signal_3825}), .b ({signal_4751, signal_4333}), .c ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_224 ( .a ({signal_4753, signal_3824}), .b ({signal_4754, signal_4332}), .c ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_225 ( .a ({signal_4756, signal_3823}), .b ({signal_4757, signal_4331}), .c ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_226 ( .a ({signal_4759, signal_3822}), .b ({signal_4760, signal_4330}), .c ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_227 ( .a ({signal_4762, signal_3821}), .b ({signal_4763, signal_4329}), .c ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_228 ( .a ({signal_4765, signal_3866}), .b ({signal_4766, signal_4374}), .c ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_229 ( .a ({signal_4768, signal_3820}), .b ({signal_4769, signal_4328}), .c ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_230 ( .a ({signal_4771, signal_3819}), .b ({signal_4772, signal_4327}), .c ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_231 ( .a ({signal_4774, signal_3818}), .b ({signal_4775, signal_4326}), .c ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_232 ( .a ({signal_4777, signal_3817}), .b ({signal_4778, signal_4325}), .c ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_233 ( .a ({signal_4780, signal_3816}), .b ({signal_4781, signal_4324}), .c ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_234 ( .a ({signal_4783, signal_3815}), .b ({signal_4784, signal_4323}), .c ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_235 ( .a ({signal_4786, signal_3814}), .b ({signal_4787, signal_4322}), .c ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_236 ( .a ({signal_4789, signal_3813}), .b ({signal_4790, signal_4321}), .c ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_237 ( .a ({signal_4792, signal_3812}), .b ({signal_4793, signal_4320}), .c ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_238 ( .a ({signal_4795, signal_3811}), .b ({signal_4796, signal_4319}), .c ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_239 ( .a ({signal_4798, signal_3865}), .b ({signal_4799, signal_4373}), .c ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_240 ( .a ({signal_4801, signal_3810}), .b ({signal_4802, signal_4318}), .c ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_241 ( .a ({signal_4804, signal_3809}), .b ({signal_4805, signal_4317}), .c ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_242 ( .a ({signal_4807, signal_3808}), .b ({signal_4808, signal_4316}), .c ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_243 ( .a ({signal_4810, signal_3807}), .b ({signal_4811, signal_4315}), .c ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_244 ( .a ({signal_4813, signal_3806}), .b ({signal_4814, signal_4314}), .c ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_245 ( .a ({signal_4816, signal_3805}), .b ({signal_4817, signal_4313}), .c ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_246 ( .a ({signal_4819, signal_3804}), .b ({signal_4820, signal_4312}), .c ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_247 ( .a ({signal_4822, signal_3803}), .b ({signal_4823, signal_4311}), .c ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_248 ( .a ({signal_4825, signal_3802}), .b ({signal_4826, signal_4310}), .c ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_249 ( .a ({signal_4828, signal_3801}), .b ({signal_4829, signal_4309}), .c ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_250 ( .a ({signal_4831, signal_3864}), .b ({signal_4832, signal_4372}), .c ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_251 ( .a ({signal_4834, signal_3800}), .b ({signal_4835, signal_4308}), .c ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_252 ( .a ({signal_4837, signal_3799}), .b ({signal_4838, signal_4307}), .c ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_253 ( .a ({signal_4840, signal_3798}), .b ({signal_4841, signal_4306}), .c ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_254 ( .a ({signal_4843, signal_3797}), .b ({signal_4844, signal_4305}), .c ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_255 ( .a ({signal_4846, signal_3796}), .b ({signal_4847, signal_4304}), .c ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_256 ( .a ({signal_4849, signal_3795}), .b ({signal_4850, signal_4303}), .c ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_257 ( .a ({signal_4852, signal_3794}), .b ({signal_4853, signal_4302}), .c ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_258 ( .a ({signal_4855, signal_3793}), .b ({signal_4856, signal_4301}), .c ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_259 ( .a ({signal_4858, signal_3792}), .b ({signal_4859, signal_4300}), .c ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_260 ( .a ({signal_4861, signal_3791}), .b ({signal_4862, signal_4299}), .c ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_261 ( .a ({signal_4864, signal_3863}), .b ({signal_4865, signal_4371}), .c ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_262 ( .a ({signal_4867, signal_3790}), .b ({signal_4868, signal_4298}), .c ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_263 ( .a ({signal_4870, signal_3789}), .b ({signal_4871, signal_4297}), .c ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_264 ( .a ({signal_4873, signal_3788}), .b ({signal_4874, signal_4296}), .c ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_265 ( .a ({signal_4876, signal_3787}), .b ({signal_4877, signal_4295}), .c ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_266 ( .a ({signal_4879, signal_3786}), .b ({signal_4880, signal_4294}), .c ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_267 ( .a ({signal_4882, signal_3785}), .b ({signal_4883, signal_4293}), .c ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_268 ( .a ({signal_4885, signal_3784}), .b ({signal_4886, signal_4292}), .c ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_269 ( .a ({signal_4888, signal_3783}), .b ({signal_4889, signal_4291}), .c ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_270 ( .a ({signal_4891, signal_3782}), .b ({signal_4892, signal_4290}), .c ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_271 ( .a ({signal_4894, signal_3781}), .b ({signal_4895, signal_4289}), .c ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_272 ( .a ({signal_4897, signal_3862}), .b ({signal_4898, signal_4370}), .c ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_273 ( .a ({signal_4900, signal_3780}), .b ({signal_4901, signal_4288}), .c ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_274 ( .a ({signal_4903, signal_3779}), .b ({signal_4904, signal_4287}), .c ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_275 ( .a ({signal_4906, signal_3778}), .b ({signal_4907, signal_4286}), .c ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_276 ( .a ({signal_4909, signal_3777}), .b ({signal_4910, signal_4285}), .c ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_277 ( .a ({signal_4912, signal_3776}), .b ({signal_4913, signal_4284}), .c ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_278 ( .a ({signal_4915, signal_3775}), .b ({signal_4916, signal_4283}), .c ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_279 ( .a ({signal_4918, signal_3774}), .b ({signal_4919, signal_4282}), .c ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_280 ( .a ({signal_4921, signal_3773}), .b ({signal_4922, signal_4281}), .c ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_281 ( .a ({signal_4924, signal_3772}), .b ({signal_4925, signal_4280}), .c ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_282 ( .a ({signal_4927, signal_3771}), .b ({signal_4928, signal_4279}), .c ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_283 ( .a ({signal_4930, signal_3861}), .b ({signal_4931, signal_4369}), .c ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    NAND2_X1 cell_284 ( .A1 (signal_4385), .A2 (signal_414), .ZN (signal_415) ) ;
    NOR2_X1 cell_285 ( .A1 (signal_4388), .A2 (signal_415), .ZN (done) ) ;
    INV_X1 cell_286 ( .A (signal_416), .ZN (signal_417) ) ;
    NAND2_X1 cell_287 ( .A1 (signal_4386), .A2 (signal_4387), .ZN (signal_419) ) ;
    NOR2_X1 cell_288 ( .A1 (signal_417), .A2 (signal_419), .ZN (signal_393) ) ;
    INV_X1 cell_289 ( .A (signal_418), .ZN (signal_420) ) ;
    NOR2_X1 cell_290 ( .A1 (signal_420), .A2 (signal_419), .ZN (signal_394) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_679 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_4933, signal_792}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_807 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_4934, signal_912}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_935 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_4935, signal_1032}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_1063 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_4936, signal_1152}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_1191 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_4937, signal_1272}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_1319 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_4938, signal_1392}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_1447 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_4939, signal_1512}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_1575 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_4940, signal_1632}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_1703 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_4941, signal_1752}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_1831 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_4942, signal_1872}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_1959 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_4943, signal_1992}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_2087 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_4944, signal_2112}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_2215 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_4945, signal_2232}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_2343 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_4946, signal_2352}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_2471 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_4947, signal_2472}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_2599 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_4948, signal_2592}) ) ;
    INV_X1 cell_4187 ( .A (signal_3597), .ZN (signal_3607) ) ;
    MUX2_X1 cell_4188 ( .S (signal_3609), .A (signal_3598), .B (signal_3599), .Z (signal_3597) ) ;
    NOR2_X1 cell_4189 ( .A1 (reset), .A2 (signal_3600), .ZN (signal_3610) ) ;
    XNOR2_X1 cell_4190 ( .A (signal_4388), .B (signal_4387), .ZN (signal_3600) ) ;
    MUX2_X1 cell_4191 ( .S (signal_4385), .A (signal_3601), .B (signal_3602), .Z (signal_3608) ) ;
    NAND2_X1 cell_4192 ( .A1 (signal_3598), .A2 (signal_3603), .ZN (signal_3602) ) ;
    NAND2_X1 cell_4193 ( .A1 (signal_3609), .A2 (signal_3606), .ZN (signal_3603) ) ;
    NOR2_X1 cell_4194 ( .A1 (signal_3604), .A2 (signal_3612), .ZN (signal_3598) ) ;
    NOR2_X1 cell_4195 ( .A1 (signal_4387), .A2 (reset), .ZN (signal_3604) ) ;
    NOR2_X1 cell_4196 ( .A1 (signal_3609), .A2 (signal_3599), .ZN (signal_3601) ) ;
    NAND2_X1 cell_4197 ( .A1 (signal_4387), .A2 (signal_3605), .ZN (signal_3599) ) ;
    NOR2_X1 cell_4198 ( .A1 (reset), .A2 (signal_3611), .ZN (signal_3605) ) ;
    NOR2_X1 cell_4199 ( .A1 (reset), .A2 (signal_4388), .ZN (signal_3612) ) ;
    INV_X1 cell_4200 ( .A (reset), .ZN (signal_3606) ) ;
    INV_X1 cell_4201 ( .A (signal_4388), .ZN (signal_3611) ) ;
    INV_X1 cell_4205 ( .A (signal_4386), .ZN (signal_3609) ) ;
    ClockGatingController #(2) cell_4210 ( .clk (clk), .rst (reset), .GatedClk (signal_46981), .Synch (Synch) ) ;

    /* cells in depth 1 */
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_28 ( .s (signal_402), .b ({signal_5012, signal_3994}), .a ({signal_5244, signal_4122}), .c ({signal_5272, signal_3742}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_29 ( .s (signal_402), .b ({signal_5150, signal_4415}), .a ({signal_5039, signal_4022}), .c ({signal_5273, signal_3642}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_30 ( .s (signal_402), .b ({signal_5149, signal_4414}), .a ({signal_5038, signal_4021}), .c ({signal_5274, signal_3641}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_31 ( .s (signal_402), .b ({signal_5148, signal_4413}), .a ({signal_5037, signal_4020}), .c ({signal_5275, signal_3640}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_32 ( .s (signal_402), .b ({signal_5152, signal_4420}), .a ({signal_5036, signal_4019}), .c ({signal_5276, signal_3639}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_33 ( .s (signal_402), .b ({signal_4973, signal_3890}), .a ({signal_5035, signal_4018}), .c ({signal_5277, signal_3638}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_34 ( .s (signal_402), .b ({signal_5146, signal_4410}), .a ({signal_5237, signal_4017}), .c ({signal_5278, signal_3637}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_35 ( .s (signal_402), .b ({signal_4972, signal_3888}), .a ({signal_5034, signal_4016}), .c ({signal_5279, signal_3636}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_36 ( .s (signal_396), .b ({signal_4971, signal_3887}), .a ({signal_5033, signal_4015}), .c ({signal_5280, signal_3635}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_37 ( .s (signal_397), .b ({signal_5145, signal_4407}), .a ({signal_5032, signal_4014}), .c ({signal_5281, signal_3634}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_38 ( .s (signal_398), .b ({signal_5144, signal_4406}), .a ({signal_5031, signal_4013}), .c ({signal_5282, signal_3633}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_39 ( .s (signal_399), .b ({signal_5008, signal_3984}), .a ({signal_5124, signal_4112}), .c ({signal_5283, signal_3732}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_40 ( .s (signal_400), .b ({signal_5143, signal_4405}), .a ({signal_5030, signal_4012}), .c ({signal_5284, signal_3632}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_41 ( .s (signal_401), .b ({signal_5147, signal_4412}), .a ({signal_5029, signal_4011}), .c ({signal_5285, signal_3631}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_42 ( .s (signal_400), .b ({signal_4970, signal_3882}), .a ({signal_5028, signal_4010}), .c ({signal_5286, signal_3630}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_43 ( .s (signal_399), .b ({signal_5141, signal_4402}), .a ({signal_5027, signal_4009}), .c ({signal_5287, signal_3629}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_44 ( .s (signal_399), .b ({signal_4969, signal_3880}), .a ({signal_5026, signal_4008}), .c ({signal_5288, signal_3628}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_45 ( .s (signal_396), .b ({signal_4968, signal_3879}), .a ({signal_5025, signal_4007}), .c ({signal_5289, signal_3627}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_46 ( .s (signal_397), .b ({signal_5140, signal_4399}), .a ({signal_5024, signal_4006}), .c ({signal_5290, signal_3626}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_47 ( .s (signal_398), .b ({signal_5139, signal_4398}), .a ({signal_5023, signal_4005}), .c ({signal_5291, signal_3625}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_48 ( .s (signal_400), .b ({signal_5138, signal_4397}), .a ({signal_5022, signal_4004}), .c ({signal_5292, signal_3624}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_49 ( .s (signal_401), .b ({signal_5142, signal_4404}), .a ({signal_5021, signal_4003}), .c ({signal_5293, signal_3623}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_50 ( .s (signal_401), .b ({signal_5007, signal_3983}), .a ({signal_5123, signal_4111}), .c ({signal_5294, signal_3731}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_51 ( .s (signal_400), .b ({signal_4967, signal_3874}), .a ({signal_5020, signal_4002}), .c ({signal_5295, signal_3622}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_52 ( .s (signal_399), .b ({signal_5136, signal_4394}), .a ({signal_5019, signal_4001}), .c ({signal_5296, signal_3621}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_53 ( .s (signal_400), .b ({signal_4966, signal_3872}), .a ({signal_5018, signal_4000}), .c ({signal_5297, signal_3620}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_54 ( .s (signal_401), .b ({signal_4965, signal_3871}), .a ({signal_5017, signal_3999}), .c ({signal_5298, signal_3619}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_55 ( .s (signal_397), .b ({signal_5135, signal_4391}), .a ({signal_5016, signal_3998}), .c ({signal_5299, signal_3618}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_56 ( .s (signal_401), .b ({signal_5134, signal_4390}), .a ({signal_5015, signal_3997}), .c ({signal_5300, signal_3617}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_57 ( .s (signal_397), .b ({signal_5133, signal_4389}), .a ({signal_5014, signal_3996}), .c ({signal_5301, signal_3616}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_58 ( .s (signal_398), .b ({signal_5137, signal_4396}), .a ({signal_5013, signal_3995}), .c ({signal_5302, signal_3615}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_59 ( .s (signal_396), .b ({signal_5205, signal_4503}), .a ({signal_5122, signal_4110}), .c ({signal_5303, signal_3730}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_60 ( .s (signal_398), .b ({signal_5204, signal_4502}), .a ({signal_5121, signal_4109}), .c ({signal_5304, signal_3729}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_61 ( .s (signal_397), .b ({signal_5203, signal_4501}), .a ({signal_5120, signal_4108}), .c ({signal_5305, signal_3728}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_62 ( .s (signal_398), .b ({signal_5207, signal_4508}), .a ({signal_5119, signal_4107}), .c ({signal_5306, signal_3727}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_63 ( .s (signal_396), .b ({signal_5006, signal_3978}), .a ({signal_5118, signal_4106}), .c ({signal_5307, signal_3726}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_64 ( .s (signal_399), .b ({signal_5201, signal_4498}), .a ({signal_5117, signal_4105}), .c ({signal_5308, signal_3725}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_65 ( .s (signal_400), .b ({signal_5005, signal_3976}), .a ({signal_5116, signal_4104}), .c ({signal_5309, signal_3724}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_66 ( .s (signal_401), .b ({signal_5004, signal_3975}), .a ({signal_5115, signal_4103}), .c ({signal_5310, signal_3723}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_67 ( .s (signal_399), .b ({signal_5211, signal_4514}), .a ({signal_5132, signal_4121}), .c ({signal_5311, signal_3741}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_68 ( .s (signal_400), .b ({signal_5200, signal_4495}), .a ({signal_5114, signal_4102}), .c ({signal_5312, signal_3722}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_69 ( .s (signal_397), .b ({signal_5199, signal_4494}), .a ({signal_5113, signal_4101}), .c ({signal_5313, signal_3721}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_70 ( .s (signal_398), .b ({signal_5198, signal_4493}), .a ({signal_5112, signal_4100}), .c ({signal_5314, signal_3720}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_71 ( .s (signal_396), .b ({signal_5202, signal_4500}), .a ({signal_5111, signal_4099}), .c ({signal_5315, signal_3719}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_72 ( .s (signal_401), .b ({signal_5003, signal_3970}), .a ({signal_5110, signal_4098}), .c ({signal_5316, signal_3718}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_73 ( .s (signal_399), .b ({signal_5196, signal_4490}), .a ({signal_5109, signal_4097}), .c ({signal_5317, signal_3717}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_74 ( .s (signal_397), .b ({signal_5002, signal_3968}), .a ({signal_5108, signal_4096}), .c ({signal_5318, signal_3716}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_75 ( .s (signal_398), .b ({signal_5001, signal_3967}), .a ({signal_5107, signal_4095}), .c ({signal_5319, signal_3715}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_76 ( .s (signal_396), .b ({signal_5195, signal_4487}), .a ({signal_5106, signal_4094}), .c ({signal_5320, signal_3714}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_77 ( .s (signal_400), .b ({signal_5194, signal_4486}), .a ({signal_5105, signal_4093}), .c ({signal_5321, signal_3713}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_78 ( .s (signal_396), .b ({signal_5011, signal_3992}), .a ({signal_5131, signal_4120}), .c ({signal_5322, signal_3740}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_79 ( .s (signal_401), .b ({signal_5193, signal_4485}), .a ({signal_5104, signal_4092}), .c ({signal_5323, signal_3712}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_80 ( .s (signal_399), .b ({signal_5197, signal_4492}), .a ({signal_5103, signal_4091}), .c ({signal_5324, signal_3711}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_81 ( .s (signal_397), .b ({signal_5000, signal_3962}), .a ({signal_5242, signal_4090}), .c ({signal_5325, signal_3710}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_82 ( .s (signal_398), .b ({signal_5191, signal_4482}), .a ({signal_5102, signal_4089}), .c ({signal_5326, signal_3709}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_83 ( .s (signal_396), .b ({signal_4999, signal_3960}), .a ({signal_5101, signal_4088}), .c ({signal_5327, signal_3708}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_84 ( .s (signal_401), .b ({signal_4998, signal_3959}), .a ({signal_5100, signal_4087}), .c ({signal_5328, signal_3707}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_85 ( .s (signal_401), .b ({signal_5190, signal_4479}), .a ({signal_5099, signal_4086}), .c ({signal_5329, signal_3706}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_86 ( .s (signal_401), .b ({signal_5189, signal_4478}), .a ({signal_5098, signal_4085}), .c ({signal_5330, signal_3705}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_87 ( .s (signal_401), .b ({signal_5188, signal_4477}), .a ({signal_5097, signal_4084}), .c ({signal_5331, signal_3704}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_88 ( .s (signal_401), .b ({signal_5192, signal_4484}), .a ({signal_5096, signal_4083}), .c ({signal_5332, signal_3703}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_89 ( .s (signal_401), .b ({signal_5010, signal_3991}), .a ({signal_5130, signal_4119}), .c ({signal_5333, signal_3739}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_90 ( .s (signal_401), .b ({signal_4997, signal_3954}), .a ({signal_5095, signal_4082}), .c ({signal_5334, signal_3702}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_91 ( .s (signal_401), .b ({signal_5186, signal_4474}), .a ({signal_5241, signal_4081}), .c ({signal_5335, signal_3701}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_92 ( .s (signal_401), .b ({signal_4996, signal_3952}), .a ({signal_5094, signal_4080}), .c ({signal_5336, signal_3700}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_93 ( .s (signal_401), .b ({signal_4995, signal_3951}), .a ({signal_5093, signal_4079}), .c ({signal_5337, signal_3699}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_94 ( .s (signal_401), .b ({signal_5185, signal_4471}), .a ({signal_5092, signal_4078}), .c ({signal_5338, signal_3698}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_95 ( .s (signal_401), .b ({signal_5184, signal_4470}), .a ({signal_5091, signal_4077}), .c ({signal_5339, signal_3697}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_96 ( .s (signal_400), .b ({signal_5183, signal_4469}), .a ({signal_5090, signal_4076}), .c ({signal_5340, signal_3696}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_97 ( .s (signal_400), .b ({signal_5187, signal_4476}), .a ({signal_5089, signal_4075}), .c ({signal_5341, signal_3695}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_98 ( .s (signal_400), .b ({signal_4994, signal_3946}), .a ({signal_5088, signal_4074}), .c ({signal_5342, signal_3694}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_99 ( .s (signal_400), .b ({signal_5181, signal_4466}), .a ({signal_5087, signal_4073}), .c ({signal_5343, signal_3693}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_100 ( .s (signal_400), .b ({signal_5210, signal_4511}), .a ({signal_5129, signal_4118}), .c ({signal_5344, signal_3738}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_101 ( .s (signal_400), .b ({signal_4993, signal_3944}), .a ({signal_5086, signal_4072}), .c ({signal_5345, signal_3692}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_102 ( .s (signal_400), .b ({signal_4992, signal_3943}), .a ({signal_5085, signal_4071}), .c ({signal_5346, signal_3691}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_103 ( .s (signal_400), .b ({signal_5180, signal_4463}), .a ({signal_5084, signal_4070}), .c ({signal_5347, signal_3690}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_104 ( .s (signal_400), .b ({signal_5179, signal_4462}), .a ({signal_5083, signal_4069}), .c ({signal_5348, signal_3689}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_105 ( .s (signal_400), .b ({signal_5178, signal_4461}), .a ({signal_5082, signal_4068}), .c ({signal_5349, signal_3688}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_106 ( .s (signal_400), .b ({signal_5182, signal_4468}), .a ({signal_5081, signal_4067}), .c ({signal_5350, signal_3687}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_107 ( .s (signal_400), .b ({signal_4991, signal_3938}), .a ({signal_5080, signal_4066}), .c ({signal_5351, signal_3686}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_108 ( .s (signal_399), .b ({signal_5176, signal_4458}), .a ({signal_5079, signal_4065}), .c ({signal_5352, signal_3685}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_109 ( .s (signal_399), .b ({signal_4990, signal_3936}), .a ({signal_5078, signal_4064}), .c ({signal_5353, signal_3684}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_110 ( .s (signal_399), .b ({signal_4989, signal_3935}), .a ({signal_5077, signal_4063}), .c ({signal_5354, signal_3683}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_111 ( .s (signal_399), .b ({signal_5209, signal_4510}), .a ({signal_5128, signal_4117}), .c ({signal_5355, signal_3737}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_112 ( .s (signal_399), .b ({signal_5175, signal_4455}), .a ({signal_5076, signal_4062}), .c ({signal_5356, signal_3682}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_113 ( .s (signal_399), .b ({signal_5174, signal_4454}), .a ({signal_5075, signal_4061}), .c ({signal_5357, signal_3681}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_114 ( .s (signal_399), .b ({signal_5173, signal_4453}), .a ({signal_5074, signal_4060}), .c ({signal_5358, signal_3680}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_115 ( .s (signal_399), .b ({signal_5177, signal_4460}), .a ({signal_5073, signal_4059}), .c ({signal_5359, signal_3679}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_116 ( .s (signal_399), .b ({signal_4988, signal_3930}), .a ({signal_5240, signal_4058}), .c ({signal_5360, signal_3678}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_117 ( .s (signal_399), .b ({signal_5171, signal_4450}), .a ({signal_5072, signal_4057}), .c ({signal_5361, signal_3677}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_118 ( .s (signal_399), .b ({signal_4987, signal_3928}), .a ({signal_5071, signal_4056}), .c ({signal_5362, signal_3676}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_119 ( .s (signal_399), .b ({signal_4986, signal_3927}), .a ({signal_5070, signal_4055}), .c ({signal_5363, signal_3675}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_120 ( .s (signal_398), .b ({signal_5170, signal_4447}), .a ({signal_5069, signal_4054}), .c ({signal_5364, signal_3674}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_121 ( .s (signal_398), .b ({signal_5169, signal_4446}), .a ({signal_5068, signal_4053}), .c ({signal_5365, signal_3673}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_122 ( .s (signal_398), .b ({signal_5208, signal_4509}), .a ({signal_5127, signal_4116}), .c ({signal_5366, signal_3736}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_123 ( .s (signal_398), .b ({signal_5168, signal_4445}), .a ({signal_5067, signal_4052}), .c ({signal_5367, signal_3672}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_124 ( .s (signal_398), .b ({signal_5172, signal_4452}), .a ({signal_5066, signal_4051}), .c ({signal_5368, signal_3671}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_125 ( .s (signal_398), .b ({signal_4985, signal_3922}), .a ({signal_5065, signal_4050}), .c ({signal_5369, signal_3670}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_126 ( .s (signal_398), .b ({signal_5166, signal_4442}), .a ({signal_5239, signal_4049}), .c ({signal_5370, signal_3669}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_127 ( .s (signal_398), .b ({signal_4984, signal_3920}), .a ({signal_5064, signal_4048}), .c ({signal_5371, signal_3668}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_128 ( .s (signal_398), .b ({signal_4983, signal_3919}), .a ({signal_5063, signal_4047}), .c ({signal_5372, signal_3667}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_129 ( .s (signal_398), .b ({signal_5165, signal_4439}), .a ({signal_5062, signal_4046}), .c ({signal_5373, signal_3666}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_130 ( .s (signal_398), .b ({signal_5164, signal_4438}), .a ({signal_5061, signal_4045}), .c ({signal_5374, signal_3665}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_131 ( .s (signal_398), .b ({signal_5163, signal_4437}), .a ({signal_5060, signal_4044}), .c ({signal_5375, signal_3664}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_132 ( .s (signal_397), .b ({signal_5167, signal_4444}), .a ({signal_5059, signal_4043}), .c ({signal_5376, signal_3663}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_133 ( .s (signal_397), .b ({signal_5212, signal_4516}), .a ({signal_5126, signal_4115}), .c ({signal_5377, signal_3735}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_134 ( .s (signal_397), .b ({signal_4982, signal_3914}), .a ({signal_5058, signal_4042}), .c ({signal_5378, signal_3662}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_135 ( .s (signal_397), .b ({signal_5161, signal_4434}), .a ({signal_5057, signal_4041}), .c ({signal_5379, signal_3661}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_136 ( .s (signal_397), .b ({signal_4981, signal_3912}), .a ({signal_5056, signal_4040}), .c ({signal_5380, signal_3660}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_137 ( .s (signal_397), .b ({signal_4980, signal_3911}), .a ({signal_5055, signal_4039}), .c ({signal_5381, signal_3659}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_138 ( .s (signal_397), .b ({signal_5160, signal_4431}), .a ({signal_5054, signal_4038}), .c ({signal_5382, signal_3658}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_139 ( .s (signal_397), .b ({signal_5159, signal_4430}), .a ({signal_5053, signal_4037}), .c ({signal_5383, signal_3657}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_140 ( .s (signal_397), .b ({signal_5158, signal_4429}), .a ({signal_5052, signal_4036}), .c ({signal_5384, signal_3656}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_141 ( .s (signal_397), .b ({signal_5162, signal_4436}), .a ({signal_5051, signal_4035}), .c ({signal_5385, signal_3655}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_142 ( .s (signal_397), .b ({signal_4979, signal_3906}), .a ({signal_5050, signal_4034}), .c ({signal_5386, signal_3654}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_143 ( .s (signal_397), .b ({signal_5156, signal_4426}), .a ({signal_5049, signal_4033}), .c ({signal_5387, signal_3653}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_144 ( .s (signal_396), .b ({signal_5009, signal_3986}), .a ({signal_5125, signal_4114}), .c ({signal_5388, signal_3734}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_145 ( .s (signal_396), .b ({signal_4978, signal_3904}), .a ({signal_5048, signal_4032}), .c ({signal_5389, signal_3652}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_146 ( .s (signal_396), .b ({signal_4977, signal_3903}), .a ({signal_5047, signal_4031}), .c ({signal_5390, signal_3651}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_147 ( .s (signal_396), .b ({signal_5155, signal_4423}), .a ({signal_5046, signal_4030}), .c ({signal_5391, signal_3650}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_148 ( .s (signal_396), .b ({signal_5154, signal_4422}), .a ({signal_5045, signal_4029}), .c ({signal_5392, signal_3649}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_149 ( .s (signal_396), .b ({signal_5153, signal_4421}), .a ({signal_5044, signal_4028}), .c ({signal_5393, signal_3648}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_150 ( .s (signal_396), .b ({signal_5157, signal_4428}), .a ({signal_5043, signal_4027}), .c ({signal_5394, signal_3647}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_151 ( .s (signal_396), .b ({signal_4976, signal_3898}), .a ({signal_5238, signal_4026}), .c ({signal_5395, signal_3646}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_152 ( .s (signal_396), .b ({signal_5151, signal_4418}), .a ({signal_5042, signal_4025}), .c ({signal_5396, signal_3645}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_153 ( .s (signal_396), .b ({signal_4975, signal_3896}), .a ({signal_5041, signal_4024}), .c ({signal_5397, signal_3644}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_154 ( .s (signal_396), .b ({signal_4974, signal_3895}), .a ({signal_5040, signal_4023}), .c ({signal_5398, signal_3643}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_155 ( .s (signal_396), .b ({signal_5206, signal_4506}), .a ({signal_5243, signal_4113}), .c ({signal_5399, signal_3733}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_291 ( .s (reset), .b ({signal_5272, signal_3742}), .a ({plaintext_s1[0], plaintext_s0[0]}), .c ({signal_5478, signal_421}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_294 ( .s (reset), .b ({signal_5311, signal_3741}), .a ({plaintext_s1[1], plaintext_s0[1]}), .c ({signal_5480, signal_423}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_297 ( .s (reset), .b ({signal_5322, signal_3740}), .a ({plaintext_s1[2], plaintext_s0[2]}), .c ({signal_5482, signal_425}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_300 ( .s (reset), .b ({signal_5333, signal_3739}), .a ({plaintext_s1[3], plaintext_s0[3]}), .c ({signal_5484, signal_427}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_303 ( .s (reset), .b ({signal_5344, signal_3738}), .a ({plaintext_s1[4], plaintext_s0[4]}), .c ({signal_5486, signal_429}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_306 ( .s (reset), .b ({signal_5355, signal_3737}), .a ({plaintext_s1[5], plaintext_s0[5]}), .c ({signal_5488, signal_431}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_309 ( .s (reset), .b ({signal_5366, signal_3736}), .a ({plaintext_s1[6], plaintext_s0[6]}), .c ({signal_5490, signal_433}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_312 ( .s (reset), .b ({signal_5377, signal_3735}), .a ({plaintext_s1[7], plaintext_s0[7]}), .c ({signal_5492, signal_435}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_315 ( .s (reset), .b ({signal_5388, signal_3734}), .a ({plaintext_s1[8], plaintext_s0[8]}), .c ({signal_5494, signal_437}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_318 ( .s (reset), .b ({signal_5399, signal_3733}), .a ({plaintext_s1[9], plaintext_s0[9]}), .c ({signal_5496, signal_439}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_321 ( .s (reset), .b ({signal_5283, signal_3732}), .a ({plaintext_s1[10], plaintext_s0[10]}), .c ({signal_5498, signal_441}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_324 ( .s (reset), .b ({signal_5294, signal_3731}), .a ({plaintext_s1[11], plaintext_s0[11]}), .c ({signal_5500, signal_443}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_327 ( .s (reset), .b ({signal_5303, signal_3730}), .a ({plaintext_s1[12], plaintext_s0[12]}), .c ({signal_5502, signal_445}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_330 ( .s (reset), .b ({signal_5304, signal_3729}), .a ({plaintext_s1[13], plaintext_s0[13]}), .c ({signal_5504, signal_447}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_333 ( .s (reset), .b ({signal_5305, signal_3728}), .a ({plaintext_s1[14], plaintext_s0[14]}), .c ({signal_5506, signal_449}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_336 ( .s (reset), .b ({signal_5306, signal_3727}), .a ({plaintext_s1[15], plaintext_s0[15]}), .c ({signal_5508, signal_451}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_339 ( .s (reset), .b ({signal_5307, signal_3726}), .a ({plaintext_s1[16], plaintext_s0[16]}), .c ({signal_5510, signal_453}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_342 ( .s (reset), .b ({signal_5308, signal_3725}), .a ({plaintext_s1[17], plaintext_s0[17]}), .c ({signal_5512, signal_455}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_345 ( .s (reset), .b ({signal_5309, signal_3724}), .a ({plaintext_s1[18], plaintext_s0[18]}), .c ({signal_5514, signal_457}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_348 ( .s (reset), .b ({signal_5310, signal_3723}), .a ({plaintext_s1[19], plaintext_s0[19]}), .c ({signal_5516, signal_459}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_351 ( .s (reset), .b ({signal_5312, signal_3722}), .a ({plaintext_s1[20], plaintext_s0[20]}), .c ({signal_5518, signal_461}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_354 ( .s (reset), .b ({signal_5313, signal_3721}), .a ({plaintext_s1[21], plaintext_s0[21]}), .c ({signal_5520, signal_463}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_357 ( .s (reset), .b ({signal_5314, signal_3720}), .a ({plaintext_s1[22], plaintext_s0[22]}), .c ({signal_5522, signal_465}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_360 ( .s (reset), .b ({signal_5315, signal_3719}), .a ({plaintext_s1[23], plaintext_s0[23]}), .c ({signal_5524, signal_467}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_363 ( .s (reset), .b ({signal_5316, signal_3718}), .a ({plaintext_s1[24], plaintext_s0[24]}), .c ({signal_5526, signal_469}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_366 ( .s (reset), .b ({signal_5317, signal_3717}), .a ({plaintext_s1[25], plaintext_s0[25]}), .c ({signal_5528, signal_471}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_369 ( .s (reset), .b ({signal_5318, signal_3716}), .a ({plaintext_s1[26], plaintext_s0[26]}), .c ({signal_5530, signal_473}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_372 ( .s (reset), .b ({signal_5319, signal_3715}), .a ({plaintext_s1[27], plaintext_s0[27]}), .c ({signal_5532, signal_475}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_375 ( .s (reset), .b ({signal_5320, signal_3714}), .a ({plaintext_s1[28], plaintext_s0[28]}), .c ({signal_5534, signal_477}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_378 ( .s (reset), .b ({signal_5321, signal_3713}), .a ({plaintext_s1[29], plaintext_s0[29]}), .c ({signal_5536, signal_479}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_381 ( .s (reset), .b ({signal_5323, signal_3712}), .a ({plaintext_s1[30], plaintext_s0[30]}), .c ({signal_5538, signal_481}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_384 ( .s (reset), .b ({signal_5324, signal_3711}), .a ({plaintext_s1[31], plaintext_s0[31]}), .c ({signal_5540, signal_483}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_387 ( .s (reset), .b ({signal_5325, signal_3710}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({signal_5542, signal_485}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_390 ( .s (reset), .b ({signal_5326, signal_3709}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({signal_5544, signal_487}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_393 ( .s (reset), .b ({signal_5327, signal_3708}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({signal_5546, signal_489}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_396 ( .s (reset), .b ({signal_5328, signal_3707}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({signal_5548, signal_491}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_399 ( .s (reset), .b ({signal_5329, signal_3706}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({signal_5550, signal_493}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_402 ( .s (reset), .b ({signal_5330, signal_3705}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({signal_5552, signal_495}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_405 ( .s (reset), .b ({signal_5331, signal_3704}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({signal_5554, signal_497}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_408 ( .s (reset), .b ({signal_5332, signal_3703}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({signal_5556, signal_499}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_411 ( .s (reset), .b ({signal_5334, signal_3702}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({signal_5558, signal_501}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_414 ( .s (reset), .b ({signal_5335, signal_3701}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({signal_5560, signal_503}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_417 ( .s (reset), .b ({signal_5336, signal_3700}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({signal_5562, signal_505}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_420 ( .s (reset), .b ({signal_5337, signal_3699}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({signal_5564, signal_507}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_423 ( .s (reset), .b ({signal_5338, signal_3698}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({signal_5566, signal_509}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_426 ( .s (reset), .b ({signal_5339, signal_3697}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({signal_5568, signal_511}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_429 ( .s (reset), .b ({signal_5340, signal_3696}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({signal_5570, signal_513}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_432 ( .s (reset), .b ({signal_5341, signal_3695}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({signal_5572, signal_515}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_435 ( .s (reset), .b ({signal_5342, signal_3694}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({signal_5574, signal_517}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_438 ( .s (reset), .b ({signal_5343, signal_3693}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({signal_5576, signal_519}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_441 ( .s (reset), .b ({signal_5345, signal_3692}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({signal_5578, signal_521}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_444 ( .s (reset), .b ({signal_5346, signal_3691}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({signal_5580, signal_523}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_447 ( .s (reset), .b ({signal_5347, signal_3690}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({signal_5582, signal_525}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_450 ( .s (reset), .b ({signal_5348, signal_3689}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({signal_5584, signal_527}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_453 ( .s (reset), .b ({signal_5349, signal_3688}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({signal_5586, signal_529}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_456 ( .s (reset), .b ({signal_5350, signal_3687}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({signal_5588, signal_531}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_459 ( .s (reset), .b ({signal_5351, signal_3686}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({signal_5590, signal_533}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_462 ( .s (reset), .b ({signal_5352, signal_3685}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({signal_5592, signal_535}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_465 ( .s (reset), .b ({signal_5353, signal_3684}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({signal_5594, signal_537}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_468 ( .s (reset), .b ({signal_5354, signal_3683}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({signal_5596, signal_539}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_471 ( .s (reset), .b ({signal_5356, signal_3682}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({signal_5598, signal_541}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_474 ( .s (reset), .b ({signal_5357, signal_3681}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({signal_5600, signal_543}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_477 ( .s (reset), .b ({signal_5358, signal_3680}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({signal_5602, signal_545}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_480 ( .s (reset), .b ({signal_5359, signal_3679}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({signal_5604, signal_547}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_483 ( .s (reset), .b ({signal_5360, signal_3678}), .a ({plaintext_s1[64], plaintext_s0[64]}), .c ({signal_5606, signal_549}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_486 ( .s (reset), .b ({signal_5361, signal_3677}), .a ({plaintext_s1[65], plaintext_s0[65]}), .c ({signal_5608, signal_551}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_489 ( .s (reset), .b ({signal_5362, signal_3676}), .a ({plaintext_s1[66], plaintext_s0[66]}), .c ({signal_5610, signal_553}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_492 ( .s (reset), .b ({signal_5363, signal_3675}), .a ({plaintext_s1[67], plaintext_s0[67]}), .c ({signal_5612, signal_555}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_495 ( .s (reset), .b ({signal_5364, signal_3674}), .a ({plaintext_s1[68], plaintext_s0[68]}), .c ({signal_5614, signal_557}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_498 ( .s (reset), .b ({signal_5365, signal_3673}), .a ({plaintext_s1[69], plaintext_s0[69]}), .c ({signal_5616, signal_559}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_501 ( .s (reset), .b ({signal_5367, signal_3672}), .a ({plaintext_s1[70], plaintext_s0[70]}), .c ({signal_5618, signal_561}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_504 ( .s (reset), .b ({signal_5368, signal_3671}), .a ({plaintext_s1[71], plaintext_s0[71]}), .c ({signal_5620, signal_563}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_507 ( .s (reset), .b ({signal_5369, signal_3670}), .a ({plaintext_s1[72], plaintext_s0[72]}), .c ({signal_5622, signal_565}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_510 ( .s (reset), .b ({signal_5370, signal_3669}), .a ({plaintext_s1[73], plaintext_s0[73]}), .c ({signal_5624, signal_567}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_513 ( .s (reset), .b ({signal_5371, signal_3668}), .a ({plaintext_s1[74], plaintext_s0[74]}), .c ({signal_5626, signal_569}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_516 ( .s (reset), .b ({signal_5372, signal_3667}), .a ({plaintext_s1[75], plaintext_s0[75]}), .c ({signal_5628, signal_571}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_519 ( .s (reset), .b ({signal_5373, signal_3666}), .a ({plaintext_s1[76], plaintext_s0[76]}), .c ({signal_5630, signal_573}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_522 ( .s (reset), .b ({signal_5374, signal_3665}), .a ({plaintext_s1[77], plaintext_s0[77]}), .c ({signal_5632, signal_575}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_525 ( .s (reset), .b ({signal_5375, signal_3664}), .a ({plaintext_s1[78], plaintext_s0[78]}), .c ({signal_5634, signal_577}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_528 ( .s (reset), .b ({signal_5376, signal_3663}), .a ({plaintext_s1[79], plaintext_s0[79]}), .c ({signal_5636, signal_579}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_531 ( .s (reset), .b ({signal_5378, signal_3662}), .a ({plaintext_s1[80], plaintext_s0[80]}), .c ({signal_5638, signal_581}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_534 ( .s (reset), .b ({signal_5379, signal_3661}), .a ({plaintext_s1[81], plaintext_s0[81]}), .c ({signal_5640, signal_583}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_537 ( .s (reset), .b ({signal_5380, signal_3660}), .a ({plaintext_s1[82], plaintext_s0[82]}), .c ({signal_5642, signal_585}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_540 ( .s (reset), .b ({signal_5381, signal_3659}), .a ({plaintext_s1[83], plaintext_s0[83]}), .c ({signal_5644, signal_587}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_543 ( .s (reset), .b ({signal_5382, signal_3658}), .a ({plaintext_s1[84], plaintext_s0[84]}), .c ({signal_5646, signal_589}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_546 ( .s (reset), .b ({signal_5383, signal_3657}), .a ({plaintext_s1[85], plaintext_s0[85]}), .c ({signal_5648, signal_591}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_549 ( .s (reset), .b ({signal_5384, signal_3656}), .a ({plaintext_s1[86], plaintext_s0[86]}), .c ({signal_5650, signal_593}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_552 ( .s (reset), .b ({signal_5385, signal_3655}), .a ({plaintext_s1[87], plaintext_s0[87]}), .c ({signal_5652, signal_595}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_555 ( .s (reset), .b ({signal_5386, signal_3654}), .a ({plaintext_s1[88], plaintext_s0[88]}), .c ({signal_5654, signal_597}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_558 ( .s (reset), .b ({signal_5387, signal_3653}), .a ({plaintext_s1[89], plaintext_s0[89]}), .c ({signal_5656, signal_599}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_561 ( .s (reset), .b ({signal_5389, signal_3652}), .a ({plaintext_s1[90], plaintext_s0[90]}), .c ({signal_5658, signal_601}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_564 ( .s (reset), .b ({signal_5390, signal_3651}), .a ({plaintext_s1[91], plaintext_s0[91]}), .c ({signal_5660, signal_603}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_567 ( .s (reset), .b ({signal_5391, signal_3650}), .a ({plaintext_s1[92], plaintext_s0[92]}), .c ({signal_5662, signal_605}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_570 ( .s (reset), .b ({signal_5392, signal_3649}), .a ({plaintext_s1[93], plaintext_s0[93]}), .c ({signal_5664, signal_607}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_573 ( .s (reset), .b ({signal_5393, signal_3648}), .a ({plaintext_s1[94], plaintext_s0[94]}), .c ({signal_5666, signal_609}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_576 ( .s (reset), .b ({signal_5394, signal_3647}), .a ({plaintext_s1[95], plaintext_s0[95]}), .c ({signal_5668, signal_611}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_579 ( .s (reset), .b ({signal_5395, signal_3646}), .a ({plaintext_s1[96], plaintext_s0[96]}), .c ({signal_5670, signal_613}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_582 ( .s (reset), .b ({signal_5396, signal_3645}), .a ({plaintext_s1[97], plaintext_s0[97]}), .c ({signal_5672, signal_615}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_585 ( .s (reset), .b ({signal_5397, signal_3644}), .a ({plaintext_s1[98], plaintext_s0[98]}), .c ({signal_5674, signal_617}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_588 ( .s (reset), .b ({signal_5398, signal_3643}), .a ({plaintext_s1[99], plaintext_s0[99]}), .c ({signal_5676, signal_619}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_591 ( .s (reset), .b ({signal_5273, signal_3642}), .a ({plaintext_s1[100], plaintext_s0[100]}), .c ({signal_5678, signal_621}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_594 ( .s (reset), .b ({signal_5274, signal_3641}), .a ({plaintext_s1[101], plaintext_s0[101]}), .c ({signal_5680, signal_623}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_597 ( .s (reset), .b ({signal_5275, signal_3640}), .a ({plaintext_s1[102], plaintext_s0[102]}), .c ({signal_5682, signal_625}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_600 ( .s (reset), .b ({signal_5276, signal_3639}), .a ({plaintext_s1[103], plaintext_s0[103]}), .c ({signal_5684, signal_627}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_603 ( .s (reset), .b ({signal_5277, signal_3638}), .a ({plaintext_s1[104], plaintext_s0[104]}), .c ({signal_5686, signal_629}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_606 ( .s (reset), .b ({signal_5278, signal_3637}), .a ({plaintext_s1[105], plaintext_s0[105]}), .c ({signal_5688, signal_631}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_609 ( .s (reset), .b ({signal_5279, signal_3636}), .a ({plaintext_s1[106], plaintext_s0[106]}), .c ({signal_5690, signal_633}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_612 ( .s (reset), .b ({signal_5280, signal_3635}), .a ({plaintext_s1[107], plaintext_s0[107]}), .c ({signal_5692, signal_635}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_615 ( .s (reset), .b ({signal_5281, signal_3634}), .a ({plaintext_s1[108], plaintext_s0[108]}), .c ({signal_5694, signal_637}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_618 ( .s (reset), .b ({signal_5282, signal_3633}), .a ({plaintext_s1[109], plaintext_s0[109]}), .c ({signal_5696, signal_639}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_621 ( .s (reset), .b ({signal_5284, signal_3632}), .a ({plaintext_s1[110], plaintext_s0[110]}), .c ({signal_5698, signal_641}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_624 ( .s (reset), .b ({signal_5285, signal_3631}), .a ({plaintext_s1[111], plaintext_s0[111]}), .c ({signal_5700, signal_643}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_627 ( .s (reset), .b ({signal_5286, signal_3630}), .a ({plaintext_s1[112], plaintext_s0[112]}), .c ({signal_5702, signal_645}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_630 ( .s (reset), .b ({signal_5287, signal_3629}), .a ({plaintext_s1[113], plaintext_s0[113]}), .c ({signal_5704, signal_647}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_633 ( .s (reset), .b ({signal_5288, signal_3628}), .a ({plaintext_s1[114], plaintext_s0[114]}), .c ({signal_5706, signal_649}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_636 ( .s (reset), .b ({signal_5289, signal_3627}), .a ({plaintext_s1[115], plaintext_s0[115]}), .c ({signal_5708, signal_651}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_639 ( .s (reset), .b ({signal_5290, signal_3626}), .a ({plaintext_s1[116], plaintext_s0[116]}), .c ({signal_5710, signal_653}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_642 ( .s (reset), .b ({signal_5291, signal_3625}), .a ({plaintext_s1[117], plaintext_s0[117]}), .c ({signal_5712, signal_655}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_645 ( .s (reset), .b ({signal_5292, signal_3624}), .a ({plaintext_s1[118], plaintext_s0[118]}), .c ({signal_5714, signal_657}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_648 ( .s (reset), .b ({signal_5293, signal_3623}), .a ({plaintext_s1[119], plaintext_s0[119]}), .c ({signal_5716, signal_659}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_651 ( .s (reset), .b ({signal_5295, signal_3622}), .a ({plaintext_s1[120], plaintext_s0[120]}), .c ({signal_5718, signal_661}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_654 ( .s (reset), .b ({signal_5296, signal_3621}), .a ({plaintext_s1[121], plaintext_s0[121]}), .c ({signal_5720, signal_663}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_657 ( .s (reset), .b ({signal_5297, signal_3620}), .a ({plaintext_s1[122], plaintext_s0[122]}), .c ({signal_5722, signal_665}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_660 ( .s (reset), .b ({signal_5298, signal_3619}), .a ({plaintext_s1[123], plaintext_s0[123]}), .c ({signal_5724, signal_667}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_663 ( .s (reset), .b ({signal_5299, signal_3618}), .a ({plaintext_s1[124], plaintext_s0[124]}), .c ({signal_5726, signal_669}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_666 ( .s (reset), .b ({signal_5300, signal_3617}), .a ({plaintext_s1[125], plaintext_s0[125]}), .c ({signal_5728, signal_671}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_669 ( .s (reset), .b ({signal_5301, signal_3616}), .a ({plaintext_s1[126], plaintext_s0[126]}), .c ({signal_5730, signal_673}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_672 ( .s (reset), .b ({signal_5302, signal_3615}), .a ({plaintext_s1[127], plaintext_s0[127]}), .c ({signal_5732, signal_675}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(0)) cell_2723 ( .a ({signal_4949, signal_2597}), .b ({signal_5141, signal_4402}), .c ({signal_5237, signal_4017}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(0)) cell_2815 ( .a ({signal_4950, signal_2660}), .b ({signal_4973, signal_3890}), .c ({signal_5238, signal_4026}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(0)) cell_2831 ( .a ({signal_4951, signal_2661}), .b ({signal_5161, signal_4434}), .c ({signal_5239, signal_4049}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(0)) cell_2923 ( .a ({signal_4952, signal_2724}), .b ({signal_4985, signal_3922}), .c ({signal_5240, signal_4058}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(0)) cell_2939 ( .a ({signal_4953, signal_2725}), .b ({signal_5181, signal_4466}), .c ({signal_5241, signal_4081}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(0)) cell_3031 ( .a ({signal_4954, signal_2788}), .b ({signal_4997, signal_3954}), .c ({signal_5242, signal_4090}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(0)) cell_3047 ( .a ({signal_4955, signal_2789}), .b ({signal_5201, signal_4498}), .c ({signal_5243, signal_4113}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(0)) cell_3139 ( .a ({signal_4956, signal_2852}), .b ({signal_5009, signal_3986}), .c ({signal_5244, signal_4122}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3155 ( .s (reset), .b ({signal_5908, signal_4250}), .a ({key_s1[0], key_s0[0]}), .c ({signal_5910, signal_2853}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3158 ( .s (reset), .b ({signal_5894, signal_4249}), .a ({key_s1[1], key_s0[1]}), .c ({signal_5912, signal_2855}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3161 ( .s (reset), .b ({signal_5886, signal_4248}), .a ({key_s1[2], key_s0[2]}), .c ({signal_5914, signal_2857}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3164 ( .s (reset), .b ({signal_5883, signal_4247}), .a ({key_s1[3], key_s0[3]}), .c ({signal_5916, signal_2859}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3167 ( .s (reset), .b ({signal_5882, signal_4246}), .a ({key_s1[4], key_s0[4]}), .c ({signal_5918, signal_2861}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3170 ( .s (reset), .b ({signal_5881, signal_4245}), .a ({key_s1[5], key_s0[5]}), .c ({signal_5920, signal_2863}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3173 ( .s (reset), .b ({signal_5880, signal_4244}), .a ({key_s1[6], key_s0[6]}), .c ({signal_5922, signal_2865}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3176 ( .s (reset), .b ({signal_5879, signal_4243}), .a ({key_s1[7], key_s0[7]}), .c ({signal_5924, signal_2867}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3179 ( .s (reset), .b ({signal_5878, signal_4242}), .a ({key_s1[8], key_s0[8]}), .c ({signal_5926, signal_2869}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3182 ( .s (reset), .b ({signal_5877, signal_4241}), .a ({key_s1[9], key_s0[9]}), .c ({signal_5928, signal_2871}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3185 ( .s (reset), .b ({signal_5907, signal_4240}), .a ({key_s1[10], key_s0[10]}), .c ({signal_5930, signal_2873}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3188 ( .s (reset), .b ({signal_5906, signal_4239}), .a ({key_s1[11], key_s0[11]}), .c ({signal_5932, signal_2875}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3191 ( .s (reset), .b ({signal_5902, signal_4238}), .a ({key_s1[12], key_s0[12]}), .c ({signal_5934, signal_2877}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3194 ( .s (reset), .b ({signal_5901, signal_4237}), .a ({key_s1[13], key_s0[13]}), .c ({signal_5936, signal_2879}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3197 ( .s (reset), .b ({signal_5900, signal_4236}), .a ({key_s1[14], key_s0[14]}), .c ({signal_5938, signal_2881}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3200 ( .s (reset), .b ({signal_5899, signal_4235}), .a ({key_s1[15], key_s0[15]}), .c ({signal_5940, signal_2883}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3203 ( .s (reset), .b ({signal_5898, signal_4234}), .a ({key_s1[16], key_s0[16]}), .c ({signal_5942, signal_2885}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3206 ( .s (reset), .b ({signal_5897, signal_4233}), .a ({key_s1[17], key_s0[17]}), .c ({signal_5944, signal_2887}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3209 ( .s (reset), .b ({signal_5896, signal_4232}), .a ({key_s1[18], key_s0[18]}), .c ({signal_5946, signal_2889}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3212 ( .s (reset), .b ({signal_5895, signal_4231}), .a ({key_s1[19], key_s0[19]}), .c ({signal_5948, signal_2891}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3215 ( .s (reset), .b ({signal_5893, signal_4230}), .a ({key_s1[20], key_s0[20]}), .c ({signal_5950, signal_2893}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3218 ( .s (reset), .b ({signal_5892, signal_4229}), .a ({key_s1[21], key_s0[21]}), .c ({signal_5952, signal_2895}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3221 ( .s (reset), .b ({signal_5891, signal_4228}), .a ({key_s1[22], key_s0[22]}), .c ({signal_5954, signal_2897}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3224 ( .s (reset), .b ({signal_5890, signal_4227}), .a ({key_s1[23], key_s0[23]}), .c ({signal_5956, signal_2899}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3227 ( .s (reset), .b ({signal_5980, signal_4226}), .a ({key_s1[24], key_s0[24]}), .c ({signal_5982, signal_2901}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3230 ( .s (reset), .b ({signal_5979, signal_4225}), .a ({key_s1[25], key_s0[25]}), .c ({signal_5984, signal_2903}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3233 ( .s (reset), .b ({signal_6014, signal_4224}), .a ({key_s1[26], key_s0[26]}), .c ({signal_6016, signal_2905}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3236 ( .s (reset), .b ({signal_6013, signal_4223}), .a ({key_s1[27], key_s0[27]}), .c ({signal_6018, signal_2907}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3239 ( .s (reset), .b ({signal_5999, signal_4222}), .a ({key_s1[28], key_s0[28]}), .c ({signal_6003, signal_2909}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3242 ( .s (reset), .b ({signal_6012, signal_4221}), .a ({key_s1[29], key_s0[29]}), .c ({signal_6020, signal_2911}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3245 ( .s (reset), .b ({signal_5974, signal_4220}), .a ({key_s1[30], key_s0[30]}), .c ({signal_5986, signal_2913}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3248 ( .s (reset), .b ({signal_5997, signal_4219}), .a ({key_s1[31], key_s0[31]}), .c ({signal_6005, signal_2915}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3251 ( .s (reset), .b ({signal_5815, signal_4218}), .a ({key_s1[32], key_s0[32]}), .c ({signal_5820, signal_2917}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3254 ( .s (reset), .b ({signal_5802, signal_4217}), .a ({key_s1[33], key_s0[33]}), .c ({signal_5822, signal_2919}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3257 ( .s (reset), .b ({signal_5795, signal_4216}), .a ({key_s1[34], key_s0[34]}), .c ({signal_5824, signal_2921}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3260 ( .s (reset), .b ({signal_5793, signal_4215}), .a ({key_s1[35], key_s0[35]}), .c ({signal_5826, signal_2923}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3263 ( .s (reset), .b ({signal_5792, signal_4214}), .a ({key_s1[36], key_s0[36]}), .c ({signal_5828, signal_2925}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3266 ( .s (reset), .b ({signal_5791, signal_4213}), .a ({key_s1[37], key_s0[37]}), .c ({signal_5830, signal_2927}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3269 ( .s (reset), .b ({signal_5790, signal_4212}), .a ({key_s1[38], key_s0[38]}), .c ({signal_5832, signal_2929}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3272 ( .s (reset), .b ({signal_5789, signal_4211}), .a ({key_s1[39], key_s0[39]}), .c ({signal_5834, signal_2931}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3275 ( .s (reset), .b ({signal_5788, signal_4210}), .a ({key_s1[40], key_s0[40]}), .c ({signal_5836, signal_2933}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3278 ( .s (reset), .b ({signal_5787, signal_4209}), .a ({key_s1[41], key_s0[41]}), .c ({signal_5838, signal_2935}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3281 ( .s (reset), .b ({signal_5814, signal_4208}), .a ({key_s1[42], key_s0[42]}), .c ({signal_5840, signal_2937}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3284 ( .s (reset), .b ({signal_5813, signal_4207}), .a ({key_s1[43], key_s0[43]}), .c ({signal_5842, signal_2939}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3287 ( .s (reset), .b ({signal_5810, signal_4206}), .a ({key_s1[44], key_s0[44]}), .c ({signal_5844, signal_2941}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3290 ( .s (reset), .b ({signal_5809, signal_4205}), .a ({key_s1[45], key_s0[45]}), .c ({signal_5846, signal_2943}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3293 ( .s (reset), .b ({signal_5808, signal_4204}), .a ({key_s1[46], key_s0[46]}), .c ({signal_5848, signal_2945}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3296 ( .s (reset), .b ({signal_5807, signal_4203}), .a ({key_s1[47], key_s0[47]}), .c ({signal_5850, signal_2947}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3299 ( .s (reset), .b ({signal_5806, signal_4202}), .a ({key_s1[48], key_s0[48]}), .c ({signal_5852, signal_2949}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3302 ( .s (reset), .b ({signal_5805, signal_4201}), .a ({key_s1[49], key_s0[49]}), .c ({signal_5854, signal_2951}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3305 ( .s (reset), .b ({signal_5804, signal_4200}), .a ({key_s1[50], key_s0[50]}), .c ({signal_5856, signal_2953}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3308 ( .s (reset), .b ({signal_5803, signal_4199}), .a ({key_s1[51], key_s0[51]}), .c ({signal_5858, signal_2955}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3311 ( .s (reset), .b ({signal_5801, signal_4198}), .a ({key_s1[52], key_s0[52]}), .c ({signal_5860, signal_2957}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3314 ( .s (reset), .b ({signal_5800, signal_4197}), .a ({key_s1[53], key_s0[53]}), .c ({signal_5862, signal_2959}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3317 ( .s (reset), .b ({signal_5799, signal_4196}), .a ({key_s1[54], key_s0[54]}), .c ({signal_5864, signal_2961}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3320 ( .s (reset), .b ({signal_5798, signal_4195}), .a ({key_s1[55], key_s0[55]}), .c ({signal_5866, signal_2963}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3323 ( .s (reset), .b ({signal_5889, signal_4194}), .a ({key_s1[56], key_s0[56]}), .c ({signal_5958, signal_2965}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3326 ( .s (reset), .b ({signal_5888, signal_4193}), .a ({key_s1[57], key_s0[57]}), .c ({signal_5960, signal_2967}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3329 ( .s (reset), .b ({signal_6001, signal_4192}), .a ({key_s1[58], key_s0[58]}), .c ({signal_6007, signal_2969}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3332 ( .s (reset), .b ({signal_6000, signal_4191}), .a ({key_s1[59], key_s0[59]}), .c ({signal_6009, signal_2971}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3335 ( .s (reset), .b ({signal_5976, signal_4190}), .a ({key_s1[60], key_s0[60]}), .c ({signal_5988, signal_2973}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3338 ( .s (reset), .b ({signal_5998, signal_4189}), .a ({key_s1[61], key_s0[61]}), .c ({signal_6011, signal_2975}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3341 ( .s (reset), .b ({signal_5885, signal_4188}), .a ({key_s1[62], key_s0[62]}), .c ({signal_5962, signal_2977}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3344 ( .s (reset), .b ({signal_5973, signal_4187}), .a ({key_s1[63], key_s0[63]}), .c ({signal_5990, signal_2979}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3347 ( .s (reset), .b ({signal_5474, signal_4186}), .a ({key_s1[64], key_s0[64]}), .c ({signal_5734, signal_2981}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3350 ( .s (reset), .b ({signal_5460, signal_4185}), .a ({key_s1[65], key_s0[65]}), .c ({signal_5736, signal_2983}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3353 ( .s (reset), .b ({signal_5455, signal_4184}), .a ({key_s1[66], key_s0[66]}), .c ({signal_5738, signal_2985}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3356 ( .s (reset), .b ({signal_5454, signal_4183}), .a ({key_s1[67], key_s0[67]}), .c ({signal_5740, signal_2987}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3359 ( .s (reset), .b ({signal_5453, signal_4182}), .a ({key_s1[68], key_s0[68]}), .c ({signal_5742, signal_2989}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3362 ( .s (reset), .b ({signal_5452, signal_4181}), .a ({key_s1[69], key_s0[69]}), .c ({signal_5744, signal_2991}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3365 ( .s (reset), .b ({signal_5451, signal_4180}), .a ({key_s1[70], key_s0[70]}), .c ({signal_5746, signal_2993}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3368 ( .s (reset), .b ({signal_5450, signal_4179}), .a ({key_s1[71], key_s0[71]}), .c ({signal_5748, signal_2995}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3371 ( .s (reset), .b ({signal_5449, signal_4178}), .a ({key_s1[72], key_s0[72]}), .c ({signal_5750, signal_2997}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3374 ( .s (reset), .b ({signal_5448, signal_4177}), .a ({key_s1[73], key_s0[73]}), .c ({signal_5752, signal_2999}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3377 ( .s (reset), .b ({signal_5473, signal_4176}), .a ({key_s1[74], key_s0[74]}), .c ({signal_5754, signal_3001}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3380 ( .s (reset), .b ({signal_5472, signal_4175}), .a ({key_s1[75], key_s0[75]}), .c ({signal_5756, signal_3003}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3383 ( .s (reset), .b ({signal_5468, signal_4174}), .a ({key_s1[76], key_s0[76]}), .c ({signal_5758, signal_3005}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3386 ( .s (reset), .b ({signal_5467, signal_4173}), .a ({key_s1[77], key_s0[77]}), .c ({signal_5760, signal_3007}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3389 ( .s (reset), .b ({signal_5466, signal_4172}), .a ({key_s1[78], key_s0[78]}), .c ({signal_5762, signal_3009}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3392 ( .s (reset), .b ({signal_5465, signal_4171}), .a ({key_s1[79], key_s0[79]}), .c ({signal_5764, signal_3011}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3395 ( .s (reset), .b ({signal_5464, signal_4170}), .a ({key_s1[80], key_s0[80]}), .c ({signal_5766, signal_3013}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3398 ( .s (reset), .b ({signal_5463, signal_4169}), .a ({key_s1[81], key_s0[81]}), .c ({signal_5768, signal_3015}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3401 ( .s (reset), .b ({signal_5462, signal_4168}), .a ({key_s1[82], key_s0[82]}), .c ({signal_5770, signal_3017}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3404 ( .s (reset), .b ({signal_5461, signal_4167}), .a ({key_s1[83], key_s0[83]}), .c ({signal_5772, signal_3019}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3407 ( .s (reset), .b ({signal_5459, signal_4166}), .a ({key_s1[84], key_s0[84]}), .c ({signal_5774, signal_3021}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3410 ( .s (reset), .b ({signal_5458, signal_4165}), .a ({key_s1[85], key_s0[85]}), .c ({signal_5776, signal_3023}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3413 ( .s (reset), .b ({signal_5457, signal_4164}), .a ({key_s1[86], key_s0[86]}), .c ({signal_5778, signal_3025}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3416 ( .s (reset), .b ({signal_5456, signal_4163}), .a ({key_s1[87], key_s0[87]}), .c ({signal_5780, signal_3027}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3419 ( .s (reset), .b ({signal_5797, signal_4162}), .a ({key_s1[88], key_s0[88]}), .c ({signal_5868, signal_3029}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3422 ( .s (reset), .b ({signal_5796, signal_4161}), .a ({key_s1[89], key_s0[89]}), .c ({signal_5870, signal_3031}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3425 ( .s (reset), .b ({signal_5978, signal_4160}), .a ({key_s1[90], key_s0[90]}), .c ({signal_5992, signal_3033}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3428 ( .s (reset), .b ({signal_5977, signal_4159}), .a ({key_s1[91], key_s0[91]}), .c ({signal_5994, signal_3035}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3431 ( .s (reset), .b ({signal_5887, signal_4158}), .a ({key_s1[92], key_s0[92]}), .c ({signal_5964, signal_3037}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3434 ( .s (reset), .b ({signal_5975, signal_4157}), .a ({key_s1[93], key_s0[93]}), .c ({signal_5996, signal_3039}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3437 ( .s (reset), .b ({signal_5794, signal_4156}), .a ({key_s1[94], key_s0[94]}), .c ({signal_5872, signal_3041}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3440 ( .s (reset), .b ({signal_5884, signal_4155}), .a ({key_s1[95], key_s0[95]}), .c ({signal_5966, signal_3043}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3443 ( .s (reset), .b ({signal_5268, signal_4154}), .a ({key_s1[96], key_s0[96]}), .c ({signal_5401, signal_3045}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3446 ( .s (reset), .b ({signal_5247, signal_4153}), .a ({key_s1[97], key_s0[97]}), .c ({signal_5403, signal_3047}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3449 ( .s (reset), .b ({signal_5246, signal_4152}), .a ({key_s1[98], key_s0[98]}), .c ({signal_5405, signal_3049}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3452 ( .s (reset), .b ({signal_5245, signal_4151}), .a ({key_s1[99], key_s0[99]}), .c ({signal_5407, signal_3051}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3455 ( .s (reset), .b ({signal_5267, signal_4150}), .a ({key_s1[100], key_s0[100]}), .c ({signal_5409, signal_3053}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3458 ( .s (reset), .b ({signal_5266, signal_4149}), .a ({key_s1[101], key_s0[101]}), .c ({signal_5411, signal_3055}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3461 ( .s (reset), .b ({signal_5265, signal_4148}), .a ({key_s1[102], key_s0[102]}), .c ({signal_5413, signal_3057}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3464 ( .s (reset), .b ({signal_5264, signal_4147}), .a ({key_s1[103], key_s0[103]}), .c ({signal_5415, signal_3059}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3467 ( .s (reset), .b ({signal_5263, signal_4146}), .a ({key_s1[104], key_s0[104]}), .c ({signal_5417, signal_3061}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3470 ( .s (reset), .b ({signal_5262, signal_4145}), .a ({key_s1[105], key_s0[105]}), .c ({signal_5419, signal_3063}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3473 ( .s (reset), .b ({signal_5261, signal_4144}), .a ({key_s1[106], key_s0[106]}), .c ({signal_5421, signal_3065}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3476 ( .s (reset), .b ({signal_5260, signal_4143}), .a ({key_s1[107], key_s0[107]}), .c ({signal_5423, signal_3067}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3479 ( .s (reset), .b ({signal_5259, signal_4142}), .a ({key_s1[108], key_s0[108]}), .c ({signal_5425, signal_3069}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3482 ( .s (reset), .b ({signal_5258, signal_4141}), .a ({key_s1[109], key_s0[109]}), .c ({signal_5427, signal_3071}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3485 ( .s (reset), .b ({signal_5257, signal_4140}), .a ({key_s1[110], key_s0[110]}), .c ({signal_5429, signal_3073}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3488 ( .s (reset), .b ({signal_5256, signal_4139}), .a ({key_s1[111], key_s0[111]}), .c ({signal_5431, signal_3075}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3491 ( .s (reset), .b ({signal_5255, signal_4138}), .a ({key_s1[112], key_s0[112]}), .c ({signal_5433, signal_3077}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3494 ( .s (reset), .b ({signal_5254, signal_4137}), .a ({key_s1[113], key_s0[113]}), .c ({signal_5435, signal_3079}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3497 ( .s (reset), .b ({signal_5253, signal_4136}), .a ({key_s1[114], key_s0[114]}), .c ({signal_5437, signal_3081}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3500 ( .s (reset), .b ({signal_5252, signal_4135}), .a ({key_s1[115], key_s0[115]}), .c ({signal_5439, signal_3083}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3503 ( .s (reset), .b ({signal_5251, signal_4134}), .a ({key_s1[116], key_s0[116]}), .c ({signal_5441, signal_3085}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3506 ( .s (reset), .b ({signal_5250, signal_4133}), .a ({key_s1[117], key_s0[117]}), .c ({signal_5443, signal_3087}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3509 ( .s (reset), .b ({signal_5249, signal_4132}), .a ({key_s1[118], key_s0[118]}), .c ({signal_5445, signal_3089}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3512 ( .s (reset), .b ({signal_5248, signal_4131}), .a ({key_s1[119], key_s0[119]}), .c ({signal_5447, signal_3091}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3515 ( .s (reset), .b ({signal_5471, signal_4130}), .a ({key_s1[120], key_s0[120]}), .c ({signal_5782, signal_3093}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3518 ( .s (reset), .b ({signal_5470, signal_4129}), .a ({key_s1[121], key_s0[121]}), .c ({signal_5784, signal_3095}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3521 ( .s (reset), .b ({signal_5905, signal_4128}), .a ({key_s1[122], key_s0[122]}), .c ({signal_5968, signal_3097}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3524 ( .s (reset), .b ({signal_5904, signal_4127}), .a ({key_s1[123], key_s0[123]}), .c ({signal_5970, signal_3099}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3527 ( .s (reset), .b ({signal_5812, signal_4126}), .a ({key_s1[124], key_s0[124]}), .c ({signal_5874, signal_3101}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3530 ( .s (reset), .b ({signal_5903, signal_4125}), .a ({key_s1[125], key_s0[125]}), .c ({signal_5972, signal_3103}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3533 ( .s (reset), .b ({signal_5469, signal_4124}), .a ({key_s1[126], key_s0[126]}), .c ({signal_5786, signal_3105}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) cell_3536 ( .s (reset), .b ({signal_5811, signal_4123}), .a ({key_s1[127], key_s0[127]}), .c ({signal_5876, signal_3107}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3539 ( .a ({signal_4931, signal_4369}), .b ({signal_5787, signal_4209}), .c ({signal_5877, signal_4241}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3540 ( .a ({signal_4898, signal_4370}), .b ({signal_5788, signal_4210}), .c ({signal_5878, signal_4242}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3541 ( .a ({signal_4865, signal_4371}), .b ({signal_5789, signal_4211}), .c ({signal_5879, signal_4243}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3542 ( .a ({signal_4832, signal_4372}), .b ({signal_5790, signal_4212}), .c ({signal_5880, signal_4244}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3543 ( .a ({signal_4799, signal_4373}), .b ({signal_5791, signal_4213}), .c ({signal_5881, signal_4245}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3544 ( .a ({signal_4766, signal_4374}), .b ({signal_5792, signal_4214}), .c ({signal_5882, signal_4246}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3545 ( .a ({signal_4739, signal_4337}), .b ({signal_5448, signal_4177}), .c ({signal_5787, signal_4209}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3546 ( .a ({signal_4844, signal_4305}), .b ({signal_5262, signal_4145}), .c ({signal_5448, signal_4177}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3547 ( .a ({signal_4736, signal_4338}), .b ({signal_5449, signal_4178}), .c ({signal_5788, signal_4210}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3548 ( .a ({signal_4841, signal_4306}), .b ({signal_5263, signal_4146}), .c ({signal_5449, signal_4178}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3549 ( .a ({signal_4733, signal_4375}), .b ({signal_5793, signal_4215}), .c ({signal_5883, signal_4247}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3550 ( .a ({signal_4730, signal_4339}), .b ({signal_5450, signal_4179}), .c ({signal_5789, signal_4211}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3551 ( .a ({signal_4838, signal_4307}), .b ({signal_5264, signal_4147}), .c ({signal_5450, signal_4179}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3552 ( .a ({signal_4727, signal_4340}), .b ({signal_5451, signal_4180}), .c ({signal_5790, signal_4212}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3553 ( .a ({signal_4835, signal_4308}), .b ({signal_5265, signal_4148}), .c ({signal_5451, signal_4180}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3554 ( .a ({signal_4724, signal_4341}), .b ({signal_5452, signal_4181}), .c ({signal_5791, signal_4213}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3555 ( .a ({signal_4829, signal_4309}), .b ({signal_5266, signal_4149}), .c ({signal_5452, signal_4181}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3556 ( .a ({signal_4721, signal_4342}), .b ({signal_5453, signal_4182}), .c ({signal_5792, signal_4214}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3557 ( .a ({signal_4826, signal_4310}), .b ({signal_5267, signal_4150}), .c ({signal_5453, signal_4182}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3558 ( .a ({signal_4718, signal_4343}), .b ({signal_5454, signal_4183}), .c ({signal_5793, signal_4215}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3559 ( .a ({signal_4823, signal_4311}), .b ({signal_5245, signal_4151}), .c ({signal_5454, signal_4183}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3560 ( .a ({signal_4928, signal_4279}), .b ({signal_5233, signal_4545}), .c ({signal_5245, signal_4151}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3561 ( .a ({signal_4706, signal_4347}), .b ({signal_5973, signal_4187}), .c ({signal_5997, signal_4219}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3562 ( .a ({signal_4811, signal_4315}), .b ({signal_5884, signal_4155}), .c ({signal_5973, signal_4187}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3563 ( .a ({signal_4916, signal_4283}), .b ({signal_5811, signal_4123}), .c ({signal_5884, signal_4155}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3564 ( .a ({signal_4703, signal_4348}), .b ({signal_5885, signal_4188}), .c ({signal_5974, signal_4220}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3565 ( .a ({signal_4808, signal_4316}), .b ({signal_5794, signal_4156}), .c ({signal_5885, signal_4188}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3566 ( .a ({signal_4913, signal_4284}), .b ({signal_5469, signal_4124}), .c ({signal_5794, signal_4156}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3567 ( .a ({signal_4700, signal_4376}), .b ({signal_5795, signal_4216}), .c ({signal_5886, signal_4248}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3568 ( .a ({signal_4715, signal_4344}), .b ({signal_5455, signal_4184}), .c ({signal_5795, signal_4216}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3569 ( .a ({signal_4820, signal_4312}), .b ({signal_5246, signal_4152}), .c ({signal_5455, signal_4184}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3570 ( .a ({signal_4925, signal_4280}), .b ({signal_5234, signal_4546}), .c ({signal_5246, signal_4152}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3571 ( .a ({signal_4697, signal_4349}), .b ({signal_5998, signal_4189}), .c ({signal_6012, signal_4221}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3572 ( .a ({signal_4805, signal_4317}), .b ({signal_5975, signal_4157}), .c ({signal_5998, signal_4189}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3573 ( .a ({signal_4910, signal_4285}), .b ({signal_5903, signal_4125}), .c ({signal_5975, signal_4157}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3574 ( .a ({signal_4694, signal_4350}), .b ({signal_5976, signal_4190}), .c ({signal_5999, signal_4222}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3575 ( .a ({signal_4802, signal_4318}), .b ({signal_5887, signal_4158}), .c ({signal_5976, signal_4190}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3576 ( .a ({signal_4907, signal_4286}), .b ({signal_5812, signal_4126}), .c ({signal_5887, signal_4158}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3577 ( .a ({signal_4691, signal_4351}), .b ({signal_6000, signal_4191}), .c ({signal_6013, signal_4223}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3578 ( .a ({signal_4796, signal_4319}), .b ({signal_5977, signal_4159}), .c ({signal_6000, signal_4191}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3579 ( .a ({signal_4904, signal_4287}), .b ({signal_5904, signal_4127}), .c ({signal_5977, signal_4159}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3580 ( .a ({signal_4688, signal_4352}), .b ({signal_6001, signal_4192}), .c ({signal_6014, signal_4224}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3581 ( .a ({signal_4793, signal_4320}), .b ({signal_5978, signal_4160}), .c ({signal_6001, signal_4192}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3582 ( .a ({signal_4901, signal_4288}), .b ({signal_5905, signal_4128}), .c ({signal_5978, signal_4160}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3583 ( .a ({signal_4685, signal_4353}), .b ({signal_5888, signal_4193}), .c ({signal_5979, signal_4225}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3584 ( .a ({signal_4790, signal_4321}), .b ({signal_5796, signal_4161}), .c ({signal_5888, signal_4193}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3585 ( .a ({signal_4895, signal_4289}), .b ({signal_5470, signal_4129}), .c ({signal_5796, signal_4161}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3586 ( .a ({signal_4682, signal_4354}), .b ({signal_5889, signal_4194}), .c ({signal_5980, signal_4226}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3587 ( .a ({signal_4787, signal_4322}), .b ({signal_5797, signal_4162}), .c ({signal_5889, signal_4194}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3588 ( .a ({signal_4892, signal_4290}), .b ({signal_5471, signal_4130}), .c ({signal_5797, signal_4162}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3589 ( .a ({signal_4679, signal_4355}), .b ({signal_5798, signal_4195}), .c ({signal_5890, signal_4227}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3590 ( .a ({signal_4784, signal_4323}), .b ({signal_5456, signal_4163}), .c ({signal_5798, signal_4195}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3591 ( .a ({signal_4889, signal_4291}), .b ({signal_5248, signal_4131}), .c ({signal_5456, signal_4163}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3592 ( .a ({signal_4676, signal_4356}), .b ({signal_5799, signal_4196}), .c ({signal_5891, signal_4228}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3593 ( .a ({signal_4781, signal_4324}), .b ({signal_5457, signal_4164}), .c ({signal_5799, signal_4196}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3594 ( .a ({signal_4886, signal_4292}), .b ({signal_5249, signal_4132}), .c ({signal_5457, signal_4164}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3595 ( .a ({signal_4673, signal_4357}), .b ({signal_5800, signal_4197}), .c ({signal_5892, signal_4229}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3596 ( .a ({signal_4778, signal_4325}), .b ({signal_5458, signal_4165}), .c ({signal_5800, signal_4197}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3597 ( .a ({signal_4883, signal_4293}), .b ({signal_5250, signal_4133}), .c ({signal_5458, signal_4165}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3598 ( .a ({signal_4670, signal_4358}), .b ({signal_5801, signal_4198}), .c ({signal_5893, signal_4230}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3599 ( .a ({signal_4775, signal_4326}), .b ({signal_5459, signal_4166}), .c ({signal_5801, signal_4198}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3600 ( .a ({signal_4880, signal_4294}), .b ({signal_5251, signal_4134}), .c ({signal_5459, signal_4166}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3601 ( .a ({signal_4667, signal_4377}), .b ({signal_5802, signal_4217}), .c ({signal_5894, signal_4249}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3602 ( .a ({signal_4712, signal_4345}), .b ({signal_5460, signal_4185}), .c ({signal_5802, signal_4217}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3603 ( .a ({signal_4817, signal_4313}), .b ({signal_5247, signal_4153}), .c ({signal_5460, signal_4185}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3604 ( .a ({signal_4922, signal_4281}), .b ({signal_5235, signal_4547}), .c ({signal_5247, signal_4153}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3605 ( .a ({signal_4664, signal_4359}), .b ({signal_5803, signal_4199}), .c ({signal_5895, signal_4231}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3606 ( .a ({signal_4772, signal_4327}), .b ({signal_5461, signal_4167}), .c ({signal_5803, signal_4199}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3607 ( .a ({signal_4877, signal_4295}), .b ({signal_5252, signal_4135}), .c ({signal_5461, signal_4167}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3608 ( .a ({signal_4661, signal_4360}), .b ({signal_5804, signal_4200}), .c ({signal_5896, signal_4232}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3609 ( .a ({signal_4769, signal_4328}), .b ({signal_5462, signal_4168}), .c ({signal_5804, signal_4200}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3610 ( .a ({signal_4874, signal_4296}), .b ({signal_5253, signal_4136}), .c ({signal_5462, signal_4168}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3611 ( .a ({signal_4658, signal_4361}), .b ({signal_5805, signal_4201}), .c ({signal_5897, signal_4233}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3612 ( .a ({signal_4763, signal_4329}), .b ({signal_5463, signal_4169}), .c ({signal_5805, signal_4201}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3613 ( .a ({signal_4871, signal_4297}), .b ({signal_5254, signal_4137}), .c ({signal_5463, signal_4169}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3614 ( .a ({signal_4655, signal_4362}), .b ({signal_5806, signal_4202}), .c ({signal_5898, signal_4234}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3615 ( .a ({signal_4760, signal_4330}), .b ({signal_5464, signal_4170}), .c ({signal_5806, signal_4202}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3616 ( .a ({signal_4868, signal_4298}), .b ({signal_5255, signal_4138}), .c ({signal_5464, signal_4170}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3617 ( .a ({signal_4652, signal_4363}), .b ({signal_5807, signal_4203}), .c ({signal_5899, signal_4235}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3618 ( .a ({signal_4757, signal_4331}), .b ({signal_5465, signal_4171}), .c ({signal_5807, signal_4203}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3619 ( .a ({signal_4862, signal_4299}), .b ({signal_5256, signal_4139}), .c ({signal_5465, signal_4171}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3620 ( .a ({signal_4649, signal_4364}), .b ({signal_5808, signal_4204}), .c ({signal_5900, signal_4236}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3621 ( .a ({signal_4754, signal_4332}), .b ({signal_5466, signal_4172}), .c ({signal_5808, signal_4204}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3622 ( .a ({signal_4859, signal_4300}), .b ({signal_5257, signal_4140}), .c ({signal_5466, signal_4172}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3623 ( .a ({signal_4646, signal_4365}), .b ({signal_5809, signal_4205}), .c ({signal_5901, signal_4237}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3624 ( .a ({signal_4751, signal_4333}), .b ({signal_5467, signal_4173}), .c ({signal_5809, signal_4205}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3625 ( .a ({signal_4856, signal_4301}), .b ({signal_5258, signal_4141}), .c ({signal_5467, signal_4173}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3626 ( .a ({signal_4643, signal_4366}), .b ({signal_5810, signal_4206}), .c ({signal_5902, signal_4238}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3627 ( .a ({signal_4748, signal_4334}), .b ({signal_5468, signal_4174}), .c ({signal_5810, signal_4206}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3628 ( .a ({signal_4853, signal_4302}), .b ({signal_5259, signal_4142}), .c ({signal_5468, signal_4174}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3629 ( .a ({signal_4640, signal_4251}), .b ({signal_5475, signal_4517}), .c ({signal_5811, signal_4123}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3630 ( .a ({signal_4637, signal_4252}), .b ({signal_5269, signal_4518}), .c ({signal_5469, signal_4124}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3631 ( .a ({signal_4634, signal_4253}), .b ({signal_5816, signal_4519}), .c ({signal_5903, signal_4125}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3632 ( .a ({signal_4631, signal_4254}), .b ({signal_5476, signal_4520}), .c ({signal_5812, signal_4126}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3633 ( .a ({signal_4628, signal_4255}), .b ({signal_5817, signal_4521}), .c ({signal_5904, signal_4127}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3634 ( .a ({signal_4625, signal_4256}), .b ({signal_5818, signal_4522}), .c ({signal_5905, signal_4128}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3635 ( .a ({signal_4622, signal_4257}), .b ({signal_5270, signal_4523}), .c ({signal_5470, signal_4129}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3636 ( .a ({signal_4619, signal_4258}), .b ({signal_5271, signal_4524}), .c ({signal_5471, signal_4130}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3637 ( .a ({signal_4616, signal_4367}), .b ({signal_5813, signal_4207}), .c ({signal_5906, signal_4239}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3638 ( .a ({signal_4745, signal_4335}), .b ({signal_5472, signal_4175}), .c ({signal_5813, signal_4207}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3639 ( .a ({signal_4850, signal_4303}), .b ({signal_5260, signal_4143}), .c ({signal_5472, signal_4175}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3640 ( .a ({signal_4613, signal_4259}), .b ({signal_5213, signal_4525}), .c ({signal_5248, signal_4131}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3641 ( .a ({signal_4610, signal_4260}), .b ({signal_5214, signal_4526}), .c ({signal_5249, signal_4132}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3642 ( .a ({signal_4607, signal_4261}), .b ({signal_5215, signal_4527}), .c ({signal_5250, signal_4133}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3643 ( .a ({signal_4604, signal_4262}), .b ({signal_5216, signal_4528}), .c ({signal_5251, signal_4134}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3644 ( .a ({signal_4601, signal_4263}), .b ({signal_5217, signal_4529}), .c ({signal_5252, signal_4135}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3645 ( .a ({signal_4598, signal_4264}), .b ({signal_5218, signal_4530}), .c ({signal_5253, signal_4136}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3646 ( .a ({signal_4595, signal_4265}), .b ({signal_5219, signal_4531}), .c ({signal_5254, signal_4137}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3647 ( .a ({signal_4592, signal_4266}), .b ({signal_5220, signal_4532}), .c ({signal_5255, signal_4138}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3648 ( .a ({signal_4589, signal_4267}), .b ({signal_5221, signal_4533}), .c ({signal_5256, signal_4139}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3649 ( .a ({signal_4586, signal_4268}), .b ({signal_5222, signal_4534}), .c ({signal_5257, signal_4140}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3650 ( .a ({signal_4583, signal_4368}), .b ({signal_5814, signal_4208}), .c ({signal_5907, signal_4240}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3651 ( .a ({signal_4742, signal_4336}), .b ({signal_5473, signal_4176}), .c ({signal_5814, signal_4208}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3652 ( .a ({signal_4847, signal_4304}), .b ({signal_5261, signal_4144}), .c ({signal_5473, signal_4176}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3653 ( .a ({signal_4580, signal_4269}), .b ({signal_5223, signal_4535}), .c ({signal_5258, signal_4141}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3654 ( .a ({signal_4577, signal_4270}), .b ({signal_5224, signal_4536}), .c ({signal_5259, signal_4142}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3655 ( .a ({signal_4574, signal_4271}), .b ({signal_5225, signal_4537}), .c ({signal_5260, signal_4143}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3656 ( .a ({signal_4571, signal_4272}), .b ({signal_5226, signal_4538}), .c ({signal_5261, signal_4144}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3657 ( .a ({signal_4568, signal_4273}), .b ({signal_5227, signal_4539}), .c ({signal_5262, signal_4145}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3658 ( .a ({signal_4565, signal_4274}), .b ({signal_5228, signal_4540}), .c ({signal_5263, signal_4146}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3659 ( .a ({signal_4562, signal_4275}), .b ({signal_5229, signal_4541}), .c ({signal_5264, signal_4147}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3660 ( .a ({signal_4559, signal_4276}), .b ({signal_5230, signal_4542}), .c ({signal_5265, signal_4148}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3661 ( .a ({signal_4556, signal_4277}), .b ({signal_5231, signal_4543}), .c ({signal_5266, signal_4149}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3662 ( .a ({signal_4553, signal_4278}), .b ({signal_5232, signal_4544}), .c ({signal_5267, signal_4150}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3663 ( .a ({signal_4550, signal_4378}), .b ({signal_5815, signal_4218}), .c ({signal_5908, signal_4250}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3664 ( .a ({signal_4709, signal_4346}), .b ({signal_5474, signal_4186}), .c ({signal_5815, signal_4218}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3665 ( .a ({signal_4814, signal_4314}), .b ({signal_5268, signal_4154}), .c ({signal_5474, signal_4186}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3666 ( .a ({signal_4919, signal_4282}), .b ({signal_5236, signal_4548}), .c ({signal_5268, signal_4154}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3667 ( .a ({signal_4964, signal_3116}), .b ({1'b0, signal_393}), .c ({signal_5475, signal_4517}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3668 ( .a ({signal_4963, signal_3115}), .b ({1'b0, signal_394}), .c ({signal_5269, signal_4518}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3669 ( .a ({signal_4962, signal_3114}), .b ({1'b0, signal_4379}), .c ({signal_5816, signal_4519}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3670 ( .a ({signal_4961, signal_3113}), .b ({1'b0, signal_4380}), .c ({signal_5476, signal_4520}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3671 ( .a ({signal_4960, signal_3112}), .b ({1'b0, signal_4381}), .c ({signal_5817, signal_4521}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3672 ( .a ({signal_4959, signal_3111}), .b ({1'b0, signal_4382}), .c ({signal_5818, signal_4522}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3673 ( .a ({signal_4958, signal_3110}), .b ({1'b0, signal_4383}), .c ({signal_5270, signal_4523}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(0)) cell_3674 ( .a ({signal_4957, signal_3109}), .b ({1'b0, signal_4384}), .c ({signal_5271, signal_4524}) ) ;
    AES_step2_ANF #(.low_latency(1), .pipeline(0)) cell_4209 ( .in0 ({signal_912, signal_792, signal_4378, signal_4377, signal_4376, signal_4375, signal_4374, signal_4373, signal_4372, signal_4371, signal_4370, signal_4369, signal_4368, signal_4367, signal_4366, signal_4365, signal_4364, signal_4363, signal_4362, signal_4361, signal_4360, signal_4359, signal_4358, signal_4357, signal_4356, signal_4355, signal_4354, signal_4353, signal_4352, signal_4351, signal_4350, signal_4349, signal_4348, signal_4347, ciphertext_s0[0], ciphertext_s0[1], ciphertext_s0[2], ciphertext_s0[4], ciphertext_s0[5], ciphertext_s0[6], ciphertext_s0[7], ciphertext_s0[8], ciphertext_s0[9], ciphertext_s0[10], ciphertext_s0[12], ciphertext_s0[13], ciphertext_s0[14], ciphertext_s0[15], ciphertext_s0[16], ciphertext_s0[17], ciphertext_s0[18], ciphertext_s0[20], ciphertext_s0[21], ciphertext_s0[22], ciphertext_s0[23], ciphertext_s0[24], ciphertext_s0[25], ciphertext_s0[26], ciphertext_s0[28], ciphertext_s0[29], ciphertext_s0[30], ciphertext_s0[31], ciphertext_s0[32], ciphertext_s0[33], ciphertext_s0[34], ciphertext_s0[36], ciphertext_s0[37], ciphertext_s0[38], ciphertext_s0[39], ciphertext_s0[40], ciphertext_s0[41], ciphertext_s0[42], ciphertext_s0[44], ciphertext_s0[45], ciphertext_s0[46], ciphertext_s0[47], ciphertext_s0[48], ciphertext_s0[49], ciphertext_s0[50], ciphertext_s0[52], ciphertext_s0[53], ciphertext_s0[54], ciphertext_s0[55], ciphertext_s0[56], ciphertext_s0[57], ciphertext_s0[58], ciphertext_s0[60], ciphertext_s0[61], ciphertext_s0[62], ciphertext_s0[63], ciphertext_s0[64], ciphertext_s0[65], ciphertext_s0[66], ciphertext_s0[68], ciphertext_s0[69], ciphertext_s0[70], ciphertext_s0[71], ciphertext_s0[72], ciphertext_s0[73], ciphertext_s0[74], ciphertext_s0[76], ciphertext_s0[77], ciphertext_s0[78], ciphertext_s0[79], ciphertext_s0[80], ciphertext_s0[81], ciphertext_s0[82], ciphertext_s0[84], ciphertext_s0[85], ciphertext_s0[86], ciphertext_s0[87], ciphertext_s0[88], ciphertext_s0[89], ciphertext_s0[90], ciphertext_s0[92], ciphertext_s0[93], ciphertext_s0[94], ciphertext_s0[95], ciphertext_s0[96], ciphertext_s0[97], ciphertext_s0[98], ciphertext_s0[100], ciphertext_s0[101], ciphertext_s0[102], ciphertext_s0[103], ciphertext_s0[104], ciphertext_s0[105], ciphertext_s0[106], ciphertext_s0[108], ciphertext_s0[109], ciphertext_s0[110], ciphertext_s0[111], ciphertext_s0[112], ciphertext_s0[113], ciphertext_s0[114], ciphertext_s0[116], ciphertext_s0[117], ciphertext_s0[118], ciphertext_s0[119], ciphertext_s0[120], ciphertext_s0[121], ciphertext_s0[122], ciphertext_s0[124], ciphertext_s0[125], ciphertext_s0[126], ciphertext_s0[127], signal_2592, signal_2472, signal_2352, signal_2232, signal_2112, signal_1992, signal_1872, signal_1752, signal_1632, signal_1512, signal_1392, signal_1272, signal_1152, signal_1032}), .in1 ({signal_4934, signal_4933, signal_4550, signal_4667, signal_4700, signal_4733, signal_4766, signal_4799, signal_4832, signal_4865, signal_4898, signal_4931, signal_4583, signal_4616, signal_4643, signal_4646, signal_4649, signal_4652, signal_4655, signal_4658, signal_4661, signal_4664, signal_4670, signal_4673, signal_4676, signal_4679, signal_4682, signal_4685, signal_4688, signal_4691, signal_4694, signal_4697, signal_4703, signal_4706, ciphertext_s1[0], ciphertext_s1[1], ciphertext_s1[2], ciphertext_s1[4], ciphertext_s1[5], ciphertext_s1[6], ciphertext_s1[7], ciphertext_s1[8], ciphertext_s1[9], ciphertext_s1[10], ciphertext_s1[12], ciphertext_s1[13], ciphertext_s1[14], ciphertext_s1[15], ciphertext_s1[16], ciphertext_s1[17], ciphertext_s1[18], ciphertext_s1[20], ciphertext_s1[21], ciphertext_s1[22], ciphertext_s1[23], ciphertext_s1[24], ciphertext_s1[25], ciphertext_s1[26], ciphertext_s1[28], ciphertext_s1[29], ciphertext_s1[30], ciphertext_s1[31], ciphertext_s1[32], ciphertext_s1[33], ciphertext_s1[34], ciphertext_s1[36], ciphertext_s1[37], ciphertext_s1[38], ciphertext_s1[39], ciphertext_s1[40], ciphertext_s1[41], ciphertext_s1[42], ciphertext_s1[44], ciphertext_s1[45], ciphertext_s1[46], ciphertext_s1[47], ciphertext_s1[48], ciphertext_s1[49], ciphertext_s1[50], ciphertext_s1[52], ciphertext_s1[53], ciphertext_s1[54], ciphertext_s1[55], ciphertext_s1[56], ciphertext_s1[57], ciphertext_s1[58], ciphertext_s1[60], ciphertext_s1[61], ciphertext_s1[62], ciphertext_s1[63], ciphertext_s1[64], ciphertext_s1[65], ciphertext_s1[66], ciphertext_s1[68], ciphertext_s1[69], ciphertext_s1[70], ciphertext_s1[71], ciphertext_s1[72], ciphertext_s1[73], ciphertext_s1[74], ciphertext_s1[76], ciphertext_s1[77], ciphertext_s1[78], ciphertext_s1[79], ciphertext_s1[80], ciphertext_s1[81], ciphertext_s1[82], ciphertext_s1[84], ciphertext_s1[85], ciphertext_s1[86], ciphertext_s1[87], ciphertext_s1[88], ciphertext_s1[89], ciphertext_s1[90], ciphertext_s1[92], ciphertext_s1[93], ciphertext_s1[94], ciphertext_s1[95], ciphertext_s1[96], ciphertext_s1[97], ciphertext_s1[98], ciphertext_s1[100], ciphertext_s1[101], ciphertext_s1[102], ciphertext_s1[103], ciphertext_s1[104], ciphertext_s1[105], ciphertext_s1[106], ciphertext_s1[108], ciphertext_s1[109], ciphertext_s1[110], ciphertext_s1[111], ciphertext_s1[112], ciphertext_s1[113], ciphertext_s1[114], ciphertext_s1[116], ciphertext_s1[117], ciphertext_s1[118], ciphertext_s1[119], ciphertext_s1[120], ciphertext_s1[121], ciphertext_s1[122], ciphertext_s1[124], ciphertext_s1[125], ciphertext_s1[126], ciphertext_s1[127], signal_4948, signal_4947, signal_4946, signal_4945, signal_4944, signal_4943, signal_4942, signal_4941, signal_4940, signal_4939, signal_4938, signal_4937, signal_4936, signal_4935}), .clk (clk), .r ({Fresh[40959], Fresh[40958], Fresh[40957], Fresh[40956], Fresh[40955], Fresh[40954], Fresh[40953], Fresh[40952], Fresh[40951], Fresh[40950], Fresh[40949], Fresh[40948], Fresh[40947], Fresh[40946], Fresh[40945], Fresh[40944], Fresh[40943], Fresh[40942], Fresh[40941], Fresh[40940], Fresh[40939], Fresh[40938], Fresh[40937], Fresh[40936], Fresh[40935], Fresh[40934], Fresh[40933], Fresh[40932], Fresh[40931], Fresh[40930], Fresh[40929], Fresh[40928], Fresh[40927], Fresh[40926], Fresh[40925], Fresh[40924], Fresh[40923], Fresh[40922], Fresh[40921], Fresh[40920], Fresh[40919], Fresh[40918], Fresh[40917], Fresh[40916], Fresh[40915], Fresh[40914], Fresh[40913], Fresh[40912], Fresh[40911], Fresh[40910], Fresh[40909], Fresh[40908], Fresh[40907], Fresh[40906], Fresh[40905], Fresh[40904], Fresh[40903], Fresh[40902], Fresh[40901], Fresh[40900], Fresh[40899], Fresh[40898], Fresh[40897], Fresh[40896], Fresh[40895], Fresh[40894], Fresh[40893], Fresh[40892], Fresh[40891], Fresh[40890], Fresh[40889], Fresh[40888], Fresh[40887], Fresh[40886], Fresh[40885], Fresh[40884], Fresh[40883], Fresh[40882], Fresh[40881], Fresh[40880], Fresh[40879], Fresh[40878], Fresh[40877], Fresh[40876], Fresh[40875], Fresh[40874], Fresh[40873], Fresh[40872], Fresh[40871], Fresh[40870], Fresh[40869], Fresh[40868], Fresh[40867], Fresh[40866], Fresh[40865], Fresh[40864], Fresh[40863], Fresh[40862], Fresh[40861], Fresh[40860], Fresh[40859], Fresh[40858], Fresh[40857], Fresh[40856], Fresh[40855], Fresh[40854], Fresh[40853], Fresh[40852], Fresh[40851], Fresh[40850], Fresh[40849], Fresh[40848], Fresh[40847], Fresh[40846], Fresh[40845], Fresh[40844], Fresh[40843], Fresh[40842], Fresh[40841], Fresh[40840], Fresh[40839], Fresh[40838], Fresh[40837], Fresh[40836], Fresh[40835], Fresh[40834], Fresh[40833], Fresh[40832], Fresh[40831], Fresh[40830], Fresh[40829], Fresh[40828], Fresh[40827], Fresh[40826], Fresh[40825], Fresh[40824], Fresh[40823], Fresh[40822], Fresh[40821], Fresh[40820], Fresh[40819], Fresh[40818], Fresh[40817], Fresh[40816], Fresh[40815], Fresh[40814], Fresh[40813], Fresh[40812], Fresh[40811], Fresh[40810], Fresh[40809], Fresh[40808], Fresh[40807], Fresh[40806], Fresh[40805], Fresh[40804], Fresh[40803], Fresh[40802], Fresh[40801], Fresh[40800], Fresh[40799], Fresh[40798], Fresh[40797], Fresh[40796], Fresh[40795], Fresh[40794], Fresh[40793], Fresh[40792], Fresh[40791], Fresh[40790], Fresh[40789], Fresh[40788], Fresh[40787], Fresh[40786], Fresh[40785], Fresh[40784], Fresh[40783], Fresh[40782], Fresh[40781], Fresh[40780], Fresh[40779], Fresh[40778], Fresh[40777], Fresh[40776], Fresh[40775], Fresh[40774], Fresh[40773], Fresh[40772], Fresh[40771], Fresh[40770], Fresh[40769], Fresh[40768], Fresh[40767], Fresh[40766], Fresh[40765], Fresh[40764], Fresh[40763], Fresh[40762], Fresh[40761], Fresh[40760], Fresh[40759], Fresh[40758], Fresh[40757], Fresh[40756], Fresh[40755], Fresh[40754], Fresh[40753], Fresh[40752], Fresh[40751], Fresh[40750], Fresh[40749], Fresh[40748], Fresh[40747], Fresh[40746], Fresh[40745], Fresh[40744], Fresh[40743], Fresh[40742], Fresh[40741], Fresh[40740], Fresh[40739], Fresh[40738], Fresh[40737], Fresh[40736], Fresh[40735], Fresh[40734], Fresh[40733], Fresh[40732], Fresh[40731], Fresh[40730], Fresh[40729], Fresh[40728], Fresh[40727], Fresh[40726], Fresh[40725], Fresh[40724], Fresh[40723], Fresh[40722], Fresh[40721], Fresh[40720], Fresh[40719], Fresh[40718], Fresh[40717], Fresh[40716], Fresh[40715], Fresh[40714], Fresh[40713], Fresh[40712], Fresh[40711], Fresh[40710], Fresh[40709], Fresh[40708], Fresh[40707], Fresh[40706], Fresh[40705], Fresh[40704], Fresh[40703], Fresh[40702], Fresh[40701], Fresh[40700], Fresh[40699], Fresh[40698], Fresh[40697], Fresh[40696], Fresh[40695], Fresh[40694], Fresh[40693], Fresh[40692], Fresh[40691], Fresh[40690], Fresh[40689], Fresh[40688], Fresh[40687], Fresh[40686], Fresh[40685], Fresh[40684], Fresh[40683], Fresh[40682], Fresh[40681], Fresh[40680], Fresh[40679], Fresh[40678], Fresh[40677], Fresh[40676], Fresh[40675], Fresh[40674], Fresh[40673], Fresh[40672], Fresh[40671], Fresh[40670], Fresh[40669], Fresh[40668], Fresh[40667], Fresh[40666], Fresh[40665], Fresh[40664], Fresh[40663], Fresh[40662], Fresh[40661], Fresh[40660], Fresh[40659], Fresh[40658], Fresh[40657], Fresh[40656], Fresh[40655], Fresh[40654], Fresh[40653], Fresh[40652], Fresh[40651], Fresh[40650], Fresh[40649], Fresh[40648], Fresh[40647], Fresh[40646], Fresh[40645], Fresh[40644], Fresh[40643], Fresh[40642], Fresh[40641], Fresh[40640], Fresh[40639], Fresh[40638], Fresh[40637], Fresh[40636], Fresh[40635], Fresh[40634], Fresh[40633], Fresh[40632], Fresh[40631], Fresh[40630], Fresh[40629], Fresh[40628], Fresh[40627], Fresh[40626], Fresh[40625], Fresh[40624], Fresh[40623], Fresh[40622], Fresh[40621], Fresh[40620], Fresh[40619], Fresh[40618], Fresh[40617], Fresh[40616], Fresh[40615], Fresh[40614], Fresh[40613], Fresh[40612], Fresh[40611], Fresh[40610], Fresh[40609], Fresh[40608], Fresh[40607], Fresh[40606], Fresh[40605], Fresh[40604], Fresh[40603], Fresh[40602], Fresh[40601], Fresh[40600], Fresh[40599], Fresh[40598], Fresh[40597], Fresh[40596], Fresh[40595], Fresh[40594], Fresh[40593], Fresh[40592], Fresh[40591], Fresh[40590], Fresh[40589], Fresh[40588], Fresh[40587], Fresh[40586], Fresh[40585], Fresh[40584], Fresh[40583], Fresh[40582], Fresh[40581], Fresh[40580], Fresh[40579], Fresh[40578], Fresh[40577], Fresh[40576], Fresh[40575], Fresh[40574], Fresh[40573], Fresh[40572], Fresh[40571], Fresh[40570], Fresh[40569], Fresh[40568], Fresh[40567], Fresh[40566], Fresh[40565], Fresh[40564], Fresh[40563], Fresh[40562], Fresh[40561], Fresh[40560], Fresh[40559], Fresh[40558], Fresh[40557], Fresh[40556], Fresh[40555], Fresh[40554], Fresh[40553], Fresh[40552], Fresh[40551], Fresh[40550], Fresh[40549], Fresh[40548], Fresh[40547], Fresh[40546], Fresh[40545], Fresh[40544], Fresh[40543], Fresh[40542], Fresh[40541], Fresh[40540], Fresh[40539], Fresh[40538], Fresh[40537], Fresh[40536], Fresh[40535], Fresh[40534], Fresh[40533], Fresh[40532], Fresh[40531], Fresh[40530], Fresh[40529], Fresh[40528], Fresh[40527], Fresh[40526], Fresh[40525], Fresh[40524], Fresh[40523], Fresh[40522], Fresh[40521], Fresh[40520], Fresh[40519], Fresh[40518], Fresh[40517], Fresh[40516], Fresh[40515], Fresh[40514], Fresh[40513], Fresh[40512], Fresh[40511], Fresh[40510], Fresh[40509], Fresh[40508], Fresh[40507], Fresh[40506], Fresh[40505], Fresh[40504], Fresh[40503], Fresh[40502], Fresh[40501], Fresh[40500], Fresh[40499], Fresh[40498], Fresh[40497], Fresh[40496], Fresh[40495], Fresh[40494], Fresh[40493], Fresh[40492], Fresh[40491], Fresh[40490], Fresh[40489], Fresh[40488], Fresh[40487], Fresh[40486], Fresh[40485], Fresh[40484], Fresh[40483], Fresh[40482], Fresh[40481], Fresh[40480], Fresh[40479], Fresh[40478], Fresh[40477], Fresh[40476], Fresh[40475], Fresh[40474], Fresh[40473], Fresh[40472], Fresh[40471], Fresh[40470], Fresh[40469], Fresh[40468], Fresh[40467], Fresh[40466], Fresh[40465], Fresh[40464], Fresh[40463], Fresh[40462], Fresh[40461], Fresh[40460], Fresh[40459], Fresh[40458], Fresh[40457], Fresh[40456], Fresh[40455], Fresh[40454], Fresh[40453], Fresh[40452], Fresh[40451], Fresh[40450], Fresh[40449], Fresh[40448], Fresh[40447], Fresh[40446], Fresh[40445], Fresh[40444], Fresh[40443], Fresh[40442], Fresh[40441], Fresh[40440], Fresh[40439], Fresh[40438], Fresh[40437], Fresh[40436], Fresh[40435], Fresh[40434], Fresh[40433], Fresh[40432], Fresh[40431], Fresh[40430], Fresh[40429], Fresh[40428], Fresh[40427], Fresh[40426], Fresh[40425], Fresh[40424], Fresh[40423], Fresh[40422], Fresh[40421], Fresh[40420], Fresh[40419], Fresh[40418], Fresh[40417], Fresh[40416], Fresh[40415], Fresh[40414], Fresh[40413], Fresh[40412], Fresh[40411], Fresh[40410], Fresh[40409], Fresh[40408], Fresh[40407], Fresh[40406], Fresh[40405], Fresh[40404], Fresh[40403], Fresh[40402], Fresh[40401], Fresh[40400], Fresh[40399], Fresh[40398], Fresh[40397], Fresh[40396], Fresh[40395], Fresh[40394], Fresh[40393], Fresh[40392], Fresh[40391], Fresh[40390], Fresh[40389], Fresh[40388], Fresh[40387], Fresh[40386], Fresh[40385], Fresh[40384], Fresh[40383], Fresh[40382], Fresh[40381], Fresh[40380], Fresh[40379], Fresh[40378], Fresh[40377], Fresh[40376], Fresh[40375], Fresh[40374], Fresh[40373], Fresh[40372], Fresh[40371], Fresh[40370], Fresh[40369], Fresh[40368], Fresh[40367], Fresh[40366], Fresh[40365], Fresh[40364], Fresh[40363], Fresh[40362], Fresh[40361], Fresh[40360], Fresh[40359], Fresh[40358], Fresh[40357], Fresh[40356], Fresh[40355], Fresh[40354], Fresh[40353], Fresh[40352], Fresh[40351], Fresh[40350], Fresh[40349], Fresh[40348], Fresh[40347], Fresh[40346], Fresh[40345], Fresh[40344], Fresh[40343], Fresh[40342], Fresh[40341], Fresh[40340], Fresh[40339], Fresh[40338], Fresh[40337], Fresh[40336], Fresh[40335], Fresh[40334], Fresh[40333], Fresh[40332], Fresh[40331], Fresh[40330], Fresh[40329], Fresh[40328], Fresh[40327], Fresh[40326], Fresh[40325], Fresh[40324], Fresh[40323], Fresh[40322], Fresh[40321], Fresh[40320], Fresh[40319], Fresh[40318], Fresh[40317], Fresh[40316], Fresh[40315], Fresh[40314], Fresh[40313], Fresh[40312], Fresh[40311], Fresh[40310], Fresh[40309], Fresh[40308], Fresh[40307], Fresh[40306], Fresh[40305], Fresh[40304], Fresh[40303], Fresh[40302], Fresh[40301], Fresh[40300], Fresh[40299], Fresh[40298], Fresh[40297], Fresh[40296], Fresh[40295], Fresh[40294], Fresh[40293], Fresh[40292], Fresh[40291], Fresh[40290], Fresh[40289], Fresh[40288], Fresh[40287], Fresh[40286], Fresh[40285], Fresh[40284], Fresh[40283], Fresh[40282], Fresh[40281], Fresh[40280], Fresh[40279], Fresh[40278], Fresh[40277], Fresh[40276], Fresh[40275], Fresh[40274], Fresh[40273], Fresh[40272], Fresh[40271], Fresh[40270], Fresh[40269], Fresh[40268], Fresh[40267], Fresh[40266], Fresh[40265], Fresh[40264], Fresh[40263], Fresh[40262], Fresh[40261], Fresh[40260], Fresh[40259], Fresh[40258], Fresh[40257], Fresh[40256], Fresh[40255], Fresh[40254], Fresh[40253], Fresh[40252], Fresh[40251], Fresh[40250], Fresh[40249], Fresh[40248], Fresh[40247], Fresh[40246], Fresh[40245], Fresh[40244], Fresh[40243], Fresh[40242], Fresh[40241], Fresh[40240], Fresh[40239], Fresh[40238], Fresh[40237], Fresh[40236], Fresh[40235], Fresh[40234], Fresh[40233], Fresh[40232], Fresh[40231], Fresh[40230], Fresh[40229], Fresh[40228], Fresh[40227], Fresh[40226], Fresh[40225], Fresh[40224], Fresh[40223], Fresh[40222], Fresh[40221], Fresh[40220], Fresh[40219], Fresh[40218], Fresh[40217], Fresh[40216], Fresh[40215], Fresh[40214], Fresh[40213], Fresh[40212], Fresh[40211], Fresh[40210], Fresh[40209], Fresh[40208], Fresh[40207], Fresh[40206], Fresh[40205], Fresh[40204], Fresh[40203], Fresh[40202], Fresh[40201], Fresh[40200], Fresh[40199], Fresh[40198], Fresh[40197], Fresh[40196], Fresh[40195], Fresh[40194], Fresh[40193], Fresh[40192], Fresh[40191], Fresh[40190], Fresh[40189], Fresh[40188], Fresh[40187], Fresh[40186], Fresh[40185], Fresh[40184], Fresh[40183], Fresh[40182], Fresh[40181], Fresh[40180], Fresh[40179], Fresh[40178], Fresh[40177], Fresh[40176], Fresh[40175], Fresh[40174], Fresh[40173], Fresh[40172], Fresh[40171], Fresh[40170], Fresh[40169], Fresh[40168], Fresh[40167], Fresh[40166], Fresh[40165], Fresh[40164], Fresh[40163], Fresh[40162], Fresh[40161], Fresh[40160], Fresh[40159], Fresh[40158], Fresh[40157], Fresh[40156], Fresh[40155], Fresh[40154], Fresh[40153], Fresh[40152], Fresh[40151], Fresh[40150], Fresh[40149], Fresh[40148], Fresh[40147], Fresh[40146], Fresh[40145], Fresh[40144], Fresh[40143], Fresh[40142], Fresh[40141], Fresh[40140], Fresh[40139], Fresh[40138], Fresh[40137], Fresh[40136], Fresh[40135], Fresh[40134], Fresh[40133], Fresh[40132], Fresh[40131], Fresh[40130], Fresh[40129], Fresh[40128], Fresh[40127], Fresh[40126], Fresh[40125], Fresh[40124], Fresh[40123], Fresh[40122], Fresh[40121], Fresh[40120], Fresh[40119], Fresh[40118], Fresh[40117], Fresh[40116], Fresh[40115], Fresh[40114], Fresh[40113], Fresh[40112], Fresh[40111], Fresh[40110], Fresh[40109], Fresh[40108], Fresh[40107], Fresh[40106], Fresh[40105], Fresh[40104], Fresh[40103], Fresh[40102], Fresh[40101], Fresh[40100], Fresh[40099], Fresh[40098], Fresh[40097], Fresh[40096], Fresh[40095], Fresh[40094], Fresh[40093], Fresh[40092], Fresh[40091], Fresh[40090], Fresh[40089], Fresh[40088], Fresh[40087], Fresh[40086], Fresh[40085], Fresh[40084], Fresh[40083], Fresh[40082], Fresh[40081], Fresh[40080], Fresh[40079], Fresh[40078], Fresh[40077], Fresh[40076], Fresh[40075], Fresh[40074], Fresh[40073], Fresh[40072], Fresh[40071], Fresh[40070], Fresh[40069], Fresh[40068], Fresh[40067], Fresh[40066], Fresh[40065], Fresh[40064], Fresh[40063], Fresh[40062], Fresh[40061], Fresh[40060], Fresh[40059], Fresh[40058], Fresh[40057], Fresh[40056], Fresh[40055], Fresh[40054], Fresh[40053], Fresh[40052], Fresh[40051], Fresh[40050], Fresh[40049], Fresh[40048], Fresh[40047], Fresh[40046], Fresh[40045], Fresh[40044], Fresh[40043], Fresh[40042], Fresh[40041], Fresh[40040], Fresh[40039], Fresh[40038], Fresh[40037], Fresh[40036], Fresh[40035], Fresh[40034], Fresh[40033], Fresh[40032], Fresh[40031], Fresh[40030], Fresh[40029], Fresh[40028], Fresh[40027], Fresh[40026], Fresh[40025], Fresh[40024], Fresh[40023], Fresh[40022], Fresh[40021], Fresh[40020], Fresh[40019], Fresh[40018], Fresh[40017], Fresh[40016], Fresh[40015], Fresh[40014], Fresh[40013], Fresh[40012], Fresh[40011], Fresh[40010], Fresh[40009], Fresh[40008], Fresh[40007], Fresh[40006], Fresh[40005], Fresh[40004], Fresh[40003], Fresh[40002], Fresh[40001], Fresh[40000], Fresh[39999], Fresh[39998], Fresh[39997], Fresh[39996], Fresh[39995], Fresh[39994], Fresh[39993], Fresh[39992], Fresh[39991], Fresh[39990], Fresh[39989], Fresh[39988], Fresh[39987], Fresh[39986], Fresh[39985], Fresh[39984], Fresh[39983], Fresh[39982], Fresh[39981], Fresh[39980], Fresh[39979], Fresh[39978], Fresh[39977], Fresh[39976], Fresh[39975], Fresh[39974], Fresh[39973], Fresh[39972], Fresh[39971], Fresh[39970], Fresh[39969], Fresh[39968], Fresh[39967], Fresh[39966], Fresh[39965], Fresh[39964], Fresh[39963], Fresh[39962], Fresh[39961], Fresh[39960], Fresh[39959], Fresh[39958], Fresh[39957], Fresh[39956], Fresh[39955], Fresh[39954], Fresh[39953], Fresh[39952], Fresh[39951], Fresh[39950], Fresh[39949], Fresh[39948], Fresh[39947], Fresh[39946], Fresh[39945], Fresh[39944], Fresh[39943], Fresh[39942], Fresh[39941], Fresh[39940], Fresh[39939], Fresh[39938], Fresh[39937], Fresh[39936], Fresh[39935], Fresh[39934], Fresh[39933], Fresh[39932], Fresh[39931], Fresh[39930], Fresh[39929], Fresh[39928], Fresh[39927], Fresh[39926], Fresh[39925], Fresh[39924], Fresh[39923], Fresh[39922], Fresh[39921], Fresh[39920], Fresh[39919], Fresh[39918], Fresh[39917], Fresh[39916], Fresh[39915], Fresh[39914], Fresh[39913], Fresh[39912], Fresh[39911], Fresh[39910], Fresh[39909], Fresh[39908], Fresh[39907], Fresh[39906], Fresh[39905], Fresh[39904], Fresh[39903], Fresh[39902], Fresh[39901], Fresh[39900], Fresh[39899], Fresh[39898], Fresh[39897], Fresh[39896], Fresh[39895], Fresh[39894], Fresh[39893], Fresh[39892], Fresh[39891], Fresh[39890], Fresh[39889], Fresh[39888], Fresh[39887], Fresh[39886], Fresh[39885], Fresh[39884], Fresh[39883], Fresh[39882], Fresh[39881], Fresh[39880], Fresh[39879], Fresh[39878], Fresh[39877], Fresh[39876], Fresh[39875], Fresh[39874], Fresh[39873], Fresh[39872], Fresh[39871], Fresh[39870], Fresh[39869], Fresh[39868], Fresh[39867], Fresh[39866], Fresh[39865], Fresh[39864], Fresh[39863], Fresh[39862], Fresh[39861], Fresh[39860], Fresh[39859], Fresh[39858], Fresh[39857], Fresh[39856], Fresh[39855], Fresh[39854], Fresh[39853], Fresh[39852], Fresh[39851], Fresh[39850], Fresh[39849], Fresh[39848], Fresh[39847], Fresh[39846], Fresh[39845], Fresh[39844], Fresh[39843], Fresh[39842], Fresh[39841], Fresh[39840], Fresh[39839], Fresh[39838], Fresh[39837], Fresh[39836], Fresh[39835], Fresh[39834], Fresh[39833], Fresh[39832], Fresh[39831], Fresh[39830], Fresh[39829], Fresh[39828], Fresh[39827], Fresh[39826], Fresh[39825], Fresh[39824], Fresh[39823], Fresh[39822], Fresh[39821], Fresh[39820], Fresh[39819], Fresh[39818], Fresh[39817], Fresh[39816], Fresh[39815], Fresh[39814], Fresh[39813], Fresh[39812], Fresh[39811], Fresh[39810], Fresh[39809], Fresh[39808], Fresh[39807], Fresh[39806], Fresh[39805], Fresh[39804], Fresh[39803], Fresh[39802], Fresh[39801], Fresh[39800], Fresh[39799], Fresh[39798], Fresh[39797], Fresh[39796], Fresh[39795], Fresh[39794], Fresh[39793], Fresh[39792], Fresh[39791], Fresh[39790], Fresh[39789], Fresh[39788], Fresh[39787], Fresh[39786], Fresh[39785], Fresh[39784], Fresh[39783], Fresh[39782], Fresh[39781], Fresh[39780], Fresh[39779], Fresh[39778], Fresh[39777], Fresh[39776], Fresh[39775], Fresh[39774], Fresh[39773], Fresh[39772], Fresh[39771], Fresh[39770], Fresh[39769], Fresh[39768], Fresh[39767], Fresh[39766], Fresh[39765], Fresh[39764], Fresh[39763], Fresh[39762], Fresh[39761], Fresh[39760], Fresh[39759], Fresh[39758], Fresh[39757], Fresh[39756], Fresh[39755], Fresh[39754], Fresh[39753], Fresh[39752], Fresh[39751], Fresh[39750], Fresh[39749], Fresh[39748], Fresh[39747], Fresh[39746], Fresh[39745], Fresh[39744], Fresh[39743], Fresh[39742], Fresh[39741], Fresh[39740], Fresh[39739], Fresh[39738], Fresh[39737], Fresh[39736], Fresh[39735], Fresh[39734], Fresh[39733], Fresh[39732], Fresh[39731], Fresh[39730], Fresh[39729], Fresh[39728], Fresh[39727], Fresh[39726], Fresh[39725], Fresh[39724], Fresh[39723], Fresh[39722], Fresh[39721], Fresh[39720], Fresh[39719], Fresh[39718], Fresh[39717], Fresh[39716], Fresh[39715], Fresh[39714], Fresh[39713], Fresh[39712], Fresh[39711], Fresh[39710], Fresh[39709], Fresh[39708], Fresh[39707], Fresh[39706], Fresh[39705], Fresh[39704], Fresh[39703], Fresh[39702], Fresh[39701], Fresh[39700], Fresh[39699], Fresh[39698], Fresh[39697], Fresh[39696], Fresh[39695], Fresh[39694], Fresh[39693], Fresh[39692], Fresh[39691], Fresh[39690], Fresh[39689], Fresh[39688], Fresh[39687], Fresh[39686], Fresh[39685], Fresh[39684], Fresh[39683], Fresh[39682], Fresh[39681], Fresh[39680], Fresh[39679], Fresh[39678], Fresh[39677], Fresh[39676], Fresh[39675], Fresh[39674], Fresh[39673], Fresh[39672], Fresh[39671], Fresh[39670], Fresh[39669], Fresh[39668], Fresh[39667], Fresh[39666], Fresh[39665], Fresh[39664], Fresh[39663], Fresh[39662], Fresh[39661], Fresh[39660], Fresh[39659], Fresh[39658], Fresh[39657], Fresh[39656], Fresh[39655], Fresh[39654], Fresh[39653], Fresh[39652], Fresh[39651], Fresh[39650], Fresh[39649], Fresh[39648], Fresh[39647], Fresh[39646], Fresh[39645], Fresh[39644], Fresh[39643], Fresh[39642], Fresh[39641], Fresh[39640], Fresh[39639], Fresh[39638], Fresh[39637], Fresh[39636], Fresh[39635], Fresh[39634], Fresh[39633], Fresh[39632], Fresh[39631], Fresh[39630], Fresh[39629], Fresh[39628], Fresh[39627], Fresh[39626], Fresh[39625], Fresh[39624], Fresh[39623], Fresh[39622], Fresh[39621], Fresh[39620], Fresh[39619], Fresh[39618], Fresh[39617], Fresh[39616], Fresh[39615], Fresh[39614], Fresh[39613], Fresh[39612], Fresh[39611], Fresh[39610], Fresh[39609], Fresh[39608], Fresh[39607], Fresh[39606], Fresh[39605], Fresh[39604], Fresh[39603], Fresh[39602], Fresh[39601], Fresh[39600], Fresh[39599], Fresh[39598], Fresh[39597], Fresh[39596], Fresh[39595], Fresh[39594], Fresh[39593], Fresh[39592], Fresh[39591], Fresh[39590], Fresh[39589], Fresh[39588], Fresh[39587], Fresh[39586], Fresh[39585], Fresh[39584], Fresh[39583], Fresh[39582], Fresh[39581], Fresh[39580], Fresh[39579], Fresh[39578], Fresh[39577], Fresh[39576], Fresh[39575], Fresh[39574], Fresh[39573], Fresh[39572], Fresh[39571], Fresh[39570], Fresh[39569], Fresh[39568], Fresh[39567], Fresh[39566], Fresh[39565], Fresh[39564], Fresh[39563], Fresh[39562], Fresh[39561], Fresh[39560], Fresh[39559], Fresh[39558], Fresh[39557], Fresh[39556], Fresh[39555], Fresh[39554], Fresh[39553], Fresh[39552], Fresh[39551], Fresh[39550], Fresh[39549], Fresh[39548], Fresh[39547], Fresh[39546], Fresh[39545], Fresh[39544], Fresh[39543], Fresh[39542], Fresh[39541], Fresh[39540], Fresh[39539], Fresh[39538], Fresh[39537], Fresh[39536], Fresh[39535], Fresh[39534], Fresh[39533], Fresh[39532], Fresh[39531], Fresh[39530], Fresh[39529], Fresh[39528], Fresh[39527], Fresh[39526], Fresh[39525], Fresh[39524], Fresh[39523], Fresh[39522], Fresh[39521], Fresh[39520], Fresh[39519], Fresh[39518], Fresh[39517], Fresh[39516], Fresh[39515], Fresh[39514], Fresh[39513], Fresh[39512], Fresh[39511], Fresh[39510], Fresh[39509], Fresh[39508], Fresh[39507], Fresh[39506], Fresh[39505], Fresh[39504], Fresh[39503], Fresh[39502], Fresh[39501], Fresh[39500], Fresh[39499], Fresh[39498], Fresh[39497], Fresh[39496], Fresh[39495], Fresh[39494], Fresh[39493], Fresh[39492], Fresh[39491], Fresh[39490], Fresh[39489], Fresh[39488], Fresh[39487], Fresh[39486], Fresh[39485], Fresh[39484], Fresh[39483], Fresh[39482], Fresh[39481], Fresh[39480], Fresh[39479], Fresh[39478], Fresh[39477], Fresh[39476], Fresh[39475], Fresh[39474], Fresh[39473], Fresh[39472], Fresh[39471], Fresh[39470], Fresh[39469], Fresh[39468], Fresh[39467], Fresh[39466], Fresh[39465], Fresh[39464], Fresh[39463], Fresh[39462], Fresh[39461], Fresh[39460], Fresh[39459], Fresh[39458], Fresh[39457], Fresh[39456], Fresh[39455], Fresh[39454], Fresh[39453], Fresh[39452], Fresh[39451], Fresh[39450], Fresh[39449], Fresh[39448], Fresh[39447], Fresh[39446], Fresh[39445], Fresh[39444], Fresh[39443], Fresh[39442], Fresh[39441], Fresh[39440], Fresh[39439], Fresh[39438], Fresh[39437], Fresh[39436], Fresh[39435], Fresh[39434], Fresh[39433], Fresh[39432], Fresh[39431], Fresh[39430], Fresh[39429], Fresh[39428], Fresh[39427], Fresh[39426], Fresh[39425], Fresh[39424], Fresh[39423], Fresh[39422], Fresh[39421], Fresh[39420], Fresh[39419], Fresh[39418], Fresh[39417], Fresh[39416], Fresh[39415], Fresh[39414], Fresh[39413], Fresh[39412], Fresh[39411], Fresh[39410], Fresh[39409], Fresh[39408], Fresh[39407], Fresh[39406], Fresh[39405], Fresh[39404], Fresh[39403], Fresh[39402], Fresh[39401], Fresh[39400], Fresh[39399], Fresh[39398], Fresh[39397], Fresh[39396], Fresh[39395], Fresh[39394], Fresh[39393], Fresh[39392], Fresh[39391], Fresh[39390], Fresh[39389], Fresh[39388], Fresh[39387], Fresh[39386], Fresh[39385], Fresh[39384], Fresh[39383], Fresh[39382], Fresh[39381], Fresh[39380], Fresh[39379], Fresh[39378], Fresh[39377], Fresh[39376], Fresh[39375], Fresh[39374], Fresh[39373], Fresh[39372], Fresh[39371], Fresh[39370], Fresh[39369], Fresh[39368], Fresh[39367], Fresh[39366], Fresh[39365], Fresh[39364], Fresh[39363], Fresh[39362], Fresh[39361], Fresh[39360], Fresh[39359], Fresh[39358], Fresh[39357], Fresh[39356], Fresh[39355], Fresh[39354], Fresh[39353], Fresh[39352], Fresh[39351], Fresh[39350], Fresh[39349], Fresh[39348], Fresh[39347], Fresh[39346], Fresh[39345], Fresh[39344], Fresh[39343], Fresh[39342], Fresh[39341], Fresh[39340], Fresh[39339], Fresh[39338], Fresh[39337], Fresh[39336], Fresh[39335], Fresh[39334], Fresh[39333], Fresh[39332], Fresh[39331], Fresh[39330], Fresh[39329], Fresh[39328], Fresh[39327], Fresh[39326], Fresh[39325], Fresh[39324], Fresh[39323], Fresh[39322], Fresh[39321], Fresh[39320], Fresh[39319], Fresh[39318], Fresh[39317], Fresh[39316], Fresh[39315], Fresh[39314], Fresh[39313], Fresh[39312], Fresh[39311], Fresh[39310], Fresh[39309], Fresh[39308], Fresh[39307], Fresh[39306], Fresh[39305], Fresh[39304], Fresh[39303], Fresh[39302], Fresh[39301], Fresh[39300], Fresh[39299], Fresh[39298], Fresh[39297], Fresh[39296], Fresh[39295], Fresh[39294], Fresh[39293], Fresh[39292], Fresh[39291], Fresh[39290], Fresh[39289], Fresh[39288], Fresh[39287], Fresh[39286], Fresh[39285], Fresh[39284], Fresh[39283], Fresh[39282], Fresh[39281], Fresh[39280], Fresh[39279], Fresh[39278], Fresh[39277], Fresh[39276], Fresh[39275], Fresh[39274], Fresh[39273], Fresh[39272], Fresh[39271], Fresh[39270], Fresh[39269], Fresh[39268], Fresh[39267], Fresh[39266], Fresh[39265], Fresh[39264], Fresh[39263], Fresh[39262], Fresh[39261], Fresh[39260], Fresh[39259], Fresh[39258], Fresh[39257], Fresh[39256], Fresh[39255], Fresh[39254], Fresh[39253], Fresh[39252], Fresh[39251], Fresh[39250], Fresh[39249], Fresh[39248], Fresh[39247], Fresh[39246], Fresh[39245], Fresh[39244], Fresh[39243], Fresh[39242], Fresh[39241], Fresh[39240], Fresh[39239], Fresh[39238], Fresh[39237], Fresh[39236], Fresh[39235], Fresh[39234], Fresh[39233], Fresh[39232], Fresh[39231], Fresh[39230], Fresh[39229], Fresh[39228], Fresh[39227], Fresh[39226], Fresh[39225], Fresh[39224], Fresh[39223], Fresh[39222], Fresh[39221], Fresh[39220], Fresh[39219], Fresh[39218], Fresh[39217], Fresh[39216], Fresh[39215], Fresh[39214], Fresh[39213], Fresh[39212], Fresh[39211], Fresh[39210], Fresh[39209], Fresh[39208], Fresh[39207], Fresh[39206], Fresh[39205], Fresh[39204], Fresh[39203], Fresh[39202], Fresh[39201], Fresh[39200], Fresh[39199], Fresh[39198], Fresh[39197], Fresh[39196], Fresh[39195], Fresh[39194], Fresh[39193], Fresh[39192], Fresh[39191], Fresh[39190], Fresh[39189], Fresh[39188], Fresh[39187], Fresh[39186], Fresh[39185], Fresh[39184], Fresh[39183], Fresh[39182], Fresh[39181], Fresh[39180], Fresh[39179], Fresh[39178], Fresh[39177], Fresh[39176], Fresh[39175], Fresh[39174], Fresh[39173], Fresh[39172], Fresh[39171], Fresh[39170], Fresh[39169], Fresh[39168], Fresh[39167], Fresh[39166], Fresh[39165], Fresh[39164], Fresh[39163], Fresh[39162], Fresh[39161], Fresh[39160], Fresh[39159], Fresh[39158], Fresh[39157], Fresh[39156], Fresh[39155], Fresh[39154], Fresh[39153], Fresh[39152], Fresh[39151], Fresh[39150], Fresh[39149], Fresh[39148], Fresh[39147], Fresh[39146], Fresh[39145], Fresh[39144], Fresh[39143], Fresh[39142], Fresh[39141], Fresh[39140], Fresh[39139], Fresh[39138], Fresh[39137], Fresh[39136], Fresh[39135], Fresh[39134], Fresh[39133], Fresh[39132], Fresh[39131], Fresh[39130], Fresh[39129], Fresh[39128], Fresh[39127], Fresh[39126], Fresh[39125], Fresh[39124], Fresh[39123], Fresh[39122], Fresh[39121], Fresh[39120], Fresh[39119], Fresh[39118], Fresh[39117], Fresh[39116], Fresh[39115], Fresh[39114], Fresh[39113], Fresh[39112], Fresh[39111], Fresh[39110], Fresh[39109], Fresh[39108], Fresh[39107], Fresh[39106], Fresh[39105], Fresh[39104], Fresh[39103], Fresh[39102], Fresh[39101], Fresh[39100], Fresh[39099], Fresh[39098], Fresh[39097], Fresh[39096], Fresh[39095], Fresh[39094], Fresh[39093], Fresh[39092], Fresh[39091], Fresh[39090], Fresh[39089], Fresh[39088], Fresh[39087], Fresh[39086], Fresh[39085], Fresh[39084], Fresh[39083], Fresh[39082], Fresh[39081], Fresh[39080], Fresh[39079], Fresh[39078], Fresh[39077], Fresh[39076], Fresh[39075], Fresh[39074], Fresh[39073], Fresh[39072], Fresh[39071], Fresh[39070], Fresh[39069], Fresh[39068], Fresh[39067], Fresh[39066], Fresh[39065], Fresh[39064], Fresh[39063], Fresh[39062], Fresh[39061], Fresh[39060], Fresh[39059], Fresh[39058], Fresh[39057], Fresh[39056], Fresh[39055], Fresh[39054], Fresh[39053], Fresh[39052], Fresh[39051], Fresh[39050], Fresh[39049], Fresh[39048], Fresh[39047], Fresh[39046], Fresh[39045], Fresh[39044], Fresh[39043], Fresh[39042], Fresh[39041], Fresh[39040], Fresh[39039], Fresh[39038], Fresh[39037], Fresh[39036], Fresh[39035], Fresh[39034], Fresh[39033], Fresh[39032], Fresh[39031], Fresh[39030], Fresh[39029], Fresh[39028], Fresh[39027], Fresh[39026], Fresh[39025], Fresh[39024], Fresh[39023], Fresh[39022], Fresh[39021], Fresh[39020], Fresh[39019], Fresh[39018], Fresh[39017], Fresh[39016], Fresh[39015], Fresh[39014], Fresh[39013], Fresh[39012], Fresh[39011], Fresh[39010], Fresh[39009], Fresh[39008], Fresh[39007], Fresh[39006], Fresh[39005], Fresh[39004], Fresh[39003], Fresh[39002], Fresh[39001], Fresh[39000], Fresh[38999], Fresh[38998], Fresh[38997], Fresh[38996], Fresh[38995], Fresh[38994], Fresh[38993], Fresh[38992], Fresh[38991], Fresh[38990], Fresh[38989], Fresh[38988], Fresh[38987], Fresh[38986], Fresh[38985], Fresh[38984], Fresh[38983], Fresh[38982], Fresh[38981], Fresh[38980], Fresh[38979], Fresh[38978], Fresh[38977], Fresh[38976], Fresh[38975], Fresh[38974], Fresh[38973], Fresh[38972], Fresh[38971], Fresh[38970], Fresh[38969], Fresh[38968], Fresh[38967], Fresh[38966], Fresh[38965], Fresh[38964], Fresh[38963], Fresh[38962], Fresh[38961], Fresh[38960], Fresh[38959], Fresh[38958], Fresh[38957], Fresh[38956], Fresh[38955], Fresh[38954], Fresh[38953], Fresh[38952], Fresh[38951], Fresh[38950], Fresh[38949], Fresh[38948], Fresh[38947], Fresh[38946], Fresh[38945], Fresh[38944], Fresh[38943], Fresh[38942], Fresh[38941], Fresh[38940], Fresh[38939], Fresh[38938], Fresh[38937], Fresh[38936], Fresh[38935], Fresh[38934], Fresh[38933], Fresh[38932], Fresh[38931], Fresh[38930], Fresh[38929], Fresh[38928], Fresh[38927], Fresh[38926], Fresh[38925], Fresh[38924], Fresh[38923], Fresh[38922], Fresh[38921], Fresh[38920], Fresh[38919], Fresh[38918], Fresh[38917], Fresh[38916], Fresh[38915], Fresh[38914], Fresh[38913], Fresh[38912], Fresh[38911], Fresh[38910], Fresh[38909], Fresh[38908], Fresh[38907], Fresh[38906], Fresh[38905], Fresh[38904], Fresh[38903], Fresh[38902], Fresh[38901], Fresh[38900], Fresh[38899], Fresh[38898], Fresh[38897], Fresh[38896], Fresh[38895], Fresh[38894], Fresh[38893], Fresh[38892], Fresh[38891], Fresh[38890], Fresh[38889], Fresh[38888], Fresh[38887], Fresh[38886], Fresh[38885], Fresh[38884], Fresh[38883], Fresh[38882], Fresh[38881], Fresh[38880], Fresh[38879], Fresh[38878], Fresh[38877], Fresh[38876], Fresh[38875], Fresh[38874], Fresh[38873], Fresh[38872], Fresh[38871], Fresh[38870], Fresh[38869], Fresh[38868], Fresh[38867], Fresh[38866], Fresh[38865], Fresh[38864], Fresh[38863], Fresh[38862], Fresh[38861], Fresh[38860], Fresh[38859], Fresh[38858], Fresh[38857], Fresh[38856], Fresh[38855], Fresh[38854], Fresh[38853], Fresh[38852], Fresh[38851], Fresh[38850], Fresh[38849], Fresh[38848], Fresh[38847], Fresh[38846], Fresh[38845], Fresh[38844], Fresh[38843], Fresh[38842], Fresh[38841], Fresh[38840], Fresh[38839], Fresh[38838], Fresh[38837], Fresh[38836], Fresh[38835], Fresh[38834], Fresh[38833], Fresh[38832], Fresh[38831], Fresh[38830], Fresh[38829], Fresh[38828], Fresh[38827], Fresh[38826], Fresh[38825], Fresh[38824], Fresh[38823], Fresh[38822], Fresh[38821], Fresh[38820], Fresh[38819], Fresh[38818], Fresh[38817], Fresh[38816], Fresh[38815], Fresh[38814], Fresh[38813], Fresh[38812], Fresh[38811], Fresh[38810], Fresh[38809], Fresh[38808], Fresh[38807], Fresh[38806], Fresh[38805], Fresh[38804], Fresh[38803], Fresh[38802], Fresh[38801], Fresh[38800], Fresh[38799], Fresh[38798], Fresh[38797], Fresh[38796], Fresh[38795], Fresh[38794], Fresh[38793], Fresh[38792], Fresh[38791], Fresh[38790], Fresh[38789], Fresh[38788], Fresh[38787], Fresh[38786], Fresh[38785], Fresh[38784], Fresh[38783], Fresh[38782], Fresh[38781], Fresh[38780], Fresh[38779], Fresh[38778], Fresh[38777], Fresh[38776], Fresh[38775], Fresh[38774], Fresh[38773], Fresh[38772], Fresh[38771], Fresh[38770], Fresh[38769], Fresh[38768], Fresh[38767], Fresh[38766], Fresh[38765], Fresh[38764], Fresh[38763], Fresh[38762], Fresh[38761], Fresh[38760], Fresh[38759], Fresh[38758], Fresh[38757], Fresh[38756], Fresh[38755], Fresh[38754], Fresh[38753], Fresh[38752], Fresh[38751], Fresh[38750], Fresh[38749], Fresh[38748], Fresh[38747], Fresh[38746], Fresh[38745], Fresh[38744], Fresh[38743], Fresh[38742], Fresh[38741], Fresh[38740], Fresh[38739], Fresh[38738], Fresh[38737], Fresh[38736], Fresh[38735], Fresh[38734], Fresh[38733], Fresh[38732], Fresh[38731], Fresh[38730], Fresh[38729], Fresh[38728], Fresh[38727], Fresh[38726], Fresh[38725], Fresh[38724], Fresh[38723], Fresh[38722], Fresh[38721], Fresh[38720], Fresh[38719], Fresh[38718], Fresh[38717], Fresh[38716], Fresh[38715], Fresh[38714], Fresh[38713], Fresh[38712], Fresh[38711], Fresh[38710], Fresh[38709], Fresh[38708], Fresh[38707], Fresh[38706], Fresh[38705], Fresh[38704], Fresh[38703], Fresh[38702], Fresh[38701], Fresh[38700], Fresh[38699], Fresh[38698], Fresh[38697], Fresh[38696], Fresh[38695], Fresh[38694], Fresh[38693], Fresh[38692], Fresh[38691], Fresh[38690], Fresh[38689], Fresh[38688], Fresh[38687], Fresh[38686], Fresh[38685], Fresh[38684], Fresh[38683], Fresh[38682], Fresh[38681], Fresh[38680], Fresh[38679], Fresh[38678], Fresh[38677], Fresh[38676], Fresh[38675], Fresh[38674], Fresh[38673], Fresh[38672], Fresh[38671], Fresh[38670], Fresh[38669], Fresh[38668], Fresh[38667], Fresh[38666], Fresh[38665], Fresh[38664], Fresh[38663], Fresh[38662], Fresh[38661], Fresh[38660], Fresh[38659], Fresh[38658], Fresh[38657], Fresh[38656], Fresh[38655], Fresh[38654], Fresh[38653], Fresh[38652], Fresh[38651], Fresh[38650], Fresh[38649], Fresh[38648], Fresh[38647], Fresh[38646], Fresh[38645], Fresh[38644], Fresh[38643], Fresh[38642], Fresh[38641], Fresh[38640], Fresh[38639], Fresh[38638], Fresh[38637], Fresh[38636], Fresh[38635], Fresh[38634], Fresh[38633], Fresh[38632], Fresh[38631], Fresh[38630], Fresh[38629], Fresh[38628], Fresh[38627], Fresh[38626], Fresh[38625], Fresh[38624], Fresh[38623], Fresh[38622], Fresh[38621], Fresh[38620], Fresh[38619], Fresh[38618], Fresh[38617], Fresh[38616], Fresh[38615], Fresh[38614], Fresh[38613], Fresh[38612], Fresh[38611], Fresh[38610], Fresh[38609], Fresh[38608], Fresh[38607], Fresh[38606], Fresh[38605], Fresh[38604], Fresh[38603], Fresh[38602], Fresh[38601], Fresh[38600], Fresh[38599], Fresh[38598], Fresh[38597], Fresh[38596], Fresh[38595], Fresh[38594], Fresh[38593], Fresh[38592], Fresh[38591], Fresh[38590], Fresh[38589], Fresh[38588], Fresh[38587], Fresh[38586], Fresh[38585], Fresh[38584], Fresh[38583], Fresh[38582], Fresh[38581], Fresh[38580], Fresh[38579], Fresh[38578], Fresh[38577], Fresh[38576], Fresh[38575], Fresh[38574], Fresh[38573], Fresh[38572], Fresh[38571], Fresh[38570], Fresh[38569], Fresh[38568], Fresh[38567], Fresh[38566], Fresh[38565], Fresh[38564], Fresh[38563], Fresh[38562], Fresh[38561], Fresh[38560], Fresh[38559], Fresh[38558], Fresh[38557], Fresh[38556], Fresh[38555], Fresh[38554], Fresh[38553], Fresh[38552], Fresh[38551], Fresh[38550], Fresh[38549], Fresh[38548], Fresh[38547], Fresh[38546], Fresh[38545], Fresh[38544], Fresh[38543], Fresh[38542], Fresh[38541], Fresh[38540], Fresh[38539], Fresh[38538], Fresh[38537], Fresh[38536], Fresh[38535], Fresh[38534], Fresh[38533], Fresh[38532], Fresh[38531], Fresh[38530], Fresh[38529], Fresh[38528], Fresh[38527], Fresh[38526], Fresh[38525], Fresh[38524], Fresh[38523], Fresh[38522], Fresh[38521], Fresh[38520], Fresh[38519], Fresh[38518], Fresh[38517], Fresh[38516], Fresh[38515], Fresh[38514], Fresh[38513], Fresh[38512], Fresh[38511], Fresh[38510], Fresh[38509], Fresh[38508], Fresh[38507], Fresh[38506], Fresh[38505], Fresh[38504], Fresh[38503], Fresh[38502], Fresh[38501], Fresh[38500], Fresh[38499], Fresh[38498], Fresh[38497], Fresh[38496], Fresh[38495], Fresh[38494], Fresh[38493], Fresh[38492], Fresh[38491], Fresh[38490], Fresh[38489], Fresh[38488], Fresh[38487], Fresh[38486], Fresh[38485], Fresh[38484], Fresh[38483], Fresh[38482], Fresh[38481], Fresh[38480], Fresh[38479], Fresh[38478], Fresh[38477], Fresh[38476], Fresh[38475], Fresh[38474], Fresh[38473], Fresh[38472], Fresh[38471], Fresh[38470], Fresh[38469], Fresh[38468], Fresh[38467], Fresh[38466], Fresh[38465], Fresh[38464], Fresh[38463], Fresh[38462], Fresh[38461], Fresh[38460], Fresh[38459], Fresh[38458], Fresh[38457], Fresh[38456], Fresh[38455], Fresh[38454], Fresh[38453], Fresh[38452], Fresh[38451], Fresh[38450], Fresh[38449], Fresh[38448], Fresh[38447], Fresh[38446], Fresh[38445], Fresh[38444], Fresh[38443], Fresh[38442], Fresh[38441], Fresh[38440], Fresh[38439], Fresh[38438], Fresh[38437], Fresh[38436], Fresh[38435], Fresh[38434], Fresh[38433], Fresh[38432], Fresh[38431], Fresh[38430], Fresh[38429], Fresh[38428], Fresh[38427], Fresh[38426], Fresh[38425], Fresh[38424], Fresh[38423], Fresh[38422], Fresh[38421], Fresh[38420], Fresh[38419], Fresh[38418], Fresh[38417], Fresh[38416], Fresh[38415], Fresh[38414], Fresh[38413], Fresh[38412], Fresh[38411], Fresh[38410], Fresh[38409], Fresh[38408], Fresh[38407], Fresh[38406], Fresh[38405], Fresh[38404], Fresh[38403], Fresh[38402], Fresh[38401], Fresh[38400], Fresh[38399], Fresh[38398], Fresh[38397], Fresh[38396], Fresh[38395], Fresh[38394], Fresh[38393], Fresh[38392], Fresh[38391], Fresh[38390], Fresh[38389], Fresh[38388], Fresh[38387], Fresh[38386], Fresh[38385], Fresh[38384], Fresh[38383], Fresh[38382], Fresh[38381], Fresh[38380], Fresh[38379], Fresh[38378], Fresh[38377], Fresh[38376], Fresh[38375], Fresh[38374], Fresh[38373], Fresh[38372], Fresh[38371], Fresh[38370], Fresh[38369], Fresh[38368], Fresh[38367], Fresh[38366], Fresh[38365], Fresh[38364], Fresh[38363], Fresh[38362], Fresh[38361], Fresh[38360], Fresh[38359], Fresh[38358], Fresh[38357], Fresh[38356], Fresh[38355], Fresh[38354], Fresh[38353], Fresh[38352], Fresh[38351], Fresh[38350], Fresh[38349], Fresh[38348], Fresh[38347], Fresh[38346], Fresh[38345], Fresh[38344], Fresh[38343], Fresh[38342], Fresh[38341], Fresh[38340], Fresh[38339], Fresh[38338], Fresh[38337], Fresh[38336], Fresh[38335], Fresh[38334], Fresh[38333], Fresh[38332], Fresh[38331], Fresh[38330], Fresh[38329], Fresh[38328], Fresh[38327], Fresh[38326], Fresh[38325], Fresh[38324], Fresh[38323], Fresh[38322], Fresh[38321], Fresh[38320], Fresh[38319], Fresh[38318], Fresh[38317], Fresh[38316], Fresh[38315], Fresh[38314], Fresh[38313], Fresh[38312], Fresh[38311], Fresh[38310], Fresh[38309], Fresh[38308], Fresh[38307], Fresh[38306], Fresh[38305], Fresh[38304], Fresh[38303], Fresh[38302], Fresh[38301], Fresh[38300], Fresh[38299], Fresh[38298], Fresh[38297], Fresh[38296], Fresh[38295], Fresh[38294], Fresh[38293], Fresh[38292], Fresh[38291], Fresh[38290], Fresh[38289], Fresh[38288], Fresh[38287], Fresh[38286], Fresh[38285], Fresh[38284], Fresh[38283], Fresh[38282], Fresh[38281], Fresh[38280], Fresh[38279], Fresh[38278], Fresh[38277], Fresh[38276], Fresh[38275], Fresh[38274], Fresh[38273], Fresh[38272], Fresh[38271], Fresh[38270], Fresh[38269], Fresh[38268], Fresh[38267], Fresh[38266], Fresh[38265], Fresh[38264], Fresh[38263], Fresh[38262], Fresh[38261], Fresh[38260], Fresh[38259], Fresh[38258], Fresh[38257], Fresh[38256], Fresh[38255], Fresh[38254], Fresh[38253], Fresh[38252], Fresh[38251], Fresh[38250], Fresh[38249], Fresh[38248], Fresh[38247], Fresh[38246], Fresh[38245], Fresh[38244], Fresh[38243], Fresh[38242], Fresh[38241], Fresh[38240], Fresh[38239], Fresh[38238], Fresh[38237], Fresh[38236], Fresh[38235], Fresh[38234], Fresh[38233], Fresh[38232], Fresh[38231], Fresh[38230], Fresh[38229], Fresh[38228], Fresh[38227], Fresh[38226], Fresh[38225], Fresh[38224], Fresh[38223], Fresh[38222], Fresh[38221], Fresh[38220], Fresh[38219], Fresh[38218], Fresh[38217], Fresh[38216], Fresh[38215], Fresh[38214], Fresh[38213], Fresh[38212], Fresh[38211], Fresh[38210], Fresh[38209], Fresh[38208], Fresh[38207], Fresh[38206], Fresh[38205], Fresh[38204], Fresh[38203], Fresh[38202], Fresh[38201], Fresh[38200], Fresh[38199], Fresh[38198], Fresh[38197], Fresh[38196], Fresh[38195], Fresh[38194], Fresh[38193], Fresh[38192], Fresh[38191], Fresh[38190], Fresh[38189], Fresh[38188], Fresh[38187], Fresh[38186], Fresh[38185], Fresh[38184], Fresh[38183], Fresh[38182], Fresh[38181], Fresh[38180], Fresh[38179], Fresh[38178], Fresh[38177], Fresh[38176], Fresh[38175], Fresh[38174], Fresh[38173], Fresh[38172], Fresh[38171], Fresh[38170], Fresh[38169], Fresh[38168], Fresh[38167], Fresh[38166], Fresh[38165], Fresh[38164], Fresh[38163], Fresh[38162], Fresh[38161], Fresh[38160], Fresh[38159], Fresh[38158], Fresh[38157], Fresh[38156], Fresh[38155], Fresh[38154], Fresh[38153], Fresh[38152], Fresh[38151], Fresh[38150], Fresh[38149], Fresh[38148], Fresh[38147], Fresh[38146], Fresh[38145], Fresh[38144], Fresh[38143], Fresh[38142], Fresh[38141], Fresh[38140], Fresh[38139], Fresh[38138], Fresh[38137], Fresh[38136], Fresh[38135], Fresh[38134], Fresh[38133], Fresh[38132], Fresh[38131], Fresh[38130], Fresh[38129], Fresh[38128], Fresh[38127], Fresh[38126], Fresh[38125], Fresh[38124], Fresh[38123], Fresh[38122], Fresh[38121], Fresh[38120], Fresh[38119], Fresh[38118], Fresh[38117], Fresh[38116], Fresh[38115], Fresh[38114], Fresh[38113], Fresh[38112], Fresh[38111], Fresh[38110], Fresh[38109], Fresh[38108], Fresh[38107], Fresh[38106], Fresh[38105], Fresh[38104], Fresh[38103], Fresh[38102], Fresh[38101], Fresh[38100], Fresh[38099], Fresh[38098], Fresh[38097], Fresh[38096], Fresh[38095], Fresh[38094], Fresh[38093], Fresh[38092], Fresh[38091], Fresh[38090], Fresh[38089], Fresh[38088], Fresh[38087], Fresh[38086], Fresh[38085], Fresh[38084], Fresh[38083], Fresh[38082], Fresh[38081], Fresh[38080], Fresh[38079], Fresh[38078], Fresh[38077], Fresh[38076], Fresh[38075], Fresh[38074], Fresh[38073], Fresh[38072], Fresh[38071], Fresh[38070], Fresh[38069], Fresh[38068], Fresh[38067], Fresh[38066], Fresh[38065], Fresh[38064], Fresh[38063], Fresh[38062], Fresh[38061], Fresh[38060], Fresh[38059], Fresh[38058], Fresh[38057], Fresh[38056], Fresh[38055], Fresh[38054], Fresh[38053], Fresh[38052], Fresh[38051], Fresh[38050], Fresh[38049], Fresh[38048], Fresh[38047], Fresh[38046], Fresh[38045], Fresh[38044], Fresh[38043], Fresh[38042], Fresh[38041], Fresh[38040], Fresh[38039], Fresh[38038], Fresh[38037], Fresh[38036], Fresh[38035], Fresh[38034], Fresh[38033], Fresh[38032], Fresh[38031], Fresh[38030], Fresh[38029], Fresh[38028], Fresh[38027], Fresh[38026], Fresh[38025], Fresh[38024], Fresh[38023], Fresh[38022], Fresh[38021], Fresh[38020], Fresh[38019], Fresh[38018], Fresh[38017], Fresh[38016], Fresh[38015], Fresh[38014], Fresh[38013], Fresh[38012], Fresh[38011], Fresh[38010], Fresh[38009], Fresh[38008], Fresh[38007], Fresh[38006], Fresh[38005], Fresh[38004], Fresh[38003], Fresh[38002], Fresh[38001], Fresh[38000], Fresh[37999], Fresh[37998], Fresh[37997], Fresh[37996], Fresh[37995], Fresh[37994], Fresh[37993], Fresh[37992], Fresh[37991], Fresh[37990], Fresh[37989], Fresh[37988], Fresh[37987], Fresh[37986], Fresh[37985], Fresh[37984], Fresh[37983], Fresh[37982], Fresh[37981], Fresh[37980], Fresh[37979], Fresh[37978], Fresh[37977], Fresh[37976], Fresh[37975], Fresh[37974], Fresh[37973], Fresh[37972], Fresh[37971], Fresh[37970], Fresh[37969], Fresh[37968], Fresh[37967], Fresh[37966], Fresh[37965], Fresh[37964], Fresh[37963], Fresh[37962], Fresh[37961], Fresh[37960], Fresh[37959], Fresh[37958], Fresh[37957], Fresh[37956], Fresh[37955], Fresh[37954], Fresh[37953], Fresh[37952], Fresh[37951], Fresh[37950], Fresh[37949], Fresh[37948], Fresh[37947], Fresh[37946], Fresh[37945], Fresh[37944], Fresh[37943], Fresh[37942], Fresh[37941], Fresh[37940], Fresh[37939], Fresh[37938], Fresh[37937], Fresh[37936], Fresh[37935], Fresh[37934], Fresh[37933], Fresh[37932], Fresh[37931], Fresh[37930], Fresh[37929], Fresh[37928], Fresh[37927], Fresh[37926], Fresh[37925], Fresh[37924], Fresh[37923], Fresh[37922], Fresh[37921], Fresh[37920], Fresh[37919], Fresh[37918], Fresh[37917], Fresh[37916], Fresh[37915], Fresh[37914], Fresh[37913], Fresh[37912], Fresh[37911], Fresh[37910], Fresh[37909], Fresh[37908], Fresh[37907], Fresh[37906], Fresh[37905], Fresh[37904], Fresh[37903], Fresh[37902], Fresh[37901], Fresh[37900], Fresh[37899], Fresh[37898], Fresh[37897], Fresh[37896], Fresh[37895], Fresh[37894], Fresh[37893], Fresh[37892], Fresh[37891], Fresh[37890], Fresh[37889], Fresh[37888], Fresh[37887], Fresh[37886], Fresh[37885], Fresh[37884], Fresh[37883], Fresh[37882], Fresh[37881], Fresh[37880], Fresh[37879], Fresh[37878], Fresh[37877], Fresh[37876], Fresh[37875], Fresh[37874], Fresh[37873], Fresh[37872], Fresh[37871], Fresh[37870], Fresh[37869], Fresh[37868], Fresh[37867], Fresh[37866], Fresh[37865], Fresh[37864], Fresh[37863], Fresh[37862], Fresh[37861], Fresh[37860], Fresh[37859], Fresh[37858], Fresh[37857], Fresh[37856], Fresh[37855], Fresh[37854], Fresh[37853], Fresh[37852], Fresh[37851], Fresh[37850], Fresh[37849], Fresh[37848], Fresh[37847], Fresh[37846], Fresh[37845], Fresh[37844], Fresh[37843], Fresh[37842], Fresh[37841], Fresh[37840], Fresh[37839], Fresh[37838], Fresh[37837], Fresh[37836], Fresh[37835], Fresh[37834], Fresh[37833], Fresh[37832], Fresh[37831], Fresh[37830], Fresh[37829], Fresh[37828], Fresh[37827], Fresh[37826], Fresh[37825], Fresh[37824], Fresh[37823], Fresh[37822], Fresh[37821], Fresh[37820], Fresh[37819], Fresh[37818], Fresh[37817], Fresh[37816], Fresh[37815], Fresh[37814], Fresh[37813], Fresh[37812], Fresh[37811], Fresh[37810], Fresh[37809], Fresh[37808], Fresh[37807], Fresh[37806], Fresh[37805], Fresh[37804], Fresh[37803], Fresh[37802], Fresh[37801], Fresh[37800], Fresh[37799], Fresh[37798], Fresh[37797], Fresh[37796], Fresh[37795], Fresh[37794], Fresh[37793], Fresh[37792], Fresh[37791], Fresh[37790], Fresh[37789], Fresh[37788], Fresh[37787], Fresh[37786], Fresh[37785], Fresh[37784], Fresh[37783], Fresh[37782], Fresh[37781], Fresh[37780], Fresh[37779], Fresh[37778], Fresh[37777], Fresh[37776], Fresh[37775], Fresh[37774], Fresh[37773], Fresh[37772], Fresh[37771], Fresh[37770], Fresh[37769], Fresh[37768], Fresh[37767], Fresh[37766], Fresh[37765], Fresh[37764], Fresh[37763], Fresh[37762], Fresh[37761], Fresh[37760], Fresh[37759], Fresh[37758], Fresh[37757], Fresh[37756], Fresh[37755], Fresh[37754], Fresh[37753], Fresh[37752], Fresh[37751], Fresh[37750], Fresh[37749], Fresh[37748], Fresh[37747], Fresh[37746], Fresh[37745], Fresh[37744], Fresh[37743], Fresh[37742], Fresh[37741], Fresh[37740], Fresh[37739], Fresh[37738], Fresh[37737], Fresh[37736], Fresh[37735], Fresh[37734], Fresh[37733], Fresh[37732], Fresh[37731], Fresh[37730], Fresh[37729], Fresh[37728], Fresh[37727], Fresh[37726], Fresh[37725], Fresh[37724], Fresh[37723], Fresh[37722], Fresh[37721], Fresh[37720], Fresh[37719], Fresh[37718], Fresh[37717], Fresh[37716], Fresh[37715], Fresh[37714], Fresh[37713], Fresh[37712], Fresh[37711], Fresh[37710], Fresh[37709], Fresh[37708], Fresh[37707], Fresh[37706], Fresh[37705], Fresh[37704], Fresh[37703], Fresh[37702], Fresh[37701], Fresh[37700], Fresh[37699], Fresh[37698], Fresh[37697], Fresh[37696], Fresh[37695], Fresh[37694], Fresh[37693], Fresh[37692], Fresh[37691], Fresh[37690], Fresh[37689], Fresh[37688], Fresh[37687], Fresh[37686], Fresh[37685], Fresh[37684], Fresh[37683], Fresh[37682], Fresh[37681], Fresh[37680], Fresh[37679], Fresh[37678], Fresh[37677], Fresh[37676], Fresh[37675], Fresh[37674], Fresh[37673], Fresh[37672], Fresh[37671], Fresh[37670], Fresh[37669], Fresh[37668], Fresh[37667], Fresh[37666], Fresh[37665], Fresh[37664], Fresh[37663], Fresh[37662], Fresh[37661], Fresh[37660], Fresh[37659], Fresh[37658], Fresh[37657], Fresh[37656], Fresh[37655], Fresh[37654], Fresh[37653], Fresh[37652], Fresh[37651], Fresh[37650], Fresh[37649], Fresh[37648], Fresh[37647], Fresh[37646], Fresh[37645], Fresh[37644], Fresh[37643], Fresh[37642], Fresh[37641], Fresh[37640], Fresh[37639], Fresh[37638], Fresh[37637], Fresh[37636], Fresh[37635], Fresh[37634], Fresh[37633], Fresh[37632], Fresh[37631], Fresh[37630], Fresh[37629], Fresh[37628], Fresh[37627], Fresh[37626], Fresh[37625], Fresh[37624], Fresh[37623], Fresh[37622], Fresh[37621], Fresh[37620], Fresh[37619], Fresh[37618], Fresh[37617], Fresh[37616], Fresh[37615], Fresh[37614], Fresh[37613], Fresh[37612], Fresh[37611], Fresh[37610], Fresh[37609], Fresh[37608], Fresh[37607], Fresh[37606], Fresh[37605], Fresh[37604], Fresh[37603], Fresh[37602], Fresh[37601], Fresh[37600], Fresh[37599], Fresh[37598], Fresh[37597], Fresh[37596], Fresh[37595], Fresh[37594], Fresh[37593], Fresh[37592], Fresh[37591], Fresh[37590], Fresh[37589], Fresh[37588], Fresh[37587], Fresh[37586], Fresh[37585], Fresh[37584], Fresh[37583], Fresh[37582], Fresh[37581], Fresh[37580], Fresh[37579], Fresh[37578], Fresh[37577], Fresh[37576], Fresh[37575], Fresh[37574], Fresh[37573], Fresh[37572], Fresh[37571], Fresh[37570], Fresh[37569], Fresh[37568], Fresh[37567], Fresh[37566], Fresh[37565], Fresh[37564], Fresh[37563], Fresh[37562], Fresh[37561], Fresh[37560], Fresh[37559], Fresh[37558], Fresh[37557], Fresh[37556], Fresh[37555], Fresh[37554], Fresh[37553], Fresh[37552], Fresh[37551], Fresh[37550], Fresh[37549], Fresh[37548], Fresh[37547], Fresh[37546], Fresh[37545], Fresh[37544], Fresh[37543], Fresh[37542], Fresh[37541], Fresh[37540], Fresh[37539], Fresh[37538], Fresh[37537], Fresh[37536], Fresh[37535], Fresh[37534], Fresh[37533], Fresh[37532], Fresh[37531], Fresh[37530], Fresh[37529], Fresh[37528], Fresh[37527], Fresh[37526], Fresh[37525], Fresh[37524], Fresh[37523], Fresh[37522], Fresh[37521], Fresh[37520], Fresh[37519], Fresh[37518], Fresh[37517], Fresh[37516], Fresh[37515], Fresh[37514], Fresh[37513], Fresh[37512], Fresh[37511], Fresh[37510], Fresh[37509], Fresh[37508], Fresh[37507], Fresh[37506], Fresh[37505], Fresh[37504], Fresh[37503], Fresh[37502], Fresh[37501], Fresh[37500], Fresh[37499], Fresh[37498], Fresh[37497], Fresh[37496], Fresh[37495], Fresh[37494], Fresh[37493], Fresh[37492], Fresh[37491], Fresh[37490], Fresh[37489], Fresh[37488], Fresh[37487], Fresh[37486], Fresh[37485], Fresh[37484], Fresh[37483], Fresh[37482], Fresh[37481], Fresh[37480], Fresh[37479], Fresh[37478], Fresh[37477], Fresh[37476], Fresh[37475], Fresh[37474], Fresh[37473], Fresh[37472], Fresh[37471], Fresh[37470], Fresh[37469], Fresh[37468], Fresh[37467], Fresh[37466], Fresh[37465], Fresh[37464], Fresh[37463], Fresh[37462], Fresh[37461], Fresh[37460], Fresh[37459], Fresh[37458], Fresh[37457], Fresh[37456], Fresh[37455], Fresh[37454], Fresh[37453], Fresh[37452], Fresh[37451], Fresh[37450], Fresh[37449], Fresh[37448], Fresh[37447], Fresh[37446], Fresh[37445], Fresh[37444], Fresh[37443], Fresh[37442], Fresh[37441], Fresh[37440], Fresh[37439], Fresh[37438], Fresh[37437], Fresh[37436], Fresh[37435], Fresh[37434], Fresh[37433], Fresh[37432], Fresh[37431], Fresh[37430], Fresh[37429], Fresh[37428], Fresh[37427], Fresh[37426], Fresh[37425], Fresh[37424], Fresh[37423], Fresh[37422], Fresh[37421], Fresh[37420], Fresh[37419], Fresh[37418], Fresh[37417], Fresh[37416], Fresh[37415], Fresh[37414], Fresh[37413], Fresh[37412], Fresh[37411], Fresh[37410], Fresh[37409], Fresh[37408], Fresh[37407], Fresh[37406], Fresh[37405], Fresh[37404], Fresh[37403], Fresh[37402], Fresh[37401], Fresh[37400], Fresh[37399], Fresh[37398], Fresh[37397], Fresh[37396], Fresh[37395], Fresh[37394], Fresh[37393], Fresh[37392], Fresh[37391], Fresh[37390], Fresh[37389], Fresh[37388], Fresh[37387], Fresh[37386], Fresh[37385], Fresh[37384], Fresh[37383], Fresh[37382], Fresh[37381], Fresh[37380], Fresh[37379], Fresh[37378], Fresh[37377], Fresh[37376], Fresh[37375], Fresh[37374], Fresh[37373], Fresh[37372], Fresh[37371], Fresh[37370], Fresh[37369], Fresh[37368], Fresh[37367], Fresh[37366], Fresh[37365], Fresh[37364], Fresh[37363], Fresh[37362], Fresh[37361], Fresh[37360], Fresh[37359], Fresh[37358], Fresh[37357], Fresh[37356], Fresh[37355], Fresh[37354], Fresh[37353], Fresh[37352], Fresh[37351], Fresh[37350], Fresh[37349], Fresh[37348], Fresh[37347], Fresh[37346], Fresh[37345], Fresh[37344], Fresh[37343], Fresh[37342], Fresh[37341], Fresh[37340], Fresh[37339], Fresh[37338], Fresh[37337], Fresh[37336], Fresh[37335], Fresh[37334], Fresh[37333], Fresh[37332], Fresh[37331], Fresh[37330], Fresh[37329], Fresh[37328], Fresh[37327], Fresh[37326], Fresh[37325], Fresh[37324], Fresh[37323], Fresh[37322], Fresh[37321], Fresh[37320], Fresh[37319], Fresh[37318], Fresh[37317], Fresh[37316], Fresh[37315], Fresh[37314], Fresh[37313], Fresh[37312], Fresh[37311], Fresh[37310], Fresh[37309], Fresh[37308], Fresh[37307], Fresh[37306], Fresh[37305], Fresh[37304], Fresh[37303], Fresh[37302], Fresh[37301], Fresh[37300], Fresh[37299], Fresh[37298], Fresh[37297], Fresh[37296], Fresh[37295], Fresh[37294], Fresh[37293], Fresh[37292], Fresh[37291], Fresh[37290], Fresh[37289], Fresh[37288], Fresh[37287], Fresh[37286], Fresh[37285], Fresh[37284], Fresh[37283], Fresh[37282], Fresh[37281], Fresh[37280], Fresh[37279], Fresh[37278], Fresh[37277], Fresh[37276], Fresh[37275], Fresh[37274], Fresh[37273], Fresh[37272], Fresh[37271], Fresh[37270], Fresh[37269], Fresh[37268], Fresh[37267], Fresh[37266], Fresh[37265], Fresh[37264], Fresh[37263], Fresh[37262], Fresh[37261], Fresh[37260], Fresh[37259], Fresh[37258], Fresh[37257], Fresh[37256], Fresh[37255], Fresh[37254], Fresh[37253], Fresh[37252], Fresh[37251], Fresh[37250], Fresh[37249], Fresh[37248], Fresh[37247], Fresh[37246], Fresh[37245], Fresh[37244], Fresh[37243], Fresh[37242], Fresh[37241], Fresh[37240], Fresh[37239], Fresh[37238], Fresh[37237], Fresh[37236], Fresh[37235], Fresh[37234], Fresh[37233], Fresh[37232], Fresh[37231], Fresh[37230], Fresh[37229], Fresh[37228], Fresh[37227], Fresh[37226], Fresh[37225], Fresh[37224], Fresh[37223], Fresh[37222], Fresh[37221], Fresh[37220], Fresh[37219], Fresh[37218], Fresh[37217], Fresh[37216], Fresh[37215], Fresh[37214], Fresh[37213], Fresh[37212], Fresh[37211], Fresh[37210], Fresh[37209], Fresh[37208], Fresh[37207], Fresh[37206], Fresh[37205], Fresh[37204], Fresh[37203], Fresh[37202], Fresh[37201], Fresh[37200], Fresh[37199], Fresh[37198], Fresh[37197], Fresh[37196], Fresh[37195], Fresh[37194], Fresh[37193], Fresh[37192], Fresh[37191], Fresh[37190], Fresh[37189], Fresh[37188], Fresh[37187], Fresh[37186], Fresh[37185], Fresh[37184], Fresh[37183], Fresh[37182], Fresh[37181], Fresh[37180], Fresh[37179], Fresh[37178], Fresh[37177], Fresh[37176], Fresh[37175], Fresh[37174], Fresh[37173], Fresh[37172], Fresh[37171], Fresh[37170], Fresh[37169], Fresh[37168], Fresh[37167], Fresh[37166], Fresh[37165], Fresh[37164], Fresh[37163], Fresh[37162], Fresh[37161], Fresh[37160], Fresh[37159], Fresh[37158], Fresh[37157], Fresh[37156], Fresh[37155], Fresh[37154], Fresh[37153], Fresh[37152], Fresh[37151], Fresh[37150], Fresh[37149], Fresh[37148], Fresh[37147], Fresh[37146], Fresh[37145], Fresh[37144], Fresh[37143], Fresh[37142], Fresh[37141], Fresh[37140], Fresh[37139], Fresh[37138], Fresh[37137], Fresh[37136], Fresh[37135], Fresh[37134], Fresh[37133], Fresh[37132], Fresh[37131], Fresh[37130], Fresh[37129], Fresh[37128], Fresh[37127], Fresh[37126], Fresh[37125], Fresh[37124], Fresh[37123], Fresh[37122], Fresh[37121], Fresh[37120], Fresh[37119], Fresh[37118], Fresh[37117], Fresh[37116], Fresh[37115], Fresh[37114], Fresh[37113], Fresh[37112], Fresh[37111], Fresh[37110], Fresh[37109], Fresh[37108], Fresh[37107], Fresh[37106], Fresh[37105], Fresh[37104], Fresh[37103], Fresh[37102], Fresh[37101], Fresh[37100], Fresh[37099], Fresh[37098], Fresh[37097], Fresh[37096], Fresh[37095], Fresh[37094], Fresh[37093], Fresh[37092], Fresh[37091], Fresh[37090], Fresh[37089], Fresh[37088], Fresh[37087], Fresh[37086], Fresh[37085], Fresh[37084], Fresh[37083], Fresh[37082], Fresh[37081], Fresh[37080], Fresh[37079], Fresh[37078], Fresh[37077], Fresh[37076], Fresh[37075], Fresh[37074], Fresh[37073], Fresh[37072], Fresh[37071], Fresh[37070], Fresh[37069], Fresh[37068], Fresh[37067], Fresh[37066], Fresh[37065], Fresh[37064], Fresh[37063], Fresh[37062], Fresh[37061], Fresh[37060], Fresh[37059], Fresh[37058], Fresh[37057], Fresh[37056], Fresh[37055], Fresh[37054], Fresh[37053], Fresh[37052], Fresh[37051], Fresh[37050], Fresh[37049], Fresh[37048], Fresh[37047], Fresh[37046], Fresh[37045], Fresh[37044], Fresh[37043], Fresh[37042], Fresh[37041], Fresh[37040], Fresh[37039], Fresh[37038], Fresh[37037], Fresh[37036], Fresh[37035], Fresh[37034], Fresh[37033], Fresh[37032], Fresh[37031], Fresh[37030], Fresh[37029], Fresh[37028], Fresh[37027], Fresh[37026], Fresh[37025], Fresh[37024], Fresh[37023], Fresh[37022], Fresh[37021], Fresh[37020], Fresh[37019], Fresh[37018], Fresh[37017], Fresh[37016], Fresh[37015], Fresh[37014], Fresh[37013], Fresh[37012], Fresh[37011], Fresh[37010], Fresh[37009], Fresh[37008], Fresh[37007], Fresh[37006], Fresh[37005], Fresh[37004], Fresh[37003], Fresh[37002], Fresh[37001], Fresh[37000], Fresh[36999], Fresh[36998], Fresh[36997], Fresh[36996], Fresh[36995], Fresh[36994], Fresh[36993], Fresh[36992], Fresh[36991], Fresh[36990], Fresh[36989], Fresh[36988], Fresh[36987], Fresh[36986], Fresh[36985], Fresh[36984], Fresh[36983], Fresh[36982], Fresh[36981], Fresh[36980], Fresh[36979], Fresh[36978], Fresh[36977], Fresh[36976], Fresh[36975], Fresh[36974], Fresh[36973], Fresh[36972], Fresh[36971], Fresh[36970], Fresh[36969], Fresh[36968], Fresh[36967], Fresh[36966], Fresh[36965], Fresh[36964], Fresh[36963], Fresh[36962], Fresh[36961], Fresh[36960], Fresh[36959], Fresh[36958], Fresh[36957], Fresh[36956], Fresh[36955], Fresh[36954], Fresh[36953], Fresh[36952], Fresh[36951], Fresh[36950], Fresh[36949], Fresh[36948], Fresh[36947], Fresh[36946], Fresh[36945], Fresh[36944], Fresh[36943], Fresh[36942], Fresh[36941], Fresh[36940], Fresh[36939], Fresh[36938], Fresh[36937], Fresh[36936], Fresh[36935], Fresh[36934], Fresh[36933], Fresh[36932], Fresh[36931], Fresh[36930], Fresh[36929], Fresh[36928], Fresh[36927], Fresh[36926], Fresh[36925], Fresh[36924], Fresh[36923], Fresh[36922], Fresh[36921], Fresh[36920], Fresh[36919], Fresh[36918], Fresh[36917], Fresh[36916], Fresh[36915], Fresh[36914], Fresh[36913], Fresh[36912], Fresh[36911], Fresh[36910], Fresh[36909], Fresh[36908], Fresh[36907], Fresh[36906], Fresh[36905], Fresh[36904], Fresh[36903], Fresh[36902], Fresh[36901], Fresh[36900], Fresh[36899], Fresh[36898], Fresh[36897], Fresh[36896], Fresh[36895], Fresh[36894], Fresh[36893], Fresh[36892], Fresh[36891], Fresh[36890], Fresh[36889], Fresh[36888], Fresh[36887], Fresh[36886], Fresh[36885], Fresh[36884], Fresh[36883], Fresh[36882], Fresh[36881], Fresh[36880], Fresh[36879], Fresh[36878], Fresh[36877], Fresh[36876], Fresh[36875], Fresh[36874], Fresh[36873], Fresh[36872], Fresh[36871], Fresh[36870], Fresh[36869], Fresh[36868], Fresh[36867], Fresh[36866], Fresh[36865], Fresh[36864], Fresh[36863], Fresh[36862], Fresh[36861], Fresh[36860], Fresh[36859], Fresh[36858], Fresh[36857], Fresh[36856], Fresh[36855], Fresh[36854], Fresh[36853], Fresh[36852], Fresh[36851], Fresh[36850], Fresh[36849], Fresh[36848], Fresh[36847], Fresh[36846], Fresh[36845], Fresh[36844], Fresh[36843], Fresh[36842], Fresh[36841], Fresh[36840], Fresh[36839], Fresh[36838], Fresh[36837], Fresh[36836], Fresh[36835], Fresh[36834], Fresh[36833], Fresh[36832], Fresh[36831], Fresh[36830], Fresh[36829], Fresh[36828], Fresh[36827], Fresh[36826], Fresh[36825], Fresh[36824], Fresh[36823], Fresh[36822], Fresh[36821], Fresh[36820], Fresh[36819], Fresh[36818], Fresh[36817], Fresh[36816], Fresh[36815], Fresh[36814], Fresh[36813], Fresh[36812], Fresh[36811], Fresh[36810], Fresh[36809], Fresh[36808], Fresh[36807], Fresh[36806], Fresh[36805], Fresh[36804], Fresh[36803], Fresh[36802], Fresh[36801], Fresh[36800], Fresh[36799], Fresh[36798], Fresh[36797], Fresh[36796], Fresh[36795], Fresh[36794], Fresh[36793], Fresh[36792], Fresh[36791], Fresh[36790], Fresh[36789], Fresh[36788], Fresh[36787], Fresh[36786], Fresh[36785], Fresh[36784], Fresh[36783], Fresh[36782], Fresh[36781], Fresh[36780], Fresh[36779], Fresh[36778], Fresh[36777], Fresh[36776], Fresh[36775], Fresh[36774], Fresh[36773], Fresh[36772], Fresh[36771], Fresh[36770], Fresh[36769], Fresh[36768], Fresh[36767], Fresh[36766], Fresh[36765], Fresh[36764], Fresh[36763], Fresh[36762], Fresh[36761], Fresh[36760], Fresh[36759], Fresh[36758], Fresh[36757], Fresh[36756], Fresh[36755], Fresh[36754], Fresh[36753], Fresh[36752], Fresh[36751], Fresh[36750], Fresh[36749], Fresh[36748], Fresh[36747], Fresh[36746], Fresh[36745], Fresh[36744], Fresh[36743], Fresh[36742], Fresh[36741], Fresh[36740], Fresh[36739], Fresh[36738], Fresh[36737], Fresh[36736], Fresh[36735], Fresh[36734], Fresh[36733], Fresh[36732], Fresh[36731], Fresh[36730], Fresh[36729], Fresh[36728], Fresh[36727], Fresh[36726], Fresh[36725], Fresh[36724], Fresh[36723], Fresh[36722], Fresh[36721], Fresh[36720], Fresh[36719], Fresh[36718], Fresh[36717], Fresh[36716], Fresh[36715], Fresh[36714], Fresh[36713], Fresh[36712], Fresh[36711], Fresh[36710], Fresh[36709], Fresh[36708], Fresh[36707], Fresh[36706], Fresh[36705], Fresh[36704], Fresh[36703], Fresh[36702], Fresh[36701], Fresh[36700], Fresh[36699], Fresh[36698], Fresh[36697], Fresh[36696], Fresh[36695], Fresh[36694], Fresh[36693], Fresh[36692], Fresh[36691], Fresh[36690], Fresh[36689], Fresh[36688], Fresh[36687], Fresh[36686], Fresh[36685], Fresh[36684], Fresh[36683], Fresh[36682], Fresh[36681], Fresh[36680], Fresh[36679], Fresh[36678], Fresh[36677], Fresh[36676], Fresh[36675], Fresh[36674], Fresh[36673], Fresh[36672], Fresh[36671], Fresh[36670], Fresh[36669], Fresh[36668], Fresh[36667], Fresh[36666], Fresh[36665], Fresh[36664], Fresh[36663], Fresh[36662], Fresh[36661], Fresh[36660], Fresh[36659], Fresh[36658], Fresh[36657], Fresh[36656], Fresh[36655], Fresh[36654], Fresh[36653], Fresh[36652], Fresh[36651], Fresh[36650], Fresh[36649], Fresh[36648], Fresh[36647], Fresh[36646], Fresh[36645], Fresh[36644], Fresh[36643], Fresh[36642], Fresh[36641], Fresh[36640], Fresh[36639], Fresh[36638], Fresh[36637], Fresh[36636], Fresh[36635], Fresh[36634], Fresh[36633], Fresh[36632], Fresh[36631], Fresh[36630], Fresh[36629], Fresh[36628], Fresh[36627], Fresh[36626], Fresh[36625], Fresh[36624], Fresh[36623], Fresh[36622], Fresh[36621], Fresh[36620], Fresh[36619], Fresh[36618], Fresh[36617], Fresh[36616], Fresh[36615], Fresh[36614], Fresh[36613], Fresh[36612], Fresh[36611], Fresh[36610], Fresh[36609], Fresh[36608], Fresh[36607], Fresh[36606], Fresh[36605], Fresh[36604], Fresh[36603], Fresh[36602], Fresh[36601], Fresh[36600], Fresh[36599], Fresh[36598], Fresh[36597], Fresh[36596], Fresh[36595], Fresh[36594], Fresh[36593], Fresh[36592], Fresh[36591], Fresh[36590], Fresh[36589], Fresh[36588], Fresh[36587], Fresh[36586], Fresh[36585], Fresh[36584], Fresh[36583], Fresh[36582], Fresh[36581], Fresh[36580], Fresh[36579], Fresh[36578], Fresh[36577], Fresh[36576], Fresh[36575], Fresh[36574], Fresh[36573], Fresh[36572], Fresh[36571], Fresh[36570], Fresh[36569], Fresh[36568], Fresh[36567], Fresh[36566], Fresh[36565], Fresh[36564], Fresh[36563], Fresh[36562], Fresh[36561], Fresh[36560], Fresh[36559], Fresh[36558], Fresh[36557], Fresh[36556], Fresh[36555], Fresh[36554], Fresh[36553], Fresh[36552], Fresh[36551], Fresh[36550], Fresh[36549], Fresh[36548], Fresh[36547], Fresh[36546], Fresh[36545], Fresh[36544], Fresh[36543], Fresh[36542], Fresh[36541], Fresh[36540], Fresh[36539], Fresh[36538], Fresh[36537], Fresh[36536], Fresh[36535], Fresh[36534], Fresh[36533], Fresh[36532], Fresh[36531], Fresh[36530], Fresh[36529], Fresh[36528], Fresh[36527], Fresh[36526], Fresh[36525], Fresh[36524], Fresh[36523], Fresh[36522], Fresh[36521], Fresh[36520], Fresh[36519], Fresh[36518], Fresh[36517], Fresh[36516], Fresh[36515], Fresh[36514], Fresh[36513], Fresh[36512], Fresh[36511], Fresh[36510], Fresh[36509], Fresh[36508], Fresh[36507], Fresh[36506], Fresh[36505], Fresh[36504], Fresh[36503], Fresh[36502], Fresh[36501], Fresh[36500], Fresh[36499], Fresh[36498], Fresh[36497], Fresh[36496], Fresh[36495], Fresh[36494], Fresh[36493], Fresh[36492], Fresh[36491], Fresh[36490], Fresh[36489], Fresh[36488], Fresh[36487], Fresh[36486], Fresh[36485], Fresh[36484], Fresh[36483], Fresh[36482], Fresh[36481], Fresh[36480], Fresh[36479], Fresh[36478], Fresh[36477], Fresh[36476], Fresh[36475], Fresh[36474], Fresh[36473], Fresh[36472], Fresh[36471], Fresh[36470], Fresh[36469], Fresh[36468], Fresh[36467], Fresh[36466], Fresh[36465], Fresh[36464], Fresh[36463], Fresh[36462], Fresh[36461], Fresh[36460], Fresh[36459], Fresh[36458], Fresh[36457], Fresh[36456], Fresh[36455], Fresh[36454], Fresh[36453], Fresh[36452], Fresh[36451], Fresh[36450], Fresh[36449], Fresh[36448], Fresh[36447], Fresh[36446], Fresh[36445], Fresh[36444], Fresh[36443], Fresh[36442], Fresh[36441], Fresh[36440], Fresh[36439], Fresh[36438], Fresh[36437], Fresh[36436], Fresh[36435], Fresh[36434], Fresh[36433], Fresh[36432], Fresh[36431], Fresh[36430], Fresh[36429], Fresh[36428], Fresh[36427], Fresh[36426], Fresh[36425], Fresh[36424], Fresh[36423], Fresh[36422], Fresh[36421], Fresh[36420], Fresh[36419], Fresh[36418], Fresh[36417], Fresh[36416], Fresh[36415], Fresh[36414], Fresh[36413], Fresh[36412], Fresh[36411], Fresh[36410], Fresh[36409], Fresh[36408], Fresh[36407], Fresh[36406], Fresh[36405], Fresh[36404], Fresh[36403], Fresh[36402], Fresh[36401], Fresh[36400], Fresh[36399], Fresh[36398], Fresh[36397], Fresh[36396], Fresh[36395], Fresh[36394], Fresh[36393], Fresh[36392], Fresh[36391], Fresh[36390], Fresh[36389], Fresh[36388], Fresh[36387], Fresh[36386], Fresh[36385], Fresh[36384], Fresh[36383], Fresh[36382], Fresh[36381], Fresh[36380], Fresh[36379], Fresh[36378], Fresh[36377], Fresh[36376], Fresh[36375], Fresh[36374], Fresh[36373], Fresh[36372], Fresh[36371], Fresh[36370], Fresh[36369], Fresh[36368], Fresh[36367], Fresh[36366], Fresh[36365], Fresh[36364], Fresh[36363], Fresh[36362], Fresh[36361], Fresh[36360], Fresh[36359], Fresh[36358], Fresh[36357], Fresh[36356], Fresh[36355], Fresh[36354], Fresh[36353], Fresh[36352], Fresh[36351], Fresh[36350], Fresh[36349], Fresh[36348], Fresh[36347], Fresh[36346], Fresh[36345], Fresh[36344], Fresh[36343], Fresh[36342], Fresh[36341], Fresh[36340], Fresh[36339], Fresh[36338], Fresh[36337], Fresh[36336], Fresh[36335], Fresh[36334], Fresh[36333], Fresh[36332], Fresh[36331], Fresh[36330], Fresh[36329], Fresh[36328], Fresh[36327], Fresh[36326], Fresh[36325], Fresh[36324], Fresh[36323], Fresh[36322], Fresh[36321], Fresh[36320], Fresh[36319], Fresh[36318], Fresh[36317], Fresh[36316], Fresh[36315], Fresh[36314], Fresh[36313], Fresh[36312], Fresh[36311], Fresh[36310], Fresh[36309], Fresh[36308], Fresh[36307], Fresh[36306], Fresh[36305], Fresh[36304], Fresh[36303], Fresh[36302], Fresh[36301], Fresh[36300], Fresh[36299], Fresh[36298], Fresh[36297], Fresh[36296], Fresh[36295], Fresh[36294], Fresh[36293], Fresh[36292], Fresh[36291], Fresh[36290], Fresh[36289], Fresh[36288], Fresh[36287], Fresh[36286], Fresh[36285], Fresh[36284], Fresh[36283], Fresh[36282], Fresh[36281], Fresh[36280], Fresh[36279], Fresh[36278], Fresh[36277], Fresh[36276], Fresh[36275], Fresh[36274], Fresh[36273], Fresh[36272], Fresh[36271], Fresh[36270], Fresh[36269], Fresh[36268], Fresh[36267], Fresh[36266], Fresh[36265], Fresh[36264], Fresh[36263], Fresh[36262], Fresh[36261], Fresh[36260], Fresh[36259], Fresh[36258], Fresh[36257], Fresh[36256], Fresh[36255], Fresh[36254], Fresh[36253], Fresh[36252], Fresh[36251], Fresh[36250], Fresh[36249], Fresh[36248], Fresh[36247], Fresh[36246], Fresh[36245], Fresh[36244], Fresh[36243], Fresh[36242], Fresh[36241], Fresh[36240], Fresh[36239], Fresh[36238], Fresh[36237], Fresh[36236], Fresh[36235], Fresh[36234], Fresh[36233], Fresh[36232], Fresh[36231], Fresh[36230], Fresh[36229], Fresh[36228], Fresh[36227], Fresh[36226], Fresh[36225], Fresh[36224], Fresh[36223], Fresh[36222], Fresh[36221], Fresh[36220], Fresh[36219], Fresh[36218], Fresh[36217], Fresh[36216], Fresh[36215], Fresh[36214], Fresh[36213], Fresh[36212], Fresh[36211], Fresh[36210], Fresh[36209], Fresh[36208], Fresh[36207], Fresh[36206], Fresh[36205], Fresh[36204], Fresh[36203], Fresh[36202], Fresh[36201], Fresh[36200], Fresh[36199], Fresh[36198], Fresh[36197], Fresh[36196], Fresh[36195], Fresh[36194], Fresh[36193], Fresh[36192], Fresh[36191], Fresh[36190], Fresh[36189], Fresh[36188], Fresh[36187], Fresh[36186], Fresh[36185], Fresh[36184], Fresh[36183], Fresh[36182], Fresh[36181], Fresh[36180], Fresh[36179], Fresh[36178], Fresh[36177], Fresh[36176], Fresh[36175], Fresh[36174], Fresh[36173], Fresh[36172], Fresh[36171], Fresh[36170], Fresh[36169], Fresh[36168], Fresh[36167], Fresh[36166], Fresh[36165], Fresh[36164], Fresh[36163], Fresh[36162], Fresh[36161], Fresh[36160], Fresh[36159], Fresh[36158], Fresh[36157], Fresh[36156], Fresh[36155], Fresh[36154], Fresh[36153], Fresh[36152], Fresh[36151], Fresh[36150], Fresh[36149], Fresh[36148], Fresh[36147], Fresh[36146], Fresh[36145], Fresh[36144], Fresh[36143], Fresh[36142], Fresh[36141], Fresh[36140], Fresh[36139], Fresh[36138], Fresh[36137], Fresh[36136], Fresh[36135], Fresh[36134], Fresh[36133], Fresh[36132], Fresh[36131], Fresh[36130], Fresh[36129], Fresh[36128], Fresh[36127], Fresh[36126], Fresh[36125], Fresh[36124], Fresh[36123], Fresh[36122], Fresh[36121], Fresh[36120], Fresh[36119], Fresh[36118], Fresh[36117], Fresh[36116], Fresh[36115], Fresh[36114], Fresh[36113], Fresh[36112], Fresh[36111], Fresh[36110], Fresh[36109], Fresh[36108], Fresh[36107], Fresh[36106], Fresh[36105], Fresh[36104], Fresh[36103], Fresh[36102], Fresh[36101], Fresh[36100], Fresh[36099], Fresh[36098], Fresh[36097], Fresh[36096], Fresh[36095], Fresh[36094], Fresh[36093], Fresh[36092], Fresh[36091], Fresh[36090], Fresh[36089], Fresh[36088], Fresh[36087], Fresh[36086], Fresh[36085], Fresh[36084], Fresh[36083], Fresh[36082], Fresh[36081], Fresh[36080], Fresh[36079], Fresh[36078], Fresh[36077], Fresh[36076], Fresh[36075], Fresh[36074], Fresh[36073], Fresh[36072], Fresh[36071], Fresh[36070], Fresh[36069], Fresh[36068], Fresh[36067], Fresh[36066], Fresh[36065], Fresh[36064], Fresh[36063], Fresh[36062], Fresh[36061], Fresh[36060], Fresh[36059], Fresh[36058], Fresh[36057], Fresh[36056], Fresh[36055], Fresh[36054], Fresh[36053], Fresh[36052], Fresh[36051], Fresh[36050], Fresh[36049], Fresh[36048], Fresh[36047], Fresh[36046], Fresh[36045], Fresh[36044], Fresh[36043], Fresh[36042], Fresh[36041], Fresh[36040], Fresh[36039], Fresh[36038], Fresh[36037], Fresh[36036], Fresh[36035], Fresh[36034], Fresh[36033], Fresh[36032], Fresh[36031], Fresh[36030], Fresh[36029], Fresh[36028], Fresh[36027], Fresh[36026], Fresh[36025], Fresh[36024], Fresh[36023], Fresh[36022], Fresh[36021], Fresh[36020], Fresh[36019], Fresh[36018], Fresh[36017], Fresh[36016], Fresh[36015], Fresh[36014], Fresh[36013], Fresh[36012], Fresh[36011], Fresh[36010], Fresh[36009], Fresh[36008], Fresh[36007], Fresh[36006], Fresh[36005], Fresh[36004], Fresh[36003], Fresh[36002], Fresh[36001], Fresh[36000], Fresh[35999], Fresh[35998], Fresh[35997], Fresh[35996], Fresh[35995], Fresh[35994], Fresh[35993], Fresh[35992], Fresh[35991], Fresh[35990], Fresh[35989], Fresh[35988], Fresh[35987], Fresh[35986], Fresh[35985], Fresh[35984], Fresh[35983], Fresh[35982], Fresh[35981], Fresh[35980], Fresh[35979], Fresh[35978], Fresh[35977], Fresh[35976], Fresh[35975], Fresh[35974], Fresh[35973], Fresh[35972], Fresh[35971], Fresh[35970], Fresh[35969], Fresh[35968], Fresh[35967], Fresh[35966], Fresh[35965], Fresh[35964], Fresh[35963], Fresh[35962], Fresh[35961], Fresh[35960], Fresh[35959], Fresh[35958], Fresh[35957], Fresh[35956], Fresh[35955], Fresh[35954], Fresh[35953], Fresh[35952], Fresh[35951], Fresh[35950], Fresh[35949], Fresh[35948], Fresh[35947], Fresh[35946], Fresh[35945], Fresh[35944], Fresh[35943], Fresh[35942], Fresh[35941], Fresh[35940], Fresh[35939], Fresh[35938], Fresh[35937], Fresh[35936], Fresh[35935], Fresh[35934], Fresh[35933], Fresh[35932], Fresh[35931], Fresh[35930], Fresh[35929], Fresh[35928], Fresh[35927], Fresh[35926], Fresh[35925], Fresh[35924], Fresh[35923], Fresh[35922], Fresh[35921], Fresh[35920], Fresh[35919], Fresh[35918], Fresh[35917], Fresh[35916], Fresh[35915], Fresh[35914], Fresh[35913], Fresh[35912], Fresh[35911], Fresh[35910], Fresh[35909], Fresh[35908], Fresh[35907], Fresh[35906], Fresh[35905], Fresh[35904], Fresh[35903], Fresh[35902], Fresh[35901], Fresh[35900], Fresh[35899], Fresh[35898], Fresh[35897], Fresh[35896], Fresh[35895], Fresh[35894], Fresh[35893], Fresh[35892], Fresh[35891], Fresh[35890], Fresh[35889], Fresh[35888], Fresh[35887], Fresh[35886], Fresh[35885], Fresh[35884], Fresh[35883], Fresh[35882], Fresh[35881], Fresh[35880], Fresh[35879], Fresh[35878], Fresh[35877], Fresh[35876], Fresh[35875], Fresh[35874], Fresh[35873], Fresh[35872], Fresh[35871], Fresh[35870], Fresh[35869], Fresh[35868], Fresh[35867], Fresh[35866], Fresh[35865], Fresh[35864], Fresh[35863], Fresh[35862], Fresh[35861], Fresh[35860], Fresh[35859], Fresh[35858], Fresh[35857], Fresh[35856], Fresh[35855], Fresh[35854], Fresh[35853], Fresh[35852], Fresh[35851], Fresh[35850], Fresh[35849], Fresh[35848], Fresh[35847], Fresh[35846], Fresh[35845], Fresh[35844], Fresh[35843], Fresh[35842], Fresh[35841], Fresh[35840], Fresh[35839], Fresh[35838], Fresh[35837], Fresh[35836], Fresh[35835], Fresh[35834], Fresh[35833], Fresh[35832], Fresh[35831], Fresh[35830], Fresh[35829], Fresh[35828], Fresh[35827], Fresh[35826], Fresh[35825], Fresh[35824], Fresh[35823], Fresh[35822], Fresh[35821], Fresh[35820], Fresh[35819], Fresh[35818], Fresh[35817], Fresh[35816], Fresh[35815], Fresh[35814], Fresh[35813], Fresh[35812], Fresh[35811], Fresh[35810], Fresh[35809], Fresh[35808], Fresh[35807], Fresh[35806], Fresh[35805], Fresh[35804], Fresh[35803], Fresh[35802], Fresh[35801], Fresh[35800], Fresh[35799], Fresh[35798], Fresh[35797], Fresh[35796], Fresh[35795], Fresh[35794], Fresh[35793], Fresh[35792], Fresh[35791], Fresh[35790], Fresh[35789], Fresh[35788], Fresh[35787], Fresh[35786], Fresh[35785], Fresh[35784], Fresh[35783], Fresh[35782], Fresh[35781], Fresh[35780], Fresh[35779], Fresh[35778], Fresh[35777], Fresh[35776], Fresh[35775], Fresh[35774], Fresh[35773], Fresh[35772], Fresh[35771], Fresh[35770], Fresh[35769], Fresh[35768], Fresh[35767], Fresh[35766], Fresh[35765], Fresh[35764], Fresh[35763], Fresh[35762], Fresh[35761], Fresh[35760], Fresh[35759], Fresh[35758], Fresh[35757], Fresh[35756], Fresh[35755], Fresh[35754], Fresh[35753], Fresh[35752], Fresh[35751], Fresh[35750], Fresh[35749], Fresh[35748], Fresh[35747], Fresh[35746], Fresh[35745], Fresh[35744], Fresh[35743], Fresh[35742], Fresh[35741], Fresh[35740], Fresh[35739], Fresh[35738], Fresh[35737], Fresh[35736], Fresh[35735], Fresh[35734], Fresh[35733], Fresh[35732], Fresh[35731], Fresh[35730], Fresh[35729], Fresh[35728], Fresh[35727], Fresh[35726], Fresh[35725], Fresh[35724], Fresh[35723], Fresh[35722], Fresh[35721], Fresh[35720], Fresh[35719], Fresh[35718], Fresh[35717], Fresh[35716], Fresh[35715], Fresh[35714], Fresh[35713], Fresh[35712], Fresh[35711], Fresh[35710], Fresh[35709], Fresh[35708], Fresh[35707], Fresh[35706], Fresh[35705], Fresh[35704], Fresh[35703], Fresh[35702], Fresh[35701], Fresh[35700], Fresh[35699], Fresh[35698], Fresh[35697], Fresh[35696], Fresh[35695], Fresh[35694], Fresh[35693], Fresh[35692], Fresh[35691], Fresh[35690], Fresh[35689], Fresh[35688], Fresh[35687], Fresh[35686], Fresh[35685], Fresh[35684], Fresh[35683], Fresh[35682], Fresh[35681], Fresh[35680], Fresh[35679], Fresh[35678], Fresh[35677], Fresh[35676], Fresh[35675], Fresh[35674], Fresh[35673], Fresh[35672], Fresh[35671], Fresh[35670], Fresh[35669], Fresh[35668], Fresh[35667], Fresh[35666], Fresh[35665], Fresh[35664], Fresh[35663], Fresh[35662], Fresh[35661], Fresh[35660], Fresh[35659], Fresh[35658], Fresh[35657], Fresh[35656], Fresh[35655], Fresh[35654], Fresh[35653], Fresh[35652], Fresh[35651], Fresh[35650], Fresh[35649], Fresh[35648], Fresh[35647], Fresh[35646], Fresh[35645], Fresh[35644], Fresh[35643], Fresh[35642], Fresh[35641], Fresh[35640], Fresh[35639], Fresh[35638], Fresh[35637], Fresh[35636], Fresh[35635], Fresh[35634], Fresh[35633], Fresh[35632], Fresh[35631], Fresh[35630], Fresh[35629], Fresh[35628], Fresh[35627], Fresh[35626], Fresh[35625], Fresh[35624], Fresh[35623], Fresh[35622], Fresh[35621], Fresh[35620], Fresh[35619], Fresh[35618], Fresh[35617], Fresh[35616], Fresh[35615], Fresh[35614], Fresh[35613], Fresh[35612], Fresh[35611], Fresh[35610], Fresh[35609], Fresh[35608], Fresh[35607], Fresh[35606], Fresh[35605], Fresh[35604], Fresh[35603], Fresh[35602], Fresh[35601], Fresh[35600], Fresh[35599], Fresh[35598], Fresh[35597], Fresh[35596], Fresh[35595], Fresh[35594], Fresh[35593], Fresh[35592], Fresh[35591], Fresh[35590], Fresh[35589], Fresh[35588], Fresh[35587], Fresh[35586], Fresh[35585], Fresh[35584], Fresh[35583], Fresh[35582], Fresh[35581], Fresh[35580], Fresh[35579], Fresh[35578], Fresh[35577], Fresh[35576], Fresh[35575], Fresh[35574], Fresh[35573], Fresh[35572], Fresh[35571], Fresh[35570], Fresh[35569], Fresh[35568], Fresh[35567], Fresh[35566], Fresh[35565], Fresh[35564], Fresh[35563], Fresh[35562], Fresh[35561], Fresh[35560], Fresh[35559], Fresh[35558], Fresh[35557], Fresh[35556], Fresh[35555], Fresh[35554], Fresh[35553], Fresh[35552], Fresh[35551], Fresh[35550], Fresh[35549], Fresh[35548], Fresh[35547], Fresh[35546], Fresh[35545], Fresh[35544], Fresh[35543], Fresh[35542], Fresh[35541], Fresh[35540], Fresh[35539], Fresh[35538], Fresh[35537], Fresh[35536], Fresh[35535], Fresh[35534], Fresh[35533], Fresh[35532], Fresh[35531], Fresh[35530], Fresh[35529], Fresh[35528], Fresh[35527], Fresh[35526], Fresh[35525], Fresh[35524], Fresh[35523], Fresh[35522], Fresh[35521], Fresh[35520], Fresh[35519], Fresh[35518], Fresh[35517], Fresh[35516], Fresh[35515], Fresh[35514], Fresh[35513], Fresh[35512], Fresh[35511], Fresh[35510], Fresh[35509], Fresh[35508], Fresh[35507], Fresh[35506], Fresh[35505], Fresh[35504], Fresh[35503], Fresh[35502], Fresh[35501], Fresh[35500], Fresh[35499], Fresh[35498], Fresh[35497], Fresh[35496], Fresh[35495], Fresh[35494], Fresh[35493], Fresh[35492], Fresh[35491], Fresh[35490], Fresh[35489], Fresh[35488], Fresh[35487], Fresh[35486], Fresh[35485], Fresh[35484], Fresh[35483], Fresh[35482], Fresh[35481], Fresh[35480], Fresh[35479], Fresh[35478], Fresh[35477], Fresh[35476], Fresh[35475], Fresh[35474], Fresh[35473], Fresh[35472], Fresh[35471], Fresh[35470], Fresh[35469], Fresh[35468], Fresh[35467], Fresh[35466], Fresh[35465], Fresh[35464], Fresh[35463], Fresh[35462], Fresh[35461], Fresh[35460], Fresh[35459], Fresh[35458], Fresh[35457], Fresh[35456], Fresh[35455], Fresh[35454], Fresh[35453], Fresh[35452], Fresh[35451], Fresh[35450], Fresh[35449], Fresh[35448], Fresh[35447], Fresh[35446], Fresh[35445], Fresh[35444], Fresh[35443], Fresh[35442], Fresh[35441], Fresh[35440], Fresh[35439], Fresh[35438], Fresh[35437], Fresh[35436], Fresh[35435], Fresh[35434], Fresh[35433], Fresh[35432], Fresh[35431], Fresh[35430], Fresh[35429], Fresh[35428], Fresh[35427], Fresh[35426], Fresh[35425], Fresh[35424], Fresh[35423], Fresh[35422], Fresh[35421], Fresh[35420], Fresh[35419], Fresh[35418], Fresh[35417], Fresh[35416], Fresh[35415], Fresh[35414], Fresh[35413], Fresh[35412], Fresh[35411], Fresh[35410], Fresh[35409], Fresh[35408], Fresh[35407], Fresh[35406], Fresh[35405], Fresh[35404], Fresh[35403], Fresh[35402], Fresh[35401], Fresh[35400], Fresh[35399], Fresh[35398], Fresh[35397], Fresh[35396], Fresh[35395], Fresh[35394], Fresh[35393], Fresh[35392], Fresh[35391], Fresh[35390], Fresh[35389], Fresh[35388], Fresh[35387], Fresh[35386], Fresh[35385], Fresh[35384], Fresh[35383], Fresh[35382], Fresh[35381], Fresh[35380], Fresh[35379], Fresh[35378], Fresh[35377], Fresh[35376], Fresh[35375], Fresh[35374], Fresh[35373], Fresh[35372], Fresh[35371], Fresh[35370], Fresh[35369], Fresh[35368], Fresh[35367], Fresh[35366], Fresh[35365], Fresh[35364], Fresh[35363], Fresh[35362], Fresh[35361], Fresh[35360], Fresh[35359], Fresh[35358], Fresh[35357], Fresh[35356], Fresh[35355], Fresh[35354], Fresh[35353], Fresh[35352], Fresh[35351], Fresh[35350], Fresh[35349], Fresh[35348], Fresh[35347], Fresh[35346], Fresh[35345], Fresh[35344], Fresh[35343], Fresh[35342], Fresh[35341], Fresh[35340], Fresh[35339], Fresh[35338], Fresh[35337], Fresh[35336], Fresh[35335], Fresh[35334], Fresh[35333], Fresh[35332], Fresh[35331], Fresh[35330], Fresh[35329], Fresh[35328], Fresh[35327], Fresh[35326], Fresh[35325], Fresh[35324], Fresh[35323], Fresh[35322], Fresh[35321], Fresh[35320], Fresh[35319], Fresh[35318], Fresh[35317], Fresh[35316], Fresh[35315], Fresh[35314], Fresh[35313], Fresh[35312], Fresh[35311], Fresh[35310], Fresh[35309], Fresh[35308], Fresh[35307], Fresh[35306], Fresh[35305], Fresh[35304], Fresh[35303], Fresh[35302], Fresh[35301], Fresh[35300], Fresh[35299], Fresh[35298], Fresh[35297], Fresh[35296], Fresh[35295], Fresh[35294], Fresh[35293], Fresh[35292], Fresh[35291], Fresh[35290], Fresh[35289], Fresh[35288], Fresh[35287], Fresh[35286], Fresh[35285], Fresh[35284], Fresh[35283], Fresh[35282], Fresh[35281], Fresh[35280], Fresh[35279], Fresh[35278], Fresh[35277], Fresh[35276], Fresh[35275], Fresh[35274], Fresh[35273], Fresh[35272], Fresh[35271], Fresh[35270], Fresh[35269], Fresh[35268], Fresh[35267], Fresh[35266], Fresh[35265], Fresh[35264], Fresh[35263], Fresh[35262], Fresh[35261], Fresh[35260], Fresh[35259], Fresh[35258], Fresh[35257], Fresh[35256], Fresh[35255], Fresh[35254], Fresh[35253], Fresh[35252], Fresh[35251], Fresh[35250], Fresh[35249], Fresh[35248], Fresh[35247], Fresh[35246], Fresh[35245], Fresh[35244], Fresh[35243], Fresh[35242], Fresh[35241], Fresh[35240], Fresh[35239], Fresh[35238], Fresh[35237], Fresh[35236], Fresh[35235], Fresh[35234], Fresh[35233], Fresh[35232], Fresh[35231], Fresh[35230], Fresh[35229], Fresh[35228], Fresh[35227], Fresh[35226], Fresh[35225], Fresh[35224], Fresh[35223], Fresh[35222], Fresh[35221], Fresh[35220], Fresh[35219], Fresh[35218], Fresh[35217], Fresh[35216], Fresh[35215], Fresh[35214], Fresh[35213], Fresh[35212], Fresh[35211], Fresh[35210], Fresh[35209], Fresh[35208], Fresh[35207], Fresh[35206], Fresh[35205], Fresh[35204], Fresh[35203], Fresh[35202], Fresh[35201], Fresh[35200], Fresh[35199], Fresh[35198], Fresh[35197], Fresh[35196], Fresh[35195], Fresh[35194], Fresh[35193], Fresh[35192], Fresh[35191], Fresh[35190], Fresh[35189], Fresh[35188], Fresh[35187], Fresh[35186], Fresh[35185], Fresh[35184], Fresh[35183], Fresh[35182], Fresh[35181], Fresh[35180], Fresh[35179], Fresh[35178], Fresh[35177], Fresh[35176], Fresh[35175], Fresh[35174], Fresh[35173], Fresh[35172], Fresh[35171], Fresh[35170], Fresh[35169], Fresh[35168], Fresh[35167], Fresh[35166], Fresh[35165], Fresh[35164], Fresh[35163], Fresh[35162], Fresh[35161], Fresh[35160], Fresh[35159], Fresh[35158], Fresh[35157], Fresh[35156], Fresh[35155], Fresh[35154], Fresh[35153], Fresh[35152], Fresh[35151], Fresh[35150], Fresh[35149], Fresh[35148], Fresh[35147], Fresh[35146], Fresh[35145], Fresh[35144], Fresh[35143], Fresh[35142], Fresh[35141], Fresh[35140], Fresh[35139], Fresh[35138], Fresh[35137], Fresh[35136], Fresh[35135], Fresh[35134], Fresh[35133], Fresh[35132], Fresh[35131], Fresh[35130], Fresh[35129], Fresh[35128], Fresh[35127], Fresh[35126], Fresh[35125], Fresh[35124], Fresh[35123], Fresh[35122], Fresh[35121], Fresh[35120], Fresh[35119], Fresh[35118], Fresh[35117], Fresh[35116], Fresh[35115], Fresh[35114], Fresh[35113], Fresh[35112], Fresh[35111], Fresh[35110], Fresh[35109], Fresh[35108], Fresh[35107], Fresh[35106], Fresh[35105], Fresh[35104], Fresh[35103], Fresh[35102], Fresh[35101], Fresh[35100], Fresh[35099], Fresh[35098], Fresh[35097], Fresh[35096], Fresh[35095], Fresh[35094], Fresh[35093], Fresh[35092], Fresh[35091], Fresh[35090], Fresh[35089], Fresh[35088], Fresh[35087], Fresh[35086], Fresh[35085], Fresh[35084], Fresh[35083], Fresh[35082], Fresh[35081], Fresh[35080], Fresh[35079], Fresh[35078], Fresh[35077], Fresh[35076], Fresh[35075], Fresh[35074], Fresh[35073], Fresh[35072], Fresh[35071], Fresh[35070], Fresh[35069], Fresh[35068], Fresh[35067], Fresh[35066], Fresh[35065], Fresh[35064], Fresh[35063], Fresh[35062], Fresh[35061], Fresh[35060], Fresh[35059], Fresh[35058], Fresh[35057], Fresh[35056], Fresh[35055], Fresh[35054], Fresh[35053], Fresh[35052], Fresh[35051], Fresh[35050], Fresh[35049], Fresh[35048], Fresh[35047], Fresh[35046], Fresh[35045], Fresh[35044], Fresh[35043], Fresh[35042], Fresh[35041], Fresh[35040], Fresh[35039], Fresh[35038], Fresh[35037], Fresh[35036], Fresh[35035], Fresh[35034], Fresh[35033], Fresh[35032], Fresh[35031], Fresh[35030], Fresh[35029], Fresh[35028], Fresh[35027], Fresh[35026], Fresh[35025], Fresh[35024], Fresh[35023], Fresh[35022], Fresh[35021], Fresh[35020], Fresh[35019], Fresh[35018], Fresh[35017], Fresh[35016], Fresh[35015], Fresh[35014], Fresh[35013], Fresh[35012], Fresh[35011], Fresh[35010], Fresh[35009], Fresh[35008], Fresh[35007], Fresh[35006], Fresh[35005], Fresh[35004], Fresh[35003], Fresh[35002], Fresh[35001], Fresh[35000], Fresh[34999], Fresh[34998], Fresh[34997], Fresh[34996], Fresh[34995], Fresh[34994], Fresh[34993], Fresh[34992], Fresh[34991], Fresh[34990], Fresh[34989], Fresh[34988], Fresh[34987], Fresh[34986], Fresh[34985], Fresh[34984], Fresh[34983], Fresh[34982], Fresh[34981], Fresh[34980], Fresh[34979], Fresh[34978], Fresh[34977], Fresh[34976], Fresh[34975], Fresh[34974], Fresh[34973], Fresh[34972], Fresh[34971], Fresh[34970], Fresh[34969], Fresh[34968], Fresh[34967], Fresh[34966], Fresh[34965], Fresh[34964], Fresh[34963], Fresh[34962], Fresh[34961], Fresh[34960], Fresh[34959], Fresh[34958], Fresh[34957], Fresh[34956], Fresh[34955], Fresh[34954], Fresh[34953], Fresh[34952], Fresh[34951], Fresh[34950], Fresh[34949], Fresh[34948], Fresh[34947], Fresh[34946], Fresh[34945], Fresh[34944], Fresh[34943], Fresh[34942], Fresh[34941], Fresh[34940], Fresh[34939], Fresh[34938], Fresh[34937], Fresh[34936], Fresh[34935], Fresh[34934], Fresh[34933], Fresh[34932], Fresh[34931], Fresh[34930], Fresh[34929], Fresh[34928], Fresh[34927], Fresh[34926], Fresh[34925], Fresh[34924], Fresh[34923], Fresh[34922], Fresh[34921], Fresh[34920], Fresh[34919], Fresh[34918], Fresh[34917], Fresh[34916], Fresh[34915], Fresh[34914], Fresh[34913], Fresh[34912], Fresh[34911], Fresh[34910], Fresh[34909], Fresh[34908], Fresh[34907], Fresh[34906], Fresh[34905], Fresh[34904], Fresh[34903], Fresh[34902], Fresh[34901], Fresh[34900], Fresh[34899], Fresh[34898], Fresh[34897], Fresh[34896], Fresh[34895], Fresh[34894], Fresh[34893], Fresh[34892], Fresh[34891], Fresh[34890], Fresh[34889], Fresh[34888], Fresh[34887], Fresh[34886], Fresh[34885], Fresh[34884], Fresh[34883], Fresh[34882], Fresh[34881], Fresh[34880], Fresh[34879], Fresh[34878], Fresh[34877], Fresh[34876], Fresh[34875], Fresh[34874], Fresh[34873], Fresh[34872], Fresh[34871], Fresh[34870], Fresh[34869], Fresh[34868], Fresh[34867], Fresh[34866], Fresh[34865], Fresh[34864], Fresh[34863], Fresh[34862], Fresh[34861], Fresh[34860], Fresh[34859], Fresh[34858], Fresh[34857], Fresh[34856], Fresh[34855], Fresh[34854], Fresh[34853], Fresh[34852], Fresh[34851], Fresh[34850], Fresh[34849], Fresh[34848], Fresh[34847], Fresh[34846], Fresh[34845], Fresh[34844], Fresh[34843], Fresh[34842], Fresh[34841], Fresh[34840], Fresh[34839], Fresh[34838], Fresh[34837], Fresh[34836], Fresh[34835], Fresh[34834], Fresh[34833], Fresh[34832], Fresh[34831], Fresh[34830], Fresh[34829], Fresh[34828], Fresh[34827], Fresh[34826], Fresh[34825], Fresh[34824], Fresh[34823], Fresh[34822], Fresh[34821], Fresh[34820], Fresh[34819], Fresh[34818], Fresh[34817], Fresh[34816], Fresh[34815], Fresh[34814], Fresh[34813], Fresh[34812], Fresh[34811], Fresh[34810], Fresh[34809], Fresh[34808], Fresh[34807], Fresh[34806], Fresh[34805], Fresh[34804], Fresh[34803], Fresh[34802], Fresh[34801], Fresh[34800], Fresh[34799], Fresh[34798], Fresh[34797], Fresh[34796], Fresh[34795], Fresh[34794], Fresh[34793], Fresh[34792], Fresh[34791], Fresh[34790], Fresh[34789], Fresh[34788], Fresh[34787], Fresh[34786], Fresh[34785], Fresh[34784], Fresh[34783], Fresh[34782], Fresh[34781], Fresh[34780], Fresh[34779], Fresh[34778], Fresh[34777], Fresh[34776], Fresh[34775], Fresh[34774], Fresh[34773], Fresh[34772], Fresh[34771], Fresh[34770], Fresh[34769], Fresh[34768], Fresh[34767], Fresh[34766], Fresh[34765], Fresh[34764], Fresh[34763], Fresh[34762], Fresh[34761], Fresh[34760], Fresh[34759], Fresh[34758], Fresh[34757], Fresh[34756], Fresh[34755], Fresh[34754], Fresh[34753], Fresh[34752], Fresh[34751], Fresh[34750], Fresh[34749], Fresh[34748], Fresh[34747], Fresh[34746], Fresh[34745], Fresh[34744], Fresh[34743], Fresh[34742], Fresh[34741], Fresh[34740], Fresh[34739], Fresh[34738], Fresh[34737], Fresh[34736], Fresh[34735], Fresh[34734], Fresh[34733], Fresh[34732], Fresh[34731], Fresh[34730], Fresh[34729], Fresh[34728], Fresh[34727], Fresh[34726], Fresh[34725], Fresh[34724], Fresh[34723], Fresh[34722], Fresh[34721], Fresh[34720], Fresh[34719], Fresh[34718], Fresh[34717], Fresh[34716], Fresh[34715], Fresh[34714], Fresh[34713], Fresh[34712], Fresh[34711], Fresh[34710], Fresh[34709], Fresh[34708], Fresh[34707], Fresh[34706], Fresh[34705], Fresh[34704], Fresh[34703], Fresh[34702], Fresh[34701], Fresh[34700], Fresh[34699], Fresh[34698], Fresh[34697], Fresh[34696], Fresh[34695], Fresh[34694], Fresh[34693], Fresh[34692], Fresh[34691], Fresh[34690], Fresh[34689], Fresh[34688], Fresh[34687], Fresh[34686], Fresh[34685], Fresh[34684], Fresh[34683], Fresh[34682], Fresh[34681], Fresh[34680], Fresh[34679], Fresh[34678], Fresh[34677], Fresh[34676], Fresh[34675], Fresh[34674], Fresh[34673], Fresh[34672], Fresh[34671], Fresh[34670], Fresh[34669], Fresh[34668], Fresh[34667], Fresh[34666], Fresh[34665], Fresh[34664], Fresh[34663], Fresh[34662], Fresh[34661], Fresh[34660], Fresh[34659], Fresh[34658], Fresh[34657], Fresh[34656], Fresh[34655], Fresh[34654], Fresh[34653], Fresh[34652], Fresh[34651], Fresh[34650], Fresh[34649], Fresh[34648], Fresh[34647], Fresh[34646], Fresh[34645], Fresh[34644], Fresh[34643], Fresh[34642], Fresh[34641], Fresh[34640], Fresh[34639], Fresh[34638], Fresh[34637], Fresh[34636], Fresh[34635], Fresh[34634], Fresh[34633], Fresh[34632], Fresh[34631], Fresh[34630], Fresh[34629], Fresh[34628], Fresh[34627], Fresh[34626], Fresh[34625], Fresh[34624], Fresh[34623], Fresh[34622], Fresh[34621], Fresh[34620], Fresh[34619], Fresh[34618], Fresh[34617], Fresh[34616], Fresh[34615], Fresh[34614], Fresh[34613], Fresh[34612], Fresh[34611], Fresh[34610], Fresh[34609], Fresh[34608], Fresh[34607], Fresh[34606], Fresh[34605], Fresh[34604], Fresh[34603], Fresh[34602], Fresh[34601], Fresh[34600], Fresh[34599], Fresh[34598], Fresh[34597], Fresh[34596], Fresh[34595], Fresh[34594], Fresh[34593], Fresh[34592], Fresh[34591], Fresh[34590], Fresh[34589], Fresh[34588], Fresh[34587], Fresh[34586], Fresh[34585], Fresh[34584], Fresh[34583], Fresh[34582], Fresh[34581], Fresh[34580], Fresh[34579], Fresh[34578], Fresh[34577], Fresh[34576], Fresh[34575], Fresh[34574], Fresh[34573], Fresh[34572], Fresh[34571], Fresh[34570], Fresh[34569], Fresh[34568], Fresh[34567], Fresh[34566], Fresh[34565], Fresh[34564], Fresh[34563], Fresh[34562], Fresh[34561], Fresh[34560], Fresh[34559], Fresh[34558], Fresh[34557], Fresh[34556], Fresh[34555], Fresh[34554], Fresh[34553], Fresh[34552], Fresh[34551], Fresh[34550], Fresh[34549], Fresh[34548], Fresh[34547], Fresh[34546], Fresh[34545], Fresh[34544], Fresh[34543], Fresh[34542], Fresh[34541], Fresh[34540], Fresh[34539], Fresh[34538], Fresh[34537], Fresh[34536], Fresh[34535], Fresh[34534], Fresh[34533], Fresh[34532], Fresh[34531], Fresh[34530], Fresh[34529], Fresh[34528], Fresh[34527], Fresh[34526], Fresh[34525], Fresh[34524], Fresh[34523], Fresh[34522], Fresh[34521], Fresh[34520], Fresh[34519], Fresh[34518], Fresh[34517], Fresh[34516], Fresh[34515], Fresh[34514], Fresh[34513], Fresh[34512], Fresh[34511], Fresh[34510], Fresh[34509], Fresh[34508], Fresh[34507], Fresh[34506], Fresh[34505], Fresh[34504], Fresh[34503], Fresh[34502], Fresh[34501], Fresh[34500], Fresh[34499], Fresh[34498], Fresh[34497], Fresh[34496], Fresh[34495], Fresh[34494], Fresh[34493], Fresh[34492], Fresh[34491], Fresh[34490], Fresh[34489], Fresh[34488], Fresh[34487], Fresh[34486], Fresh[34485], Fresh[34484], Fresh[34483], Fresh[34482], Fresh[34481], Fresh[34480], Fresh[34479], Fresh[34478], Fresh[34477], Fresh[34476], Fresh[34475], Fresh[34474], Fresh[34473], Fresh[34472], Fresh[34471], Fresh[34470], Fresh[34469], Fresh[34468], Fresh[34467], Fresh[34466], Fresh[34465], Fresh[34464], Fresh[34463], Fresh[34462], Fresh[34461], Fresh[34460], Fresh[34459], Fresh[34458], Fresh[34457], Fresh[34456], Fresh[34455], Fresh[34454], Fresh[34453], Fresh[34452], Fresh[34451], Fresh[34450], Fresh[34449], Fresh[34448], Fresh[34447], Fresh[34446], Fresh[34445], Fresh[34444], Fresh[34443], Fresh[34442], Fresh[34441], Fresh[34440], Fresh[34439], Fresh[34438], Fresh[34437], Fresh[34436], Fresh[34435], Fresh[34434], Fresh[34433], Fresh[34432], Fresh[34431], Fresh[34430], Fresh[34429], Fresh[34428], Fresh[34427], Fresh[34426], Fresh[34425], Fresh[34424], Fresh[34423], Fresh[34422], Fresh[34421], Fresh[34420], Fresh[34419], Fresh[34418], Fresh[34417], Fresh[34416], Fresh[34415], Fresh[34414], Fresh[34413], Fresh[34412], Fresh[34411], Fresh[34410], Fresh[34409], Fresh[34408], Fresh[34407], Fresh[34406], Fresh[34405], Fresh[34404], Fresh[34403], Fresh[34402], Fresh[34401], Fresh[34400], Fresh[34399], Fresh[34398], Fresh[34397], Fresh[34396], Fresh[34395], Fresh[34394], Fresh[34393], Fresh[34392], Fresh[34391], Fresh[34390], Fresh[34389], Fresh[34388], Fresh[34387], Fresh[34386], Fresh[34385], Fresh[34384], Fresh[34383], Fresh[34382], Fresh[34381], Fresh[34380], Fresh[34379], Fresh[34378], Fresh[34377], Fresh[34376], Fresh[34375], Fresh[34374], Fresh[34373], Fresh[34372], Fresh[34371], Fresh[34370], Fresh[34369], Fresh[34368], Fresh[34367], Fresh[34366], Fresh[34365], Fresh[34364], Fresh[34363], Fresh[34362], Fresh[34361], Fresh[34360], Fresh[34359], Fresh[34358], Fresh[34357], Fresh[34356], Fresh[34355], Fresh[34354], Fresh[34353], Fresh[34352], Fresh[34351], Fresh[34350], Fresh[34349], Fresh[34348], Fresh[34347], Fresh[34346], Fresh[34345], Fresh[34344], Fresh[34343], Fresh[34342], Fresh[34341], Fresh[34340], Fresh[34339], Fresh[34338], Fresh[34337], Fresh[34336], Fresh[34335], Fresh[34334], Fresh[34333], Fresh[34332], Fresh[34331], Fresh[34330], Fresh[34329], Fresh[34328], Fresh[34327], Fresh[34326], Fresh[34325], Fresh[34324], Fresh[34323], Fresh[34322], Fresh[34321], Fresh[34320], Fresh[34319], Fresh[34318], Fresh[34317], Fresh[34316], Fresh[34315], Fresh[34314], Fresh[34313], Fresh[34312], Fresh[34311], Fresh[34310], Fresh[34309], Fresh[34308], Fresh[34307], Fresh[34306], Fresh[34305], Fresh[34304], Fresh[34303], Fresh[34302], Fresh[34301], Fresh[34300], Fresh[34299], Fresh[34298], Fresh[34297], Fresh[34296], Fresh[34295], Fresh[34294], Fresh[34293], Fresh[34292], Fresh[34291], Fresh[34290], Fresh[34289], Fresh[34288], Fresh[34287], Fresh[34286], Fresh[34285], Fresh[34284], Fresh[34283], Fresh[34282], Fresh[34281], Fresh[34280], Fresh[34279], Fresh[34278], Fresh[34277], Fresh[34276], Fresh[34275], Fresh[34274], Fresh[34273], Fresh[34272], Fresh[34271], Fresh[34270], Fresh[34269], Fresh[34268], Fresh[34267], Fresh[34266], Fresh[34265], Fresh[34264], Fresh[34263], Fresh[34262], Fresh[34261], Fresh[34260], Fresh[34259], Fresh[34258], Fresh[34257], Fresh[34256], Fresh[34255], Fresh[34254], Fresh[34253], Fresh[34252], Fresh[34251], Fresh[34250], Fresh[34249], Fresh[34248], Fresh[34247], Fresh[34246], Fresh[34245], Fresh[34244], Fresh[34243], Fresh[34242], Fresh[34241], Fresh[34240], Fresh[34239], Fresh[34238], Fresh[34237], Fresh[34236], Fresh[34235], Fresh[34234], Fresh[34233], Fresh[34232], Fresh[34231], Fresh[34230], Fresh[34229], Fresh[34228], Fresh[34227], Fresh[34226], Fresh[34225], Fresh[34224], Fresh[34223], Fresh[34222], Fresh[34221], Fresh[34220], Fresh[34219], Fresh[34218], Fresh[34217], Fresh[34216], Fresh[34215], Fresh[34214], Fresh[34213], Fresh[34212], Fresh[34211], Fresh[34210], Fresh[34209], Fresh[34208], Fresh[34207], Fresh[34206], Fresh[34205], Fresh[34204], Fresh[34203], Fresh[34202], Fresh[34201], Fresh[34200], Fresh[34199], Fresh[34198], Fresh[34197], Fresh[34196], Fresh[34195], Fresh[34194], Fresh[34193], Fresh[34192], Fresh[34191], Fresh[34190], Fresh[34189], Fresh[34188], Fresh[34187], Fresh[34186], Fresh[34185], Fresh[34184], Fresh[34183], Fresh[34182], Fresh[34181], Fresh[34180], Fresh[34179], Fresh[34178], Fresh[34177], Fresh[34176], Fresh[34175], Fresh[34174], Fresh[34173], Fresh[34172], Fresh[34171], Fresh[34170], Fresh[34169], Fresh[34168], Fresh[34167], Fresh[34166], Fresh[34165], Fresh[34164], Fresh[34163], Fresh[34162], Fresh[34161], Fresh[34160], Fresh[34159], Fresh[34158], Fresh[34157], Fresh[34156], Fresh[34155], Fresh[34154], Fresh[34153], Fresh[34152], Fresh[34151], Fresh[34150], Fresh[34149], Fresh[34148], Fresh[34147], Fresh[34146], Fresh[34145], Fresh[34144], Fresh[34143], Fresh[34142], Fresh[34141], Fresh[34140], Fresh[34139], Fresh[34138], Fresh[34137], Fresh[34136], Fresh[34135], Fresh[34134], Fresh[34133], Fresh[34132], Fresh[34131], Fresh[34130], Fresh[34129], Fresh[34128], Fresh[34127], Fresh[34126], Fresh[34125], Fresh[34124], Fresh[34123], Fresh[34122], Fresh[34121], Fresh[34120], Fresh[34119], Fresh[34118], Fresh[34117], Fresh[34116], Fresh[34115], Fresh[34114], Fresh[34113], Fresh[34112], Fresh[34111], Fresh[34110], Fresh[34109], Fresh[34108], Fresh[34107], Fresh[34106], Fresh[34105], Fresh[34104], Fresh[34103], Fresh[34102], Fresh[34101], Fresh[34100], Fresh[34099], Fresh[34098], Fresh[34097], Fresh[34096], Fresh[34095], Fresh[34094], Fresh[34093], Fresh[34092], Fresh[34091], Fresh[34090], Fresh[34089], Fresh[34088], Fresh[34087], Fresh[34086], Fresh[34085], Fresh[34084], Fresh[34083], Fresh[34082], Fresh[34081], Fresh[34080], Fresh[34079], Fresh[34078], Fresh[34077], Fresh[34076], Fresh[34075], Fresh[34074], Fresh[34073], Fresh[34072], Fresh[34071], Fresh[34070], Fresh[34069], Fresh[34068], Fresh[34067], Fresh[34066], Fresh[34065], Fresh[34064], Fresh[34063], Fresh[34062], Fresh[34061], Fresh[34060], Fresh[34059], Fresh[34058], Fresh[34057], Fresh[34056], Fresh[34055], Fresh[34054], Fresh[34053], Fresh[34052], Fresh[34051], Fresh[34050], Fresh[34049], Fresh[34048], Fresh[34047], Fresh[34046], Fresh[34045], Fresh[34044], Fresh[34043], Fresh[34042], Fresh[34041], Fresh[34040], Fresh[34039], Fresh[34038], Fresh[34037], Fresh[34036], Fresh[34035], Fresh[34034], Fresh[34033], Fresh[34032], Fresh[34031], Fresh[34030], Fresh[34029], Fresh[34028], Fresh[34027], Fresh[34026], Fresh[34025], Fresh[34024], Fresh[34023], Fresh[34022], Fresh[34021], Fresh[34020], Fresh[34019], Fresh[34018], Fresh[34017], Fresh[34016], Fresh[34015], Fresh[34014], Fresh[34013], Fresh[34012], Fresh[34011], Fresh[34010], Fresh[34009], Fresh[34008], Fresh[34007], Fresh[34006], Fresh[34005], Fresh[34004], Fresh[34003], Fresh[34002], Fresh[34001], Fresh[34000], Fresh[33999], Fresh[33998], Fresh[33997], Fresh[33996], Fresh[33995], Fresh[33994], Fresh[33993], Fresh[33992], Fresh[33991], Fresh[33990], Fresh[33989], Fresh[33988], Fresh[33987], Fresh[33986], Fresh[33985], Fresh[33984], Fresh[33983], Fresh[33982], Fresh[33981], Fresh[33980], Fresh[33979], Fresh[33978], Fresh[33977], Fresh[33976], Fresh[33975], Fresh[33974], Fresh[33973], Fresh[33972], Fresh[33971], Fresh[33970], Fresh[33969], Fresh[33968], Fresh[33967], Fresh[33966], Fresh[33965], Fresh[33964], Fresh[33963], Fresh[33962], Fresh[33961], Fresh[33960], Fresh[33959], Fresh[33958], Fresh[33957], Fresh[33956], Fresh[33955], Fresh[33954], Fresh[33953], Fresh[33952], Fresh[33951], Fresh[33950], Fresh[33949], Fresh[33948], Fresh[33947], Fresh[33946], Fresh[33945], Fresh[33944], Fresh[33943], Fresh[33942], Fresh[33941], Fresh[33940], Fresh[33939], Fresh[33938], Fresh[33937], Fresh[33936], Fresh[33935], Fresh[33934], Fresh[33933], Fresh[33932], Fresh[33931], Fresh[33930], Fresh[33929], Fresh[33928], Fresh[33927], Fresh[33926], Fresh[33925], Fresh[33924], Fresh[33923], Fresh[33922], Fresh[33921], Fresh[33920], Fresh[33919], Fresh[33918], Fresh[33917], Fresh[33916], Fresh[33915], Fresh[33914], Fresh[33913], Fresh[33912], Fresh[33911], Fresh[33910], Fresh[33909], Fresh[33908], Fresh[33907], Fresh[33906], Fresh[33905], Fresh[33904], Fresh[33903], Fresh[33902], Fresh[33901], Fresh[33900], Fresh[33899], Fresh[33898], Fresh[33897], Fresh[33896], Fresh[33895], Fresh[33894], Fresh[33893], Fresh[33892], Fresh[33891], Fresh[33890], Fresh[33889], Fresh[33888], Fresh[33887], Fresh[33886], Fresh[33885], Fresh[33884], Fresh[33883], Fresh[33882], Fresh[33881], Fresh[33880], Fresh[33879], Fresh[33878], Fresh[33877], Fresh[33876], Fresh[33875], Fresh[33874], Fresh[33873], Fresh[33872], Fresh[33871], Fresh[33870], Fresh[33869], Fresh[33868], Fresh[33867], Fresh[33866], Fresh[33865], Fresh[33864], Fresh[33863], Fresh[33862], Fresh[33861], Fresh[33860], Fresh[33859], Fresh[33858], Fresh[33857], Fresh[33856], Fresh[33855], Fresh[33854], Fresh[33853], Fresh[33852], Fresh[33851], Fresh[33850], Fresh[33849], Fresh[33848], Fresh[33847], Fresh[33846], Fresh[33845], Fresh[33844], Fresh[33843], Fresh[33842], Fresh[33841], Fresh[33840], Fresh[33839], Fresh[33838], Fresh[33837], Fresh[33836], Fresh[33835], Fresh[33834], Fresh[33833], Fresh[33832], Fresh[33831], Fresh[33830], Fresh[33829], Fresh[33828], Fresh[33827], Fresh[33826], Fresh[33825], Fresh[33824], Fresh[33823], Fresh[33822], Fresh[33821], Fresh[33820], Fresh[33819], Fresh[33818], Fresh[33817], Fresh[33816], Fresh[33815], Fresh[33814], Fresh[33813], Fresh[33812], Fresh[33811], Fresh[33810], Fresh[33809], Fresh[33808], Fresh[33807], Fresh[33806], Fresh[33805], Fresh[33804], Fresh[33803], Fresh[33802], Fresh[33801], Fresh[33800], Fresh[33799], Fresh[33798], Fresh[33797], Fresh[33796], Fresh[33795], Fresh[33794], Fresh[33793], Fresh[33792], Fresh[33791], Fresh[33790], Fresh[33789], Fresh[33788], Fresh[33787], Fresh[33786], Fresh[33785], Fresh[33784], Fresh[33783], Fresh[33782], Fresh[33781], Fresh[33780], Fresh[33779], Fresh[33778], Fresh[33777], Fresh[33776], Fresh[33775], Fresh[33774], Fresh[33773], Fresh[33772], Fresh[33771], Fresh[33770], Fresh[33769], Fresh[33768], Fresh[33767], Fresh[33766], Fresh[33765], Fresh[33764], Fresh[33763], Fresh[33762], Fresh[33761], Fresh[33760], Fresh[33759], Fresh[33758], Fresh[33757], Fresh[33756], Fresh[33755], Fresh[33754], Fresh[33753], Fresh[33752], Fresh[33751], Fresh[33750], Fresh[33749], Fresh[33748], Fresh[33747], Fresh[33746], Fresh[33745], Fresh[33744], Fresh[33743], Fresh[33742], Fresh[33741], Fresh[33740], Fresh[33739], Fresh[33738], Fresh[33737], Fresh[33736], Fresh[33735], Fresh[33734], Fresh[33733], Fresh[33732], Fresh[33731], Fresh[33730], Fresh[33729], Fresh[33728], Fresh[33727], Fresh[33726], Fresh[33725], Fresh[33724], Fresh[33723], Fresh[33722], Fresh[33721], Fresh[33720], Fresh[33719], Fresh[33718], Fresh[33717], Fresh[33716], Fresh[33715], Fresh[33714], Fresh[33713], Fresh[33712], Fresh[33711], Fresh[33710], Fresh[33709], Fresh[33708], Fresh[33707], Fresh[33706], Fresh[33705], Fresh[33704], Fresh[33703], Fresh[33702], Fresh[33701], Fresh[33700], Fresh[33699], Fresh[33698], Fresh[33697], Fresh[33696], Fresh[33695], Fresh[33694], Fresh[33693], Fresh[33692], Fresh[33691], Fresh[33690], Fresh[33689], Fresh[33688], Fresh[33687], Fresh[33686], Fresh[33685], Fresh[33684], Fresh[33683], Fresh[33682], Fresh[33681], Fresh[33680], Fresh[33679], Fresh[33678], Fresh[33677], Fresh[33676], Fresh[33675], Fresh[33674], Fresh[33673], Fresh[33672], Fresh[33671], Fresh[33670], Fresh[33669], Fresh[33668], Fresh[33667], Fresh[33666], Fresh[33665], Fresh[33664], Fresh[33663], Fresh[33662], Fresh[33661], Fresh[33660], Fresh[33659], Fresh[33658], Fresh[33657], Fresh[33656], Fresh[33655], Fresh[33654], Fresh[33653], Fresh[33652], Fresh[33651], Fresh[33650], Fresh[33649], Fresh[33648], Fresh[33647], Fresh[33646], Fresh[33645], Fresh[33644], Fresh[33643], Fresh[33642], Fresh[33641], Fresh[33640], Fresh[33639], Fresh[33638], Fresh[33637], Fresh[33636], Fresh[33635], Fresh[33634], Fresh[33633], Fresh[33632], Fresh[33631], Fresh[33630], Fresh[33629], Fresh[33628], Fresh[33627], Fresh[33626], Fresh[33625], Fresh[33624], Fresh[33623], Fresh[33622], Fresh[33621], Fresh[33620], Fresh[33619], Fresh[33618], Fresh[33617], Fresh[33616], Fresh[33615], Fresh[33614], Fresh[33613], Fresh[33612], Fresh[33611], Fresh[33610], Fresh[33609], Fresh[33608], Fresh[33607], Fresh[33606], Fresh[33605], Fresh[33604], Fresh[33603], Fresh[33602], Fresh[33601], Fresh[33600], Fresh[33599], Fresh[33598], Fresh[33597], Fresh[33596], Fresh[33595], Fresh[33594], Fresh[33593], Fresh[33592], Fresh[33591], Fresh[33590], Fresh[33589], Fresh[33588], Fresh[33587], Fresh[33586], Fresh[33585], Fresh[33584], Fresh[33583], Fresh[33582], Fresh[33581], Fresh[33580], Fresh[33579], Fresh[33578], Fresh[33577], Fresh[33576], Fresh[33575], Fresh[33574], Fresh[33573], Fresh[33572], Fresh[33571], Fresh[33570], Fresh[33569], Fresh[33568], Fresh[33567], Fresh[33566], Fresh[33565], Fresh[33564], Fresh[33563], Fresh[33562], Fresh[33561], Fresh[33560], Fresh[33559], Fresh[33558], Fresh[33557], Fresh[33556], Fresh[33555], Fresh[33554], Fresh[33553], Fresh[33552], Fresh[33551], Fresh[33550], Fresh[33549], Fresh[33548], Fresh[33547], Fresh[33546], Fresh[33545], Fresh[33544], Fresh[33543], Fresh[33542], Fresh[33541], Fresh[33540], Fresh[33539], Fresh[33538], Fresh[33537], Fresh[33536], Fresh[33535], Fresh[33534], Fresh[33533], Fresh[33532], Fresh[33531], Fresh[33530], Fresh[33529], Fresh[33528], Fresh[33527], Fresh[33526], Fresh[33525], Fresh[33524], Fresh[33523], Fresh[33522], Fresh[33521], Fresh[33520], Fresh[33519], Fresh[33518], Fresh[33517], Fresh[33516], Fresh[33515], Fresh[33514], Fresh[33513], Fresh[33512], Fresh[33511], Fresh[33510], Fresh[33509], Fresh[33508], Fresh[33507], Fresh[33506], Fresh[33505], Fresh[33504], Fresh[33503], Fresh[33502], Fresh[33501], Fresh[33500], Fresh[33499], Fresh[33498], Fresh[33497], Fresh[33496], Fresh[33495], Fresh[33494], Fresh[33493], Fresh[33492], Fresh[33491], Fresh[33490], Fresh[33489], Fresh[33488], Fresh[33487], Fresh[33486], Fresh[33485], Fresh[33484], Fresh[33483], Fresh[33482], Fresh[33481], Fresh[33480], Fresh[33479], Fresh[33478], Fresh[33477], Fresh[33476], Fresh[33475], Fresh[33474], Fresh[33473], Fresh[33472], Fresh[33471], Fresh[33470], Fresh[33469], Fresh[33468], Fresh[33467], Fresh[33466], Fresh[33465], Fresh[33464], Fresh[33463], Fresh[33462], Fresh[33461], Fresh[33460], Fresh[33459], Fresh[33458], Fresh[33457], Fresh[33456], Fresh[33455], Fresh[33454], Fresh[33453], Fresh[33452], Fresh[33451], Fresh[33450], Fresh[33449], Fresh[33448], Fresh[33447], Fresh[33446], Fresh[33445], Fresh[33444], Fresh[33443], Fresh[33442], Fresh[33441], Fresh[33440], Fresh[33439], Fresh[33438], Fresh[33437], Fresh[33436], Fresh[33435], Fresh[33434], Fresh[33433], Fresh[33432], Fresh[33431], Fresh[33430], Fresh[33429], Fresh[33428], Fresh[33427], Fresh[33426], Fresh[33425], Fresh[33424], Fresh[33423], Fresh[33422], Fresh[33421], Fresh[33420], Fresh[33419], Fresh[33418], Fresh[33417], Fresh[33416], Fresh[33415], Fresh[33414], Fresh[33413], Fresh[33412], Fresh[33411], Fresh[33410], Fresh[33409], Fresh[33408], Fresh[33407], Fresh[33406], Fresh[33405], Fresh[33404], Fresh[33403], Fresh[33402], Fresh[33401], Fresh[33400], Fresh[33399], Fresh[33398], Fresh[33397], Fresh[33396], Fresh[33395], Fresh[33394], Fresh[33393], Fresh[33392], Fresh[33391], Fresh[33390], Fresh[33389], Fresh[33388], Fresh[33387], Fresh[33386], Fresh[33385], Fresh[33384], Fresh[33383], Fresh[33382], Fresh[33381], Fresh[33380], Fresh[33379], Fresh[33378], Fresh[33377], Fresh[33376], Fresh[33375], Fresh[33374], Fresh[33373], Fresh[33372], Fresh[33371], Fresh[33370], Fresh[33369], Fresh[33368], Fresh[33367], Fresh[33366], Fresh[33365], Fresh[33364], Fresh[33363], Fresh[33362], Fresh[33361], Fresh[33360], Fresh[33359], Fresh[33358], Fresh[33357], Fresh[33356], Fresh[33355], Fresh[33354], Fresh[33353], Fresh[33352], Fresh[33351], Fresh[33350], Fresh[33349], Fresh[33348], Fresh[33347], Fresh[33346], Fresh[33345], Fresh[33344], Fresh[33343], Fresh[33342], Fresh[33341], Fresh[33340], Fresh[33339], Fresh[33338], Fresh[33337], Fresh[33336], Fresh[33335], Fresh[33334], Fresh[33333], Fresh[33332], Fresh[33331], Fresh[33330], Fresh[33329], Fresh[33328], Fresh[33327], Fresh[33326], Fresh[33325], Fresh[33324], Fresh[33323], Fresh[33322], Fresh[33321], Fresh[33320], Fresh[33319], Fresh[33318], Fresh[33317], Fresh[33316], Fresh[33315], Fresh[33314], Fresh[33313], Fresh[33312], Fresh[33311], Fresh[33310], Fresh[33309], Fresh[33308], Fresh[33307], Fresh[33306], Fresh[33305], Fresh[33304], Fresh[33303], Fresh[33302], Fresh[33301], Fresh[33300], Fresh[33299], Fresh[33298], Fresh[33297], Fresh[33296], Fresh[33295], Fresh[33294], Fresh[33293], Fresh[33292], Fresh[33291], Fresh[33290], Fresh[33289], Fresh[33288], Fresh[33287], Fresh[33286], Fresh[33285], Fresh[33284], Fresh[33283], Fresh[33282], Fresh[33281], Fresh[33280], Fresh[33279], Fresh[33278], Fresh[33277], Fresh[33276], Fresh[33275], Fresh[33274], Fresh[33273], Fresh[33272], Fresh[33271], Fresh[33270], Fresh[33269], Fresh[33268], Fresh[33267], Fresh[33266], Fresh[33265], Fresh[33264], Fresh[33263], Fresh[33262], Fresh[33261], Fresh[33260], Fresh[33259], Fresh[33258], Fresh[33257], Fresh[33256], Fresh[33255], Fresh[33254], Fresh[33253], Fresh[33252], Fresh[33251], Fresh[33250], Fresh[33249], Fresh[33248], Fresh[33247], Fresh[33246], Fresh[33245], Fresh[33244], Fresh[33243], Fresh[33242], Fresh[33241], Fresh[33240], Fresh[33239], Fresh[33238], Fresh[33237], Fresh[33236], Fresh[33235], Fresh[33234], Fresh[33233], Fresh[33232], Fresh[33231], Fresh[33230], Fresh[33229], Fresh[33228], Fresh[33227], Fresh[33226], Fresh[33225], Fresh[33224], Fresh[33223], Fresh[33222], Fresh[33221], Fresh[33220], Fresh[33219], Fresh[33218], Fresh[33217], Fresh[33216], Fresh[33215], Fresh[33214], Fresh[33213], Fresh[33212], Fresh[33211], Fresh[33210], Fresh[33209], Fresh[33208], Fresh[33207], Fresh[33206], Fresh[33205], Fresh[33204], Fresh[33203], Fresh[33202], Fresh[33201], Fresh[33200], Fresh[33199], Fresh[33198], Fresh[33197], Fresh[33196], Fresh[33195], Fresh[33194], Fresh[33193], Fresh[33192], Fresh[33191], Fresh[33190], Fresh[33189], Fresh[33188], Fresh[33187], Fresh[33186], Fresh[33185], Fresh[33184], Fresh[33183], Fresh[33182], Fresh[33181], Fresh[33180], Fresh[33179], Fresh[33178], Fresh[33177], Fresh[33176], Fresh[33175], Fresh[33174], Fresh[33173], Fresh[33172], Fresh[33171], Fresh[33170], Fresh[33169], Fresh[33168], Fresh[33167], Fresh[33166], Fresh[33165], Fresh[33164], Fresh[33163], Fresh[33162], Fresh[33161], Fresh[33160], Fresh[33159], Fresh[33158], Fresh[33157], Fresh[33156], Fresh[33155], Fresh[33154], Fresh[33153], Fresh[33152], Fresh[33151], Fresh[33150], Fresh[33149], Fresh[33148], Fresh[33147], Fresh[33146], Fresh[33145], Fresh[33144], Fresh[33143], Fresh[33142], Fresh[33141], Fresh[33140], Fresh[33139], Fresh[33138], Fresh[33137], Fresh[33136], Fresh[33135], Fresh[33134], Fresh[33133], Fresh[33132], Fresh[33131], Fresh[33130], Fresh[33129], Fresh[33128], Fresh[33127], Fresh[33126], Fresh[33125], Fresh[33124], Fresh[33123], Fresh[33122], Fresh[33121], Fresh[33120], Fresh[33119], Fresh[33118], Fresh[33117], Fresh[33116], Fresh[33115], Fresh[33114], Fresh[33113], Fresh[33112], Fresh[33111], Fresh[33110], Fresh[33109], Fresh[33108], Fresh[33107], Fresh[33106], Fresh[33105], Fresh[33104], Fresh[33103], Fresh[33102], Fresh[33101], Fresh[33100], Fresh[33099], Fresh[33098], Fresh[33097], Fresh[33096], Fresh[33095], Fresh[33094], Fresh[33093], Fresh[33092], Fresh[33091], Fresh[33090], Fresh[33089], Fresh[33088], Fresh[33087], Fresh[33086], Fresh[33085], Fresh[33084], Fresh[33083], Fresh[33082], Fresh[33081], Fresh[33080], Fresh[33079], Fresh[33078], Fresh[33077], Fresh[33076], Fresh[33075], Fresh[33074], Fresh[33073], Fresh[33072], Fresh[33071], Fresh[33070], Fresh[33069], Fresh[33068], Fresh[33067], Fresh[33066], Fresh[33065], Fresh[33064], Fresh[33063], Fresh[33062], Fresh[33061], Fresh[33060], Fresh[33059], Fresh[33058], Fresh[33057], Fresh[33056], Fresh[33055], Fresh[33054], Fresh[33053], Fresh[33052], Fresh[33051], Fresh[33050], Fresh[33049], Fresh[33048], Fresh[33047], Fresh[33046], Fresh[33045], Fresh[33044], Fresh[33043], Fresh[33042], Fresh[33041], Fresh[33040], Fresh[33039], Fresh[33038], Fresh[33037], Fresh[33036], Fresh[33035], Fresh[33034], Fresh[33033], Fresh[33032], Fresh[33031], Fresh[33030], Fresh[33029], Fresh[33028], Fresh[33027], Fresh[33026], Fresh[33025], Fresh[33024], Fresh[33023], Fresh[33022], Fresh[33021], Fresh[33020], Fresh[33019], Fresh[33018], Fresh[33017], Fresh[33016], Fresh[33015], Fresh[33014], Fresh[33013], Fresh[33012], Fresh[33011], Fresh[33010], Fresh[33009], Fresh[33008], Fresh[33007], Fresh[33006], Fresh[33005], Fresh[33004], Fresh[33003], Fresh[33002], Fresh[33001], Fresh[33000], Fresh[32999], Fresh[32998], Fresh[32997], Fresh[32996], Fresh[32995], Fresh[32994], Fresh[32993], Fresh[32992], Fresh[32991], Fresh[32990], Fresh[32989], Fresh[32988], Fresh[32987], Fresh[32986], Fresh[32985], Fresh[32984], Fresh[32983], Fresh[32982], Fresh[32981], Fresh[32980], Fresh[32979], Fresh[32978], Fresh[32977], Fresh[32976], Fresh[32975], Fresh[32974], Fresh[32973], Fresh[32972], Fresh[32971], Fresh[32970], Fresh[32969], Fresh[32968], Fresh[32967], Fresh[32966], Fresh[32965], Fresh[32964], Fresh[32963], Fresh[32962], Fresh[32961], Fresh[32960], Fresh[32959], Fresh[32958], Fresh[32957], Fresh[32956], Fresh[32955], Fresh[32954], Fresh[32953], Fresh[32952], Fresh[32951], Fresh[32950], Fresh[32949], Fresh[32948], Fresh[32947], Fresh[32946], Fresh[32945], Fresh[32944], Fresh[32943], Fresh[32942], Fresh[32941], Fresh[32940], Fresh[32939], Fresh[32938], Fresh[32937], Fresh[32936], Fresh[32935], Fresh[32934], Fresh[32933], Fresh[32932], Fresh[32931], Fresh[32930], Fresh[32929], Fresh[32928], Fresh[32927], Fresh[32926], Fresh[32925], Fresh[32924], Fresh[32923], Fresh[32922], Fresh[32921], Fresh[32920], Fresh[32919], Fresh[32918], Fresh[32917], Fresh[32916], Fresh[32915], Fresh[32914], Fresh[32913], Fresh[32912], Fresh[32911], Fresh[32910], Fresh[32909], Fresh[32908], Fresh[32907], Fresh[32906], Fresh[32905], Fresh[32904], Fresh[32903], Fresh[32902], Fresh[32901], Fresh[32900], Fresh[32899], Fresh[32898], Fresh[32897], Fresh[32896], Fresh[32895], Fresh[32894], Fresh[32893], Fresh[32892], Fresh[32891], Fresh[32890], Fresh[32889], Fresh[32888], Fresh[32887], Fresh[32886], Fresh[32885], Fresh[32884], Fresh[32883], Fresh[32882], Fresh[32881], Fresh[32880], Fresh[32879], Fresh[32878], Fresh[32877], Fresh[32876], Fresh[32875], Fresh[32874], Fresh[32873], Fresh[32872], Fresh[32871], Fresh[32870], Fresh[32869], Fresh[32868], Fresh[32867], Fresh[32866], Fresh[32865], Fresh[32864], Fresh[32863], Fresh[32862], Fresh[32861], Fresh[32860], Fresh[32859], Fresh[32858], Fresh[32857], Fresh[32856], Fresh[32855], Fresh[32854], Fresh[32853], Fresh[32852], Fresh[32851], Fresh[32850], Fresh[32849], Fresh[32848], Fresh[32847], Fresh[32846], Fresh[32845], Fresh[32844], Fresh[32843], Fresh[32842], Fresh[32841], Fresh[32840], Fresh[32839], Fresh[32838], Fresh[32837], Fresh[32836], Fresh[32835], Fresh[32834], Fresh[32833], Fresh[32832], Fresh[32831], Fresh[32830], Fresh[32829], Fresh[32828], Fresh[32827], Fresh[32826], Fresh[32825], Fresh[32824], Fresh[32823], Fresh[32822], Fresh[32821], Fresh[32820], Fresh[32819], Fresh[32818], Fresh[32817], Fresh[32816], Fresh[32815], Fresh[32814], Fresh[32813], Fresh[32812], Fresh[32811], Fresh[32810], Fresh[32809], Fresh[32808], Fresh[32807], Fresh[32806], Fresh[32805], Fresh[32804], Fresh[32803], Fresh[32802], Fresh[32801], Fresh[32800], Fresh[32799], Fresh[32798], Fresh[32797], Fresh[32796], Fresh[32795], Fresh[32794], Fresh[32793], Fresh[32792], Fresh[32791], Fresh[32790], Fresh[32789], Fresh[32788], Fresh[32787], Fresh[32786], Fresh[32785], Fresh[32784], Fresh[32783], Fresh[32782], Fresh[32781], Fresh[32780], Fresh[32779], Fresh[32778], Fresh[32777], Fresh[32776], Fresh[32775], Fresh[32774], Fresh[32773], Fresh[32772], Fresh[32771], Fresh[32770], Fresh[32769], Fresh[32768], Fresh[32767], Fresh[32766], Fresh[32765], Fresh[32764], Fresh[32763], Fresh[32762], Fresh[32761], Fresh[32760], Fresh[32759], Fresh[32758], Fresh[32757], Fresh[32756], Fresh[32755], Fresh[32754], Fresh[32753], Fresh[32752], Fresh[32751], Fresh[32750], Fresh[32749], Fresh[32748], Fresh[32747], Fresh[32746], Fresh[32745], Fresh[32744], Fresh[32743], Fresh[32742], Fresh[32741], Fresh[32740], Fresh[32739], Fresh[32738], Fresh[32737], Fresh[32736], Fresh[32735], Fresh[32734], Fresh[32733], Fresh[32732], Fresh[32731], Fresh[32730], Fresh[32729], Fresh[32728], Fresh[32727], Fresh[32726], Fresh[32725], Fresh[32724], Fresh[32723], Fresh[32722], Fresh[32721], Fresh[32720], Fresh[32719], Fresh[32718], Fresh[32717], Fresh[32716], Fresh[32715], Fresh[32714], Fresh[32713], Fresh[32712], Fresh[32711], Fresh[32710], Fresh[32709], Fresh[32708], Fresh[32707], Fresh[32706], Fresh[32705], Fresh[32704], Fresh[32703], Fresh[32702], Fresh[32701], Fresh[32700], Fresh[32699], Fresh[32698], Fresh[32697], Fresh[32696], Fresh[32695], Fresh[32694], Fresh[32693], Fresh[32692], Fresh[32691], Fresh[32690], Fresh[32689], Fresh[32688], Fresh[32687], Fresh[32686], Fresh[32685], Fresh[32684], Fresh[32683], Fresh[32682], Fresh[32681], Fresh[32680], Fresh[32679], Fresh[32678], Fresh[32677], Fresh[32676], Fresh[32675], Fresh[32674], Fresh[32673], Fresh[32672], Fresh[32671], Fresh[32670], Fresh[32669], Fresh[32668], Fresh[32667], Fresh[32666], Fresh[32665], Fresh[32664], Fresh[32663], Fresh[32662], Fresh[32661], Fresh[32660], Fresh[32659], Fresh[32658], Fresh[32657], Fresh[32656], Fresh[32655], Fresh[32654], Fresh[32653], Fresh[32652], Fresh[32651], Fresh[32650], Fresh[32649], Fresh[32648], Fresh[32647], Fresh[32646], Fresh[32645], Fresh[32644], Fresh[32643], Fresh[32642], Fresh[32641], Fresh[32640], Fresh[32639], Fresh[32638], Fresh[32637], Fresh[32636], Fresh[32635], Fresh[32634], Fresh[32633], Fresh[32632], Fresh[32631], Fresh[32630], Fresh[32629], Fresh[32628], Fresh[32627], Fresh[32626], Fresh[32625], Fresh[32624], Fresh[32623], Fresh[32622], Fresh[32621], Fresh[32620], Fresh[32619], Fresh[32618], Fresh[32617], Fresh[32616], Fresh[32615], Fresh[32614], Fresh[32613], Fresh[32612], Fresh[32611], Fresh[32610], Fresh[32609], Fresh[32608], Fresh[32607], Fresh[32606], Fresh[32605], Fresh[32604], Fresh[32603], Fresh[32602], Fresh[32601], Fresh[32600], Fresh[32599], Fresh[32598], Fresh[32597], Fresh[32596], Fresh[32595], Fresh[32594], Fresh[32593], Fresh[32592], Fresh[32591], Fresh[32590], Fresh[32589], Fresh[32588], Fresh[32587], Fresh[32586], Fresh[32585], Fresh[32584], Fresh[32583], Fresh[32582], Fresh[32581], Fresh[32580], Fresh[32579], Fresh[32578], Fresh[32577], Fresh[32576], Fresh[32575], Fresh[32574], Fresh[32573], Fresh[32572], Fresh[32571], Fresh[32570], Fresh[32569], Fresh[32568], Fresh[32567], Fresh[32566], Fresh[32565], Fresh[32564], Fresh[32563], Fresh[32562], Fresh[32561], Fresh[32560], Fresh[32559], Fresh[32558], Fresh[32557], Fresh[32556], Fresh[32555], Fresh[32554], Fresh[32553], Fresh[32552], Fresh[32551], Fresh[32550], Fresh[32549], Fresh[32548], Fresh[32547], Fresh[32546], Fresh[32545], Fresh[32544], Fresh[32543], Fresh[32542], Fresh[32541], Fresh[32540], Fresh[32539], Fresh[32538], Fresh[32537], Fresh[32536], Fresh[32535], Fresh[32534], Fresh[32533], Fresh[32532], Fresh[32531], Fresh[32530], Fresh[32529], Fresh[32528], Fresh[32527], Fresh[32526], Fresh[32525], Fresh[32524], Fresh[32523], Fresh[32522], Fresh[32521], Fresh[32520], Fresh[32519], Fresh[32518], Fresh[32517], Fresh[32516], Fresh[32515], Fresh[32514], Fresh[32513], Fresh[32512], Fresh[32511], Fresh[32510], Fresh[32509], Fresh[32508], Fresh[32507], Fresh[32506], Fresh[32505], Fresh[32504], Fresh[32503], Fresh[32502], Fresh[32501], Fresh[32500], Fresh[32499], Fresh[32498], Fresh[32497], Fresh[32496], Fresh[32495], Fresh[32494], Fresh[32493], Fresh[32492], Fresh[32491], Fresh[32490], Fresh[32489], Fresh[32488], Fresh[32487], Fresh[32486], Fresh[32485], Fresh[32484], Fresh[32483], Fresh[32482], Fresh[32481], Fresh[32480], Fresh[32479], Fresh[32478], Fresh[32477], Fresh[32476], Fresh[32475], Fresh[32474], Fresh[32473], Fresh[32472], Fresh[32471], Fresh[32470], Fresh[32469], Fresh[32468], Fresh[32467], Fresh[32466], Fresh[32465], Fresh[32464], Fresh[32463], Fresh[32462], Fresh[32461], Fresh[32460], Fresh[32459], Fresh[32458], Fresh[32457], Fresh[32456], Fresh[32455], Fresh[32454], Fresh[32453], Fresh[32452], Fresh[32451], Fresh[32450], Fresh[32449], Fresh[32448], Fresh[32447], Fresh[32446], Fresh[32445], Fresh[32444], Fresh[32443], Fresh[32442], Fresh[32441], Fresh[32440], Fresh[32439], Fresh[32438], Fresh[32437], Fresh[32436], Fresh[32435], Fresh[32434], Fresh[32433], Fresh[32432], Fresh[32431], Fresh[32430], Fresh[32429], Fresh[32428], Fresh[32427], Fresh[32426], Fresh[32425], Fresh[32424], Fresh[32423], Fresh[32422], Fresh[32421], Fresh[32420], Fresh[32419], Fresh[32418], Fresh[32417], Fresh[32416], Fresh[32415], Fresh[32414], Fresh[32413], Fresh[32412], Fresh[32411], Fresh[32410], Fresh[32409], Fresh[32408], Fresh[32407], Fresh[32406], Fresh[32405], Fresh[32404], Fresh[32403], Fresh[32402], Fresh[32401], Fresh[32400], Fresh[32399], Fresh[32398], Fresh[32397], Fresh[32396], Fresh[32395], Fresh[32394], Fresh[32393], Fresh[32392], Fresh[32391], Fresh[32390], Fresh[32389], Fresh[32388], Fresh[32387], Fresh[32386], Fresh[32385], Fresh[32384], Fresh[32383], Fresh[32382], Fresh[32381], Fresh[32380], Fresh[32379], Fresh[32378], Fresh[32377], Fresh[32376], Fresh[32375], Fresh[32374], Fresh[32373], Fresh[32372], Fresh[32371], Fresh[32370], Fresh[32369], Fresh[32368], Fresh[32367], Fresh[32366], Fresh[32365], Fresh[32364], Fresh[32363], Fresh[32362], Fresh[32361], Fresh[32360], Fresh[32359], Fresh[32358], Fresh[32357], Fresh[32356], Fresh[32355], Fresh[32354], Fresh[32353], Fresh[32352], Fresh[32351], Fresh[32350], Fresh[32349], Fresh[32348], Fresh[32347], Fresh[32346], Fresh[32345], Fresh[32344], Fresh[32343], Fresh[32342], Fresh[32341], Fresh[32340], Fresh[32339], Fresh[32338], Fresh[32337], Fresh[32336], Fresh[32335], Fresh[32334], Fresh[32333], Fresh[32332], Fresh[32331], Fresh[32330], Fresh[32329], Fresh[32328], Fresh[32327], Fresh[32326], Fresh[32325], Fresh[32324], Fresh[32323], Fresh[32322], Fresh[32321], Fresh[32320], Fresh[32319], Fresh[32318], Fresh[32317], Fresh[32316], Fresh[32315], Fresh[32314], Fresh[32313], Fresh[32312], Fresh[32311], Fresh[32310], Fresh[32309], Fresh[32308], Fresh[32307], Fresh[32306], Fresh[32305], Fresh[32304], Fresh[32303], Fresh[32302], Fresh[32301], Fresh[32300], Fresh[32299], Fresh[32298], Fresh[32297], Fresh[32296], Fresh[32295], Fresh[32294], Fresh[32293], Fresh[32292], Fresh[32291], Fresh[32290], Fresh[32289], Fresh[32288], Fresh[32287], Fresh[32286], Fresh[32285], Fresh[32284], Fresh[32283], Fresh[32282], Fresh[32281], Fresh[32280], Fresh[32279], Fresh[32278], Fresh[32277], Fresh[32276], Fresh[32275], Fresh[32274], Fresh[32273], Fresh[32272], Fresh[32271], Fresh[32270], Fresh[32269], Fresh[32268], Fresh[32267], Fresh[32266], Fresh[32265], Fresh[32264], Fresh[32263], Fresh[32262], Fresh[32261], Fresh[32260], Fresh[32259], Fresh[32258], Fresh[32257], Fresh[32256], Fresh[32255], Fresh[32254], Fresh[32253], Fresh[32252], Fresh[32251], Fresh[32250], Fresh[32249], Fresh[32248], Fresh[32247], Fresh[32246], Fresh[32245], Fresh[32244], Fresh[32243], Fresh[32242], Fresh[32241], Fresh[32240], Fresh[32239], Fresh[32238], Fresh[32237], Fresh[32236], Fresh[32235], Fresh[32234], Fresh[32233], Fresh[32232], Fresh[32231], Fresh[32230], Fresh[32229], Fresh[32228], Fresh[32227], Fresh[32226], Fresh[32225], Fresh[32224], Fresh[32223], Fresh[32222], Fresh[32221], Fresh[32220], Fresh[32219], Fresh[32218], Fresh[32217], Fresh[32216], Fresh[32215], Fresh[32214], Fresh[32213], Fresh[32212], Fresh[32211], Fresh[32210], Fresh[32209], Fresh[32208], Fresh[32207], Fresh[32206], Fresh[32205], Fresh[32204], Fresh[32203], Fresh[32202], Fresh[32201], Fresh[32200], Fresh[32199], Fresh[32198], Fresh[32197], Fresh[32196], Fresh[32195], Fresh[32194], Fresh[32193], Fresh[32192], Fresh[32191], Fresh[32190], Fresh[32189], Fresh[32188], Fresh[32187], Fresh[32186], Fresh[32185], Fresh[32184], Fresh[32183], Fresh[32182], Fresh[32181], Fresh[32180], Fresh[32179], Fresh[32178], Fresh[32177], Fresh[32176], Fresh[32175], Fresh[32174], Fresh[32173], Fresh[32172], Fresh[32171], Fresh[32170], Fresh[32169], Fresh[32168], Fresh[32167], Fresh[32166], Fresh[32165], Fresh[32164], Fresh[32163], Fresh[32162], Fresh[32161], Fresh[32160], Fresh[32159], Fresh[32158], Fresh[32157], Fresh[32156], Fresh[32155], Fresh[32154], Fresh[32153], Fresh[32152], Fresh[32151], Fresh[32150], Fresh[32149], Fresh[32148], Fresh[32147], Fresh[32146], Fresh[32145], Fresh[32144], Fresh[32143], Fresh[32142], Fresh[32141], Fresh[32140], Fresh[32139], Fresh[32138], Fresh[32137], Fresh[32136], Fresh[32135], Fresh[32134], Fresh[32133], Fresh[32132], Fresh[32131], Fresh[32130], Fresh[32129], Fresh[32128], Fresh[32127], Fresh[32126], Fresh[32125], Fresh[32124], Fresh[32123], Fresh[32122], Fresh[32121], Fresh[32120], Fresh[32119], Fresh[32118], Fresh[32117], Fresh[32116], Fresh[32115], Fresh[32114], Fresh[32113], Fresh[32112], Fresh[32111], Fresh[32110], Fresh[32109], Fresh[32108], Fresh[32107], Fresh[32106], Fresh[32105], Fresh[32104], Fresh[32103], Fresh[32102], Fresh[32101], Fresh[32100], Fresh[32099], Fresh[32098], Fresh[32097], Fresh[32096], Fresh[32095], Fresh[32094], Fresh[32093], Fresh[32092], Fresh[32091], Fresh[32090], Fresh[32089], Fresh[32088], Fresh[32087], Fresh[32086], Fresh[32085], Fresh[32084], Fresh[32083], Fresh[32082], Fresh[32081], Fresh[32080], Fresh[32079], Fresh[32078], Fresh[32077], Fresh[32076], Fresh[32075], Fresh[32074], Fresh[32073], Fresh[32072], Fresh[32071], Fresh[32070], Fresh[32069], Fresh[32068], Fresh[32067], Fresh[32066], Fresh[32065], Fresh[32064], Fresh[32063], Fresh[32062], Fresh[32061], Fresh[32060], Fresh[32059], Fresh[32058], Fresh[32057], Fresh[32056], Fresh[32055], Fresh[32054], Fresh[32053], Fresh[32052], Fresh[32051], Fresh[32050], Fresh[32049], Fresh[32048], Fresh[32047], Fresh[32046], Fresh[32045], Fresh[32044], Fresh[32043], Fresh[32042], Fresh[32041], Fresh[32040], Fresh[32039], Fresh[32038], Fresh[32037], Fresh[32036], Fresh[32035], Fresh[32034], Fresh[32033], Fresh[32032], Fresh[32031], Fresh[32030], Fresh[32029], Fresh[32028], Fresh[32027], Fresh[32026], Fresh[32025], Fresh[32024], Fresh[32023], Fresh[32022], Fresh[32021], Fresh[32020], Fresh[32019], Fresh[32018], Fresh[32017], Fresh[32016], Fresh[32015], Fresh[32014], Fresh[32013], Fresh[32012], Fresh[32011], Fresh[32010], Fresh[32009], Fresh[32008], Fresh[32007], Fresh[32006], Fresh[32005], Fresh[32004], Fresh[32003], Fresh[32002], Fresh[32001], Fresh[32000], Fresh[31999], Fresh[31998], Fresh[31997], Fresh[31996], Fresh[31995], Fresh[31994], Fresh[31993], Fresh[31992], Fresh[31991], Fresh[31990], Fresh[31989], Fresh[31988], Fresh[31987], Fresh[31986], Fresh[31985], Fresh[31984], Fresh[31983], Fresh[31982], Fresh[31981], Fresh[31980], Fresh[31979], Fresh[31978], Fresh[31977], Fresh[31976], Fresh[31975], Fresh[31974], Fresh[31973], Fresh[31972], Fresh[31971], Fresh[31970], Fresh[31969], Fresh[31968], Fresh[31967], Fresh[31966], Fresh[31965], Fresh[31964], Fresh[31963], Fresh[31962], Fresh[31961], Fresh[31960], Fresh[31959], Fresh[31958], Fresh[31957], Fresh[31956], Fresh[31955], Fresh[31954], Fresh[31953], Fresh[31952], Fresh[31951], Fresh[31950], Fresh[31949], Fresh[31948], Fresh[31947], Fresh[31946], Fresh[31945], Fresh[31944], Fresh[31943], Fresh[31942], Fresh[31941], Fresh[31940], Fresh[31939], Fresh[31938], Fresh[31937], Fresh[31936], Fresh[31935], Fresh[31934], Fresh[31933], Fresh[31932], Fresh[31931], Fresh[31930], Fresh[31929], Fresh[31928], Fresh[31927], Fresh[31926], Fresh[31925], Fresh[31924], Fresh[31923], Fresh[31922], Fresh[31921], Fresh[31920], Fresh[31919], Fresh[31918], Fresh[31917], Fresh[31916], Fresh[31915], Fresh[31914], Fresh[31913], Fresh[31912], Fresh[31911], Fresh[31910], Fresh[31909], Fresh[31908], Fresh[31907], Fresh[31906], Fresh[31905], Fresh[31904], Fresh[31903], Fresh[31902], Fresh[31901], Fresh[31900], Fresh[31899], Fresh[31898], Fresh[31897], Fresh[31896], Fresh[31895], Fresh[31894], Fresh[31893], Fresh[31892], Fresh[31891], Fresh[31890], Fresh[31889], Fresh[31888], Fresh[31887], Fresh[31886], Fresh[31885], Fresh[31884], Fresh[31883], Fresh[31882], Fresh[31881], Fresh[31880], Fresh[31879], Fresh[31878], Fresh[31877], Fresh[31876], Fresh[31875], Fresh[31874], Fresh[31873], Fresh[31872], Fresh[31871], Fresh[31870], Fresh[31869], Fresh[31868], Fresh[31867], Fresh[31866], Fresh[31865], Fresh[31864], Fresh[31863], Fresh[31862], Fresh[31861], Fresh[31860], Fresh[31859], Fresh[31858], Fresh[31857], Fresh[31856], Fresh[31855], Fresh[31854], Fresh[31853], Fresh[31852], Fresh[31851], Fresh[31850], Fresh[31849], Fresh[31848], Fresh[31847], Fresh[31846], Fresh[31845], Fresh[31844], Fresh[31843], Fresh[31842], Fresh[31841], Fresh[31840], Fresh[31839], Fresh[31838], Fresh[31837], Fresh[31836], Fresh[31835], Fresh[31834], Fresh[31833], Fresh[31832], Fresh[31831], Fresh[31830], Fresh[31829], Fresh[31828], Fresh[31827], Fresh[31826], Fresh[31825], Fresh[31824], Fresh[31823], Fresh[31822], Fresh[31821], Fresh[31820], Fresh[31819], Fresh[31818], Fresh[31817], Fresh[31816], Fresh[31815], Fresh[31814], Fresh[31813], Fresh[31812], Fresh[31811], Fresh[31810], Fresh[31809], Fresh[31808], Fresh[31807], Fresh[31806], Fresh[31805], Fresh[31804], Fresh[31803], Fresh[31802], Fresh[31801], Fresh[31800], Fresh[31799], Fresh[31798], Fresh[31797], Fresh[31796], Fresh[31795], Fresh[31794], Fresh[31793], Fresh[31792], Fresh[31791], Fresh[31790], Fresh[31789], Fresh[31788], Fresh[31787], Fresh[31786], Fresh[31785], Fresh[31784], Fresh[31783], Fresh[31782], Fresh[31781], Fresh[31780], Fresh[31779], Fresh[31778], Fresh[31777], Fresh[31776], Fresh[31775], Fresh[31774], Fresh[31773], Fresh[31772], Fresh[31771], Fresh[31770], Fresh[31769], Fresh[31768], Fresh[31767], Fresh[31766], Fresh[31765], Fresh[31764], Fresh[31763], Fresh[31762], Fresh[31761], Fresh[31760], Fresh[31759], Fresh[31758], Fresh[31757], Fresh[31756], Fresh[31755], Fresh[31754], Fresh[31753], Fresh[31752], Fresh[31751], Fresh[31750], Fresh[31749], Fresh[31748], Fresh[31747], Fresh[31746], Fresh[31745], Fresh[31744], Fresh[31743], Fresh[31742], Fresh[31741], Fresh[31740], Fresh[31739], Fresh[31738], Fresh[31737], Fresh[31736], Fresh[31735], Fresh[31734], Fresh[31733], Fresh[31732], Fresh[31731], Fresh[31730], Fresh[31729], Fresh[31728], Fresh[31727], Fresh[31726], Fresh[31725], Fresh[31724], Fresh[31723], Fresh[31722], Fresh[31721], Fresh[31720], Fresh[31719], Fresh[31718], Fresh[31717], Fresh[31716], Fresh[31715], Fresh[31714], Fresh[31713], Fresh[31712], Fresh[31711], Fresh[31710], Fresh[31709], Fresh[31708], Fresh[31707], Fresh[31706], Fresh[31705], Fresh[31704], Fresh[31703], Fresh[31702], Fresh[31701], Fresh[31700], Fresh[31699], Fresh[31698], Fresh[31697], Fresh[31696], Fresh[31695], Fresh[31694], Fresh[31693], Fresh[31692], Fresh[31691], Fresh[31690], Fresh[31689], Fresh[31688], Fresh[31687], Fresh[31686], Fresh[31685], Fresh[31684], Fresh[31683], Fresh[31682], Fresh[31681], Fresh[31680], Fresh[31679], Fresh[31678], Fresh[31677], Fresh[31676], Fresh[31675], Fresh[31674], Fresh[31673], Fresh[31672], Fresh[31671], Fresh[31670], Fresh[31669], Fresh[31668], Fresh[31667], Fresh[31666], Fresh[31665], Fresh[31664], Fresh[31663], Fresh[31662], Fresh[31661], Fresh[31660], Fresh[31659], Fresh[31658], Fresh[31657], Fresh[31656], Fresh[31655], Fresh[31654], Fresh[31653], Fresh[31652], Fresh[31651], Fresh[31650], Fresh[31649], Fresh[31648], Fresh[31647], Fresh[31646], Fresh[31645], Fresh[31644], Fresh[31643], Fresh[31642], Fresh[31641], Fresh[31640], Fresh[31639], Fresh[31638], Fresh[31637], Fresh[31636], Fresh[31635], Fresh[31634], Fresh[31633], Fresh[31632], Fresh[31631], Fresh[31630], Fresh[31629], Fresh[31628], Fresh[31627], Fresh[31626], Fresh[31625], Fresh[31624], Fresh[31623], Fresh[31622], Fresh[31621], Fresh[31620], Fresh[31619], Fresh[31618], Fresh[31617], Fresh[31616], Fresh[31615], Fresh[31614], Fresh[31613], Fresh[31612], Fresh[31611], Fresh[31610], Fresh[31609], Fresh[31608], Fresh[31607], Fresh[31606], Fresh[31605], Fresh[31604], Fresh[31603], Fresh[31602], Fresh[31601], Fresh[31600], Fresh[31599], Fresh[31598], Fresh[31597], Fresh[31596], Fresh[31595], Fresh[31594], Fresh[31593], Fresh[31592], Fresh[31591], Fresh[31590], Fresh[31589], Fresh[31588], Fresh[31587], Fresh[31586], Fresh[31585], Fresh[31584], Fresh[31583], Fresh[31582], Fresh[31581], Fresh[31580], Fresh[31579], Fresh[31578], Fresh[31577], Fresh[31576], Fresh[31575], Fresh[31574], Fresh[31573], Fresh[31572], Fresh[31571], Fresh[31570], Fresh[31569], Fresh[31568], Fresh[31567], Fresh[31566], Fresh[31565], Fresh[31564], Fresh[31563], Fresh[31562], Fresh[31561], Fresh[31560], Fresh[31559], Fresh[31558], Fresh[31557], Fresh[31556], Fresh[31555], Fresh[31554], Fresh[31553], Fresh[31552], Fresh[31551], Fresh[31550], Fresh[31549], Fresh[31548], Fresh[31547], Fresh[31546], Fresh[31545], Fresh[31544], Fresh[31543], Fresh[31542], Fresh[31541], Fresh[31540], Fresh[31539], Fresh[31538], Fresh[31537], Fresh[31536], Fresh[31535], Fresh[31534], Fresh[31533], Fresh[31532], Fresh[31531], Fresh[31530], Fresh[31529], Fresh[31528], Fresh[31527], Fresh[31526], Fresh[31525], Fresh[31524], Fresh[31523], Fresh[31522], Fresh[31521], Fresh[31520], Fresh[31519], Fresh[31518], Fresh[31517], Fresh[31516], Fresh[31515], Fresh[31514], Fresh[31513], Fresh[31512], Fresh[31511], Fresh[31510], Fresh[31509], Fresh[31508], Fresh[31507], Fresh[31506], Fresh[31505], Fresh[31504], Fresh[31503], Fresh[31502], Fresh[31501], Fresh[31500], Fresh[31499], Fresh[31498], Fresh[31497], Fresh[31496], Fresh[31495], Fresh[31494], Fresh[31493], Fresh[31492], Fresh[31491], Fresh[31490], Fresh[31489], Fresh[31488], Fresh[31487], Fresh[31486], Fresh[31485], Fresh[31484], Fresh[31483], Fresh[31482], Fresh[31481], Fresh[31480], Fresh[31479], Fresh[31478], Fresh[31477], Fresh[31476], Fresh[31475], Fresh[31474], Fresh[31473], Fresh[31472], Fresh[31471], Fresh[31470], Fresh[31469], Fresh[31468], Fresh[31467], Fresh[31466], Fresh[31465], Fresh[31464], Fresh[31463], Fresh[31462], Fresh[31461], Fresh[31460], Fresh[31459], Fresh[31458], Fresh[31457], Fresh[31456], Fresh[31455], Fresh[31454], Fresh[31453], Fresh[31452], Fresh[31451], Fresh[31450], Fresh[31449], Fresh[31448], Fresh[31447], Fresh[31446], Fresh[31445], Fresh[31444], Fresh[31443], Fresh[31442], Fresh[31441], Fresh[31440], Fresh[31439], Fresh[31438], Fresh[31437], Fresh[31436], Fresh[31435], Fresh[31434], Fresh[31433], Fresh[31432], Fresh[31431], Fresh[31430], Fresh[31429], Fresh[31428], Fresh[31427], Fresh[31426], Fresh[31425], Fresh[31424], Fresh[31423], Fresh[31422], Fresh[31421], Fresh[31420], Fresh[31419], Fresh[31418], Fresh[31417], Fresh[31416], Fresh[31415], Fresh[31414], Fresh[31413], Fresh[31412], Fresh[31411], Fresh[31410], Fresh[31409], Fresh[31408], Fresh[31407], Fresh[31406], Fresh[31405], Fresh[31404], Fresh[31403], Fresh[31402], Fresh[31401], Fresh[31400], Fresh[31399], Fresh[31398], Fresh[31397], Fresh[31396], Fresh[31395], Fresh[31394], Fresh[31393], Fresh[31392], Fresh[31391], Fresh[31390], Fresh[31389], Fresh[31388], Fresh[31387], Fresh[31386], Fresh[31385], Fresh[31384], Fresh[31383], Fresh[31382], Fresh[31381], Fresh[31380], Fresh[31379], Fresh[31378], Fresh[31377], Fresh[31376], Fresh[31375], Fresh[31374], Fresh[31373], Fresh[31372], Fresh[31371], Fresh[31370], Fresh[31369], Fresh[31368], Fresh[31367], Fresh[31366], Fresh[31365], Fresh[31364], Fresh[31363], Fresh[31362], Fresh[31361], Fresh[31360], Fresh[31359], Fresh[31358], Fresh[31357], Fresh[31356], Fresh[31355], Fresh[31354], Fresh[31353], Fresh[31352], Fresh[31351], Fresh[31350], Fresh[31349], Fresh[31348], Fresh[31347], Fresh[31346], Fresh[31345], Fresh[31344], Fresh[31343], Fresh[31342], Fresh[31341], Fresh[31340], Fresh[31339], Fresh[31338], Fresh[31337], Fresh[31336], Fresh[31335], Fresh[31334], Fresh[31333], Fresh[31332], Fresh[31331], Fresh[31330], Fresh[31329], Fresh[31328], Fresh[31327], Fresh[31326], Fresh[31325], Fresh[31324], Fresh[31323], Fresh[31322], Fresh[31321], Fresh[31320], Fresh[31319], Fresh[31318], Fresh[31317], Fresh[31316], Fresh[31315], Fresh[31314], Fresh[31313], Fresh[31312], Fresh[31311], Fresh[31310], Fresh[31309], Fresh[31308], Fresh[31307], Fresh[31306], Fresh[31305], Fresh[31304], Fresh[31303], Fresh[31302], Fresh[31301], Fresh[31300], Fresh[31299], Fresh[31298], Fresh[31297], Fresh[31296], Fresh[31295], Fresh[31294], Fresh[31293], Fresh[31292], Fresh[31291], Fresh[31290], Fresh[31289], Fresh[31288], Fresh[31287], Fresh[31286], Fresh[31285], Fresh[31284], Fresh[31283], Fresh[31282], Fresh[31281], Fresh[31280], Fresh[31279], Fresh[31278], Fresh[31277], Fresh[31276], Fresh[31275], Fresh[31274], Fresh[31273], Fresh[31272], Fresh[31271], Fresh[31270], Fresh[31269], Fresh[31268], Fresh[31267], Fresh[31266], Fresh[31265], Fresh[31264], Fresh[31263], Fresh[31262], Fresh[31261], Fresh[31260], Fresh[31259], Fresh[31258], Fresh[31257], Fresh[31256], Fresh[31255], Fresh[31254], Fresh[31253], Fresh[31252], Fresh[31251], Fresh[31250], Fresh[31249], Fresh[31248], Fresh[31247], Fresh[31246], Fresh[31245], Fresh[31244], Fresh[31243], Fresh[31242], Fresh[31241], Fresh[31240], Fresh[31239], Fresh[31238], Fresh[31237], Fresh[31236], Fresh[31235], Fresh[31234], Fresh[31233], Fresh[31232], Fresh[31231], Fresh[31230], Fresh[31229], Fresh[31228], Fresh[31227], Fresh[31226], Fresh[31225], Fresh[31224], Fresh[31223], Fresh[31222], Fresh[31221], Fresh[31220], Fresh[31219], Fresh[31218], Fresh[31217], Fresh[31216], Fresh[31215], Fresh[31214], Fresh[31213], Fresh[31212], Fresh[31211], Fresh[31210], Fresh[31209], Fresh[31208], Fresh[31207], Fresh[31206], Fresh[31205], Fresh[31204], Fresh[31203], Fresh[31202], Fresh[31201], Fresh[31200], Fresh[31199], Fresh[31198], Fresh[31197], Fresh[31196], Fresh[31195], Fresh[31194], Fresh[31193], Fresh[31192], Fresh[31191], Fresh[31190], Fresh[31189], Fresh[31188], Fresh[31187], Fresh[31186], Fresh[31185], Fresh[31184], Fresh[31183], Fresh[31182], Fresh[31181], Fresh[31180], Fresh[31179], Fresh[31178], Fresh[31177], Fresh[31176], Fresh[31175], Fresh[31174], Fresh[31173], Fresh[31172], Fresh[31171], Fresh[31170], Fresh[31169], Fresh[31168], Fresh[31167], Fresh[31166], Fresh[31165], Fresh[31164], Fresh[31163], Fresh[31162], Fresh[31161], Fresh[31160], Fresh[31159], Fresh[31158], Fresh[31157], Fresh[31156], Fresh[31155], Fresh[31154], Fresh[31153], Fresh[31152], Fresh[31151], Fresh[31150], Fresh[31149], Fresh[31148], Fresh[31147], Fresh[31146], Fresh[31145], Fresh[31144], Fresh[31143], Fresh[31142], Fresh[31141], Fresh[31140], Fresh[31139], Fresh[31138], Fresh[31137], Fresh[31136], Fresh[31135], Fresh[31134], Fresh[31133], Fresh[31132], Fresh[31131], Fresh[31130], Fresh[31129], Fresh[31128], Fresh[31127], Fresh[31126], Fresh[31125], Fresh[31124], Fresh[31123], Fresh[31122], Fresh[31121], Fresh[31120], Fresh[31119], Fresh[31118], Fresh[31117], Fresh[31116], Fresh[31115], Fresh[31114], Fresh[31113], Fresh[31112], Fresh[31111], Fresh[31110], Fresh[31109], Fresh[31108], Fresh[31107], Fresh[31106], Fresh[31105], Fresh[31104], Fresh[31103], Fresh[31102], Fresh[31101], Fresh[31100], Fresh[31099], Fresh[31098], Fresh[31097], Fresh[31096], Fresh[31095], Fresh[31094], Fresh[31093], Fresh[31092], Fresh[31091], Fresh[31090], Fresh[31089], Fresh[31088], Fresh[31087], Fresh[31086], Fresh[31085], Fresh[31084], Fresh[31083], Fresh[31082], Fresh[31081], Fresh[31080], Fresh[31079], Fresh[31078], Fresh[31077], Fresh[31076], Fresh[31075], Fresh[31074], Fresh[31073], Fresh[31072], Fresh[31071], Fresh[31070], Fresh[31069], Fresh[31068], Fresh[31067], Fresh[31066], Fresh[31065], Fresh[31064], Fresh[31063], Fresh[31062], Fresh[31061], Fresh[31060], Fresh[31059], Fresh[31058], Fresh[31057], Fresh[31056], Fresh[31055], Fresh[31054], Fresh[31053], Fresh[31052], Fresh[31051], Fresh[31050], Fresh[31049], Fresh[31048], Fresh[31047], Fresh[31046], Fresh[31045], Fresh[31044], Fresh[31043], Fresh[31042], Fresh[31041], Fresh[31040], Fresh[31039], Fresh[31038], Fresh[31037], Fresh[31036], Fresh[31035], Fresh[31034], Fresh[31033], Fresh[31032], Fresh[31031], Fresh[31030], Fresh[31029], Fresh[31028], Fresh[31027], Fresh[31026], Fresh[31025], Fresh[31024], Fresh[31023], Fresh[31022], Fresh[31021], Fresh[31020], Fresh[31019], Fresh[31018], Fresh[31017], Fresh[31016], Fresh[31015], Fresh[31014], Fresh[31013], Fresh[31012], Fresh[31011], Fresh[31010], Fresh[31009], Fresh[31008], Fresh[31007], Fresh[31006], Fresh[31005], Fresh[31004], Fresh[31003], Fresh[31002], Fresh[31001], Fresh[31000], Fresh[30999], Fresh[30998], Fresh[30997], Fresh[30996], Fresh[30995], Fresh[30994], Fresh[30993], Fresh[30992], Fresh[30991], Fresh[30990], Fresh[30989], Fresh[30988], Fresh[30987], Fresh[30986], Fresh[30985], Fresh[30984], Fresh[30983], Fresh[30982], Fresh[30981], Fresh[30980], Fresh[30979], Fresh[30978], Fresh[30977], Fresh[30976], Fresh[30975], Fresh[30974], Fresh[30973], Fresh[30972], Fresh[30971], Fresh[30970], Fresh[30969], Fresh[30968], Fresh[30967], Fresh[30966], Fresh[30965], Fresh[30964], Fresh[30963], Fresh[30962], Fresh[30961], Fresh[30960], Fresh[30959], Fresh[30958], Fresh[30957], Fresh[30956], Fresh[30955], Fresh[30954], Fresh[30953], Fresh[30952], Fresh[30951], Fresh[30950], Fresh[30949], Fresh[30948], Fresh[30947], Fresh[30946], Fresh[30945], Fresh[30944], Fresh[30943], Fresh[30942], Fresh[30941], Fresh[30940], Fresh[30939], Fresh[30938], Fresh[30937], Fresh[30936], Fresh[30935], Fresh[30934], Fresh[30933], Fresh[30932], Fresh[30931], Fresh[30930], Fresh[30929], Fresh[30928], Fresh[30927], Fresh[30926], Fresh[30925], Fresh[30924], Fresh[30923], Fresh[30922], Fresh[30921], Fresh[30920], Fresh[30919], Fresh[30918], Fresh[30917], Fresh[30916], Fresh[30915], Fresh[30914], Fresh[30913], Fresh[30912], Fresh[30911], Fresh[30910], Fresh[30909], Fresh[30908], Fresh[30907], Fresh[30906], Fresh[30905], Fresh[30904], Fresh[30903], Fresh[30902], Fresh[30901], Fresh[30900], Fresh[30899], Fresh[30898], Fresh[30897], Fresh[30896], Fresh[30895], Fresh[30894], Fresh[30893], Fresh[30892], Fresh[30891], Fresh[30890], Fresh[30889], Fresh[30888], Fresh[30887], Fresh[30886], Fresh[30885], Fresh[30884], Fresh[30883], Fresh[30882], Fresh[30881], Fresh[30880], Fresh[30879], Fresh[30878], Fresh[30877], Fresh[30876], Fresh[30875], Fresh[30874], Fresh[30873], Fresh[30872], Fresh[30871], Fresh[30870], Fresh[30869], Fresh[30868], Fresh[30867], Fresh[30866], Fresh[30865], Fresh[30864], Fresh[30863], Fresh[30862], Fresh[30861], Fresh[30860], Fresh[30859], Fresh[30858], Fresh[30857], Fresh[30856], Fresh[30855], Fresh[30854], Fresh[30853], Fresh[30852], Fresh[30851], Fresh[30850], Fresh[30849], Fresh[30848], Fresh[30847], Fresh[30846], Fresh[30845], Fresh[30844], Fresh[30843], Fresh[30842], Fresh[30841], Fresh[30840], Fresh[30839], Fresh[30838], Fresh[30837], Fresh[30836], Fresh[30835], Fresh[30834], Fresh[30833], Fresh[30832], Fresh[30831], Fresh[30830], Fresh[30829], Fresh[30828], Fresh[30827], Fresh[30826], Fresh[30825], Fresh[30824], Fresh[30823], Fresh[30822], Fresh[30821], Fresh[30820], Fresh[30819], Fresh[30818], Fresh[30817], Fresh[30816], Fresh[30815], Fresh[30814], Fresh[30813], Fresh[30812], Fresh[30811], Fresh[30810], Fresh[30809], Fresh[30808], Fresh[30807], Fresh[30806], Fresh[30805], Fresh[30804], Fresh[30803], Fresh[30802], Fresh[30801], Fresh[30800], Fresh[30799], Fresh[30798], Fresh[30797], Fresh[30796], Fresh[30795], Fresh[30794], Fresh[30793], Fresh[30792], Fresh[30791], Fresh[30790], Fresh[30789], Fresh[30788], Fresh[30787], Fresh[30786], Fresh[30785], Fresh[30784], Fresh[30783], Fresh[30782], Fresh[30781], Fresh[30780], Fresh[30779], Fresh[30778], Fresh[30777], Fresh[30776], Fresh[30775], Fresh[30774], Fresh[30773], Fresh[30772], Fresh[30771], Fresh[30770], Fresh[30769], Fresh[30768], Fresh[30767], Fresh[30766], Fresh[30765], Fresh[30764], Fresh[30763], Fresh[30762], Fresh[30761], Fresh[30760], Fresh[30759], Fresh[30758], Fresh[30757], Fresh[30756], Fresh[30755], Fresh[30754], Fresh[30753], Fresh[30752], Fresh[30751], Fresh[30750], Fresh[30749], Fresh[30748], Fresh[30747], Fresh[30746], Fresh[30745], Fresh[30744], Fresh[30743], Fresh[30742], Fresh[30741], Fresh[30740], Fresh[30739], Fresh[30738], Fresh[30737], Fresh[30736], Fresh[30735], Fresh[30734], Fresh[30733], Fresh[30732], Fresh[30731], Fresh[30730], Fresh[30729], Fresh[30728], Fresh[30727], Fresh[30726], Fresh[30725], Fresh[30724], Fresh[30723], Fresh[30722], Fresh[30721], Fresh[30720], Fresh[30719], Fresh[30718], Fresh[30717], Fresh[30716], Fresh[30715], Fresh[30714], Fresh[30713], Fresh[30712], Fresh[30711], Fresh[30710], Fresh[30709], Fresh[30708], Fresh[30707], Fresh[30706], Fresh[30705], Fresh[30704], Fresh[30703], Fresh[30702], Fresh[30701], Fresh[30700], Fresh[30699], Fresh[30698], Fresh[30697], Fresh[30696], Fresh[30695], Fresh[30694], Fresh[30693], Fresh[30692], Fresh[30691], Fresh[30690], Fresh[30689], Fresh[30688], Fresh[30687], Fresh[30686], Fresh[30685], Fresh[30684], Fresh[30683], Fresh[30682], Fresh[30681], Fresh[30680], Fresh[30679], Fresh[30678], Fresh[30677], Fresh[30676], Fresh[30675], Fresh[30674], Fresh[30673], Fresh[30672], Fresh[30671], Fresh[30670], Fresh[30669], Fresh[30668], Fresh[30667], Fresh[30666], Fresh[30665], Fresh[30664], Fresh[30663], Fresh[30662], Fresh[30661], Fresh[30660], Fresh[30659], Fresh[30658], Fresh[30657], Fresh[30656], Fresh[30655], Fresh[30654], Fresh[30653], Fresh[30652], Fresh[30651], Fresh[30650], Fresh[30649], Fresh[30648], Fresh[30647], Fresh[30646], Fresh[30645], Fresh[30644], Fresh[30643], Fresh[30642], Fresh[30641], Fresh[30640], Fresh[30639], Fresh[30638], Fresh[30637], Fresh[30636], Fresh[30635], Fresh[30634], Fresh[30633], Fresh[30632], Fresh[30631], Fresh[30630], Fresh[30629], Fresh[30628], Fresh[30627], Fresh[30626], Fresh[30625], Fresh[30624], Fresh[30623], Fresh[30622], Fresh[30621], Fresh[30620], Fresh[30619], Fresh[30618], Fresh[30617], Fresh[30616], Fresh[30615], Fresh[30614], Fresh[30613], Fresh[30612], Fresh[30611], Fresh[30610], Fresh[30609], Fresh[30608], Fresh[30607], Fresh[30606], Fresh[30605], Fresh[30604], Fresh[30603], Fresh[30602], Fresh[30601], Fresh[30600], Fresh[30599], Fresh[30598], Fresh[30597], Fresh[30596], Fresh[30595], Fresh[30594], Fresh[30593], Fresh[30592], Fresh[30591], Fresh[30590], Fresh[30589], Fresh[30588], Fresh[30587], Fresh[30586], Fresh[30585], Fresh[30584], Fresh[30583], Fresh[30582], Fresh[30581], Fresh[30580], Fresh[30579], Fresh[30578], Fresh[30577], Fresh[30576], Fresh[30575], Fresh[30574], Fresh[30573], Fresh[30572], Fresh[30571], Fresh[30570], Fresh[30569], Fresh[30568], Fresh[30567], Fresh[30566], Fresh[30565], Fresh[30564], Fresh[30563], Fresh[30562], Fresh[30561], Fresh[30560], Fresh[30559], Fresh[30558], Fresh[30557], Fresh[30556], Fresh[30555], Fresh[30554], Fresh[30553], Fresh[30552], Fresh[30551], Fresh[30550], Fresh[30549], Fresh[30548], Fresh[30547], Fresh[30546], Fresh[30545], Fresh[30544], Fresh[30543], Fresh[30542], Fresh[30541], Fresh[30540], Fresh[30539], Fresh[30538], Fresh[30537], Fresh[30536], Fresh[30535], Fresh[30534], Fresh[30533], Fresh[30532], Fresh[30531], Fresh[30530], Fresh[30529], Fresh[30528], Fresh[30527], Fresh[30526], Fresh[30525], Fresh[30524], Fresh[30523], Fresh[30522], Fresh[30521], Fresh[30520], Fresh[30519], Fresh[30518], Fresh[30517], Fresh[30516], Fresh[30515], Fresh[30514], Fresh[30513], Fresh[30512], Fresh[30511], Fresh[30510], Fresh[30509], Fresh[30508], Fresh[30507], Fresh[30506], Fresh[30505], Fresh[30504], Fresh[30503], Fresh[30502], Fresh[30501], Fresh[30500], Fresh[30499], Fresh[30498], Fresh[30497], Fresh[30496], Fresh[30495], Fresh[30494], Fresh[30493], Fresh[30492], Fresh[30491], Fresh[30490], Fresh[30489], Fresh[30488], Fresh[30487], Fresh[30486], Fresh[30485], Fresh[30484], Fresh[30483], Fresh[30482], Fresh[30481], Fresh[30480], Fresh[30479], Fresh[30478], Fresh[30477], Fresh[30476], Fresh[30475], Fresh[30474], Fresh[30473], Fresh[30472], Fresh[30471], Fresh[30470], Fresh[30469], Fresh[30468], Fresh[30467], Fresh[30466], Fresh[30465], Fresh[30464], Fresh[30463], Fresh[30462], Fresh[30461], Fresh[30460], Fresh[30459], Fresh[30458], Fresh[30457], Fresh[30456], Fresh[30455], Fresh[30454], Fresh[30453], Fresh[30452], Fresh[30451], Fresh[30450], Fresh[30449], Fresh[30448], Fresh[30447], Fresh[30446], Fresh[30445], Fresh[30444], Fresh[30443], Fresh[30442], Fresh[30441], Fresh[30440], Fresh[30439], Fresh[30438], Fresh[30437], Fresh[30436], Fresh[30435], Fresh[30434], Fresh[30433], Fresh[30432], Fresh[30431], Fresh[30430], Fresh[30429], Fresh[30428], Fresh[30427], Fresh[30426], Fresh[30425], Fresh[30424], Fresh[30423], Fresh[30422], Fresh[30421], Fresh[30420], Fresh[30419], Fresh[30418], Fresh[30417], Fresh[30416], Fresh[30415], Fresh[30414], Fresh[30413], Fresh[30412], Fresh[30411], Fresh[30410], Fresh[30409], Fresh[30408], Fresh[30407], Fresh[30406], Fresh[30405], Fresh[30404], Fresh[30403], Fresh[30402], Fresh[30401], Fresh[30400], Fresh[30399], Fresh[30398], Fresh[30397], Fresh[30396], Fresh[30395], Fresh[30394], Fresh[30393], Fresh[30392], Fresh[30391], Fresh[30390], Fresh[30389], Fresh[30388], Fresh[30387], Fresh[30386], Fresh[30385], Fresh[30384], Fresh[30383], Fresh[30382], Fresh[30381], Fresh[30380], Fresh[30379], Fresh[30378], Fresh[30377], Fresh[30376], Fresh[30375], Fresh[30374], Fresh[30373], Fresh[30372], Fresh[30371], Fresh[30370], Fresh[30369], Fresh[30368], Fresh[30367], Fresh[30366], Fresh[30365], Fresh[30364], Fresh[30363], Fresh[30362], Fresh[30361], Fresh[30360], Fresh[30359], Fresh[30358], Fresh[30357], Fresh[30356], Fresh[30355], Fresh[30354], Fresh[30353], Fresh[30352], Fresh[30351], Fresh[30350], Fresh[30349], Fresh[30348], Fresh[30347], Fresh[30346], Fresh[30345], Fresh[30344], Fresh[30343], Fresh[30342], Fresh[30341], Fresh[30340], Fresh[30339], Fresh[30338], Fresh[30337], Fresh[30336], Fresh[30335], Fresh[30334], Fresh[30333], Fresh[30332], Fresh[30331], Fresh[30330], Fresh[30329], Fresh[30328], Fresh[30327], Fresh[30326], Fresh[30325], Fresh[30324], Fresh[30323], Fresh[30322], Fresh[30321], Fresh[30320], Fresh[30319], Fresh[30318], Fresh[30317], Fresh[30316], Fresh[30315], Fresh[30314], Fresh[30313], Fresh[30312], Fresh[30311], Fresh[30310], Fresh[30309], Fresh[30308], Fresh[30307], Fresh[30306], Fresh[30305], Fresh[30304], Fresh[30303], Fresh[30302], Fresh[30301], Fresh[30300], Fresh[30299], Fresh[30298], Fresh[30297], Fresh[30296], Fresh[30295], Fresh[30294], Fresh[30293], Fresh[30292], Fresh[30291], Fresh[30290], Fresh[30289], Fresh[30288], Fresh[30287], Fresh[30286], Fresh[30285], Fresh[30284], Fresh[30283], Fresh[30282], Fresh[30281], Fresh[30280], Fresh[30279], Fresh[30278], Fresh[30277], Fresh[30276], Fresh[30275], Fresh[30274], Fresh[30273], Fresh[30272], Fresh[30271], Fresh[30270], Fresh[30269], Fresh[30268], Fresh[30267], Fresh[30266], Fresh[30265], Fresh[30264], Fresh[30263], Fresh[30262], Fresh[30261], Fresh[30260], Fresh[30259], Fresh[30258], Fresh[30257], Fresh[30256], Fresh[30255], Fresh[30254], Fresh[30253], Fresh[30252], Fresh[30251], Fresh[30250], Fresh[30249], Fresh[30248], Fresh[30247], Fresh[30246], Fresh[30245], Fresh[30244], Fresh[30243], Fresh[30242], Fresh[30241], Fresh[30240], Fresh[30239], Fresh[30238], Fresh[30237], Fresh[30236], Fresh[30235], Fresh[30234], Fresh[30233], Fresh[30232], Fresh[30231], Fresh[30230], Fresh[30229], Fresh[30228], Fresh[30227], Fresh[30226], Fresh[30225], Fresh[30224], Fresh[30223], Fresh[30222], Fresh[30221], Fresh[30220], Fresh[30219], Fresh[30218], Fresh[30217], Fresh[30216], Fresh[30215], Fresh[30214], Fresh[30213], Fresh[30212], Fresh[30211], Fresh[30210], Fresh[30209], Fresh[30208], Fresh[30207], Fresh[30206], Fresh[30205], Fresh[30204], Fresh[30203], Fresh[30202], Fresh[30201], Fresh[30200], Fresh[30199], Fresh[30198], Fresh[30197], Fresh[30196], Fresh[30195], Fresh[30194], Fresh[30193], Fresh[30192], Fresh[30191], Fresh[30190], Fresh[30189], Fresh[30188], Fresh[30187], Fresh[30186], Fresh[30185], Fresh[30184], Fresh[30183], Fresh[30182], Fresh[30181], Fresh[30180], Fresh[30179], Fresh[30178], Fresh[30177], Fresh[30176], Fresh[30175], Fresh[30174], Fresh[30173], Fresh[30172], Fresh[30171], Fresh[30170], Fresh[30169], Fresh[30168], Fresh[30167], Fresh[30166], Fresh[30165], Fresh[30164], Fresh[30163], Fresh[30162], Fresh[30161], Fresh[30160], Fresh[30159], Fresh[30158], Fresh[30157], Fresh[30156], Fresh[30155], Fresh[30154], Fresh[30153], Fresh[30152], Fresh[30151], Fresh[30150], Fresh[30149], Fresh[30148], Fresh[30147], Fresh[30146], Fresh[30145], Fresh[30144], Fresh[30143], Fresh[30142], Fresh[30141], Fresh[30140], Fresh[30139], Fresh[30138], Fresh[30137], Fresh[30136], Fresh[30135], Fresh[30134], Fresh[30133], Fresh[30132], Fresh[30131], Fresh[30130], Fresh[30129], Fresh[30128], Fresh[30127], Fresh[30126], Fresh[30125], Fresh[30124], Fresh[30123], Fresh[30122], Fresh[30121], Fresh[30120], Fresh[30119], Fresh[30118], Fresh[30117], Fresh[30116], Fresh[30115], Fresh[30114], Fresh[30113], Fresh[30112], Fresh[30111], Fresh[30110], Fresh[30109], Fresh[30108], Fresh[30107], Fresh[30106], Fresh[30105], Fresh[30104], Fresh[30103], Fresh[30102], Fresh[30101], Fresh[30100], Fresh[30099], Fresh[30098], Fresh[30097], Fresh[30096], Fresh[30095], Fresh[30094], Fresh[30093], Fresh[30092], Fresh[30091], Fresh[30090], Fresh[30089], Fresh[30088], Fresh[30087], Fresh[30086], Fresh[30085], Fresh[30084], Fresh[30083], Fresh[30082], Fresh[30081], Fresh[30080], Fresh[30079], Fresh[30078], Fresh[30077], Fresh[30076], Fresh[30075], Fresh[30074], Fresh[30073], Fresh[30072], Fresh[30071], Fresh[30070], Fresh[30069], Fresh[30068], Fresh[30067], Fresh[30066], Fresh[30065], Fresh[30064], Fresh[30063], Fresh[30062], Fresh[30061], Fresh[30060], Fresh[30059], Fresh[30058], Fresh[30057], Fresh[30056], Fresh[30055], Fresh[30054], Fresh[30053], Fresh[30052], Fresh[30051], Fresh[30050], Fresh[30049], Fresh[30048], Fresh[30047], Fresh[30046], Fresh[30045], Fresh[30044], Fresh[30043], Fresh[30042], Fresh[30041], Fresh[30040], Fresh[30039], Fresh[30038], Fresh[30037], Fresh[30036], Fresh[30035], Fresh[30034], Fresh[30033], Fresh[30032], Fresh[30031], Fresh[30030], Fresh[30029], Fresh[30028], Fresh[30027], Fresh[30026], Fresh[30025], Fresh[30024], Fresh[30023], Fresh[30022], Fresh[30021], Fresh[30020], Fresh[30019], Fresh[30018], Fresh[30017], Fresh[30016], Fresh[30015], Fresh[30014], Fresh[30013], Fresh[30012], Fresh[30011], Fresh[30010], Fresh[30009], Fresh[30008], Fresh[30007], Fresh[30006], Fresh[30005], Fresh[30004], Fresh[30003], Fresh[30002], Fresh[30001], Fresh[30000], Fresh[29999], Fresh[29998], Fresh[29997], Fresh[29996], Fresh[29995], Fresh[29994], Fresh[29993], Fresh[29992], Fresh[29991], Fresh[29990], Fresh[29989], Fresh[29988], Fresh[29987], Fresh[29986], Fresh[29985], Fresh[29984], Fresh[29983], Fresh[29982], Fresh[29981], Fresh[29980], Fresh[29979], Fresh[29978], Fresh[29977], Fresh[29976], Fresh[29975], Fresh[29974], Fresh[29973], Fresh[29972], Fresh[29971], Fresh[29970], Fresh[29969], Fresh[29968], Fresh[29967], Fresh[29966], Fresh[29965], Fresh[29964], Fresh[29963], Fresh[29962], Fresh[29961], Fresh[29960], Fresh[29959], Fresh[29958], Fresh[29957], Fresh[29956], Fresh[29955], Fresh[29954], Fresh[29953], Fresh[29952], Fresh[29951], Fresh[29950], Fresh[29949], Fresh[29948], Fresh[29947], Fresh[29946], Fresh[29945], Fresh[29944], Fresh[29943], Fresh[29942], Fresh[29941], Fresh[29940], Fresh[29939], Fresh[29938], Fresh[29937], Fresh[29936], Fresh[29935], Fresh[29934], Fresh[29933], Fresh[29932], Fresh[29931], Fresh[29930], Fresh[29929], Fresh[29928], Fresh[29927], Fresh[29926], Fresh[29925], Fresh[29924], Fresh[29923], Fresh[29922], Fresh[29921], Fresh[29920], Fresh[29919], Fresh[29918], Fresh[29917], Fresh[29916], Fresh[29915], Fresh[29914], Fresh[29913], Fresh[29912], Fresh[29911], Fresh[29910], Fresh[29909], Fresh[29908], Fresh[29907], Fresh[29906], Fresh[29905], Fresh[29904], Fresh[29903], Fresh[29902], Fresh[29901], Fresh[29900], Fresh[29899], Fresh[29898], Fresh[29897], Fresh[29896], Fresh[29895], Fresh[29894], Fresh[29893], Fresh[29892], Fresh[29891], Fresh[29890], Fresh[29889], Fresh[29888], Fresh[29887], Fresh[29886], Fresh[29885], Fresh[29884], Fresh[29883], Fresh[29882], Fresh[29881], Fresh[29880], Fresh[29879], Fresh[29878], Fresh[29877], Fresh[29876], Fresh[29875], Fresh[29874], Fresh[29873], Fresh[29872], Fresh[29871], Fresh[29870], Fresh[29869], Fresh[29868], Fresh[29867], Fresh[29866], Fresh[29865], Fresh[29864], Fresh[29863], Fresh[29862], Fresh[29861], Fresh[29860], Fresh[29859], Fresh[29858], Fresh[29857], Fresh[29856], Fresh[29855], Fresh[29854], Fresh[29853], Fresh[29852], Fresh[29851], Fresh[29850], Fresh[29849], Fresh[29848], Fresh[29847], Fresh[29846], Fresh[29845], Fresh[29844], Fresh[29843], Fresh[29842], Fresh[29841], Fresh[29840], Fresh[29839], Fresh[29838], Fresh[29837], Fresh[29836], Fresh[29835], Fresh[29834], Fresh[29833], Fresh[29832], Fresh[29831], Fresh[29830], Fresh[29829], Fresh[29828], Fresh[29827], Fresh[29826], Fresh[29825], Fresh[29824], Fresh[29823], Fresh[29822], Fresh[29821], Fresh[29820], Fresh[29819], Fresh[29818], Fresh[29817], Fresh[29816], Fresh[29815], Fresh[29814], Fresh[29813], Fresh[29812], Fresh[29811], Fresh[29810], Fresh[29809], Fresh[29808], Fresh[29807], Fresh[29806], Fresh[29805], Fresh[29804], Fresh[29803], Fresh[29802], Fresh[29801], Fresh[29800], Fresh[29799], Fresh[29798], Fresh[29797], Fresh[29796], Fresh[29795], Fresh[29794], Fresh[29793], Fresh[29792], Fresh[29791], Fresh[29790], Fresh[29789], Fresh[29788], Fresh[29787], Fresh[29786], Fresh[29785], Fresh[29784], Fresh[29783], Fresh[29782], Fresh[29781], Fresh[29780], Fresh[29779], Fresh[29778], Fresh[29777], Fresh[29776], Fresh[29775], Fresh[29774], Fresh[29773], Fresh[29772], Fresh[29771], Fresh[29770], Fresh[29769], Fresh[29768], Fresh[29767], Fresh[29766], Fresh[29765], Fresh[29764], Fresh[29763], Fresh[29762], Fresh[29761], Fresh[29760], Fresh[29759], Fresh[29758], Fresh[29757], Fresh[29756], Fresh[29755], Fresh[29754], Fresh[29753], Fresh[29752], Fresh[29751], Fresh[29750], Fresh[29749], Fresh[29748], Fresh[29747], Fresh[29746], Fresh[29745], Fresh[29744], Fresh[29743], Fresh[29742], Fresh[29741], Fresh[29740], Fresh[29739], Fresh[29738], Fresh[29737], Fresh[29736], Fresh[29735], Fresh[29734], Fresh[29733], Fresh[29732], Fresh[29731], Fresh[29730], Fresh[29729], Fresh[29728], Fresh[29727], Fresh[29726], Fresh[29725], Fresh[29724], Fresh[29723], Fresh[29722], Fresh[29721], Fresh[29720], Fresh[29719], Fresh[29718], Fresh[29717], Fresh[29716], Fresh[29715], Fresh[29714], Fresh[29713], Fresh[29712], Fresh[29711], Fresh[29710], Fresh[29709], Fresh[29708], Fresh[29707], Fresh[29706], Fresh[29705], Fresh[29704], Fresh[29703], Fresh[29702], Fresh[29701], Fresh[29700], Fresh[29699], Fresh[29698], Fresh[29697], Fresh[29696], Fresh[29695], Fresh[29694], Fresh[29693], Fresh[29692], Fresh[29691], Fresh[29690], Fresh[29689], Fresh[29688], Fresh[29687], Fresh[29686], Fresh[29685], Fresh[29684], Fresh[29683], Fresh[29682], Fresh[29681], Fresh[29680], Fresh[29679], Fresh[29678], Fresh[29677], Fresh[29676], Fresh[29675], Fresh[29674], Fresh[29673], Fresh[29672], Fresh[29671], Fresh[29670], Fresh[29669], Fresh[29668], Fresh[29667], Fresh[29666], Fresh[29665], Fresh[29664], Fresh[29663], Fresh[29662], Fresh[29661], Fresh[29660], Fresh[29659], Fresh[29658], Fresh[29657], Fresh[29656], Fresh[29655], Fresh[29654], Fresh[29653], Fresh[29652], Fresh[29651], Fresh[29650], Fresh[29649], Fresh[29648], Fresh[29647], Fresh[29646], Fresh[29645], Fresh[29644], Fresh[29643], Fresh[29642], Fresh[29641], Fresh[29640], Fresh[29639], Fresh[29638], Fresh[29637], Fresh[29636], Fresh[29635], Fresh[29634], Fresh[29633], Fresh[29632], Fresh[29631], Fresh[29630], Fresh[29629], Fresh[29628], Fresh[29627], Fresh[29626], Fresh[29625], Fresh[29624], Fresh[29623], Fresh[29622], Fresh[29621], Fresh[29620], Fresh[29619], Fresh[29618], Fresh[29617], Fresh[29616], Fresh[29615], Fresh[29614], Fresh[29613], Fresh[29612], Fresh[29611], Fresh[29610], Fresh[29609], Fresh[29608], Fresh[29607], Fresh[29606], Fresh[29605], Fresh[29604], Fresh[29603], Fresh[29602], Fresh[29601], Fresh[29600], Fresh[29599], Fresh[29598], Fresh[29597], Fresh[29596], Fresh[29595], Fresh[29594], Fresh[29593], Fresh[29592], Fresh[29591], Fresh[29590], Fresh[29589], Fresh[29588], Fresh[29587], Fresh[29586], Fresh[29585], Fresh[29584], Fresh[29583], Fresh[29582], Fresh[29581], Fresh[29580], Fresh[29579], Fresh[29578], Fresh[29577], Fresh[29576], Fresh[29575], Fresh[29574], Fresh[29573], Fresh[29572], Fresh[29571], Fresh[29570], Fresh[29569], Fresh[29568], Fresh[29567], Fresh[29566], Fresh[29565], Fresh[29564], Fresh[29563], Fresh[29562], Fresh[29561], Fresh[29560], Fresh[29559], Fresh[29558], Fresh[29557], Fresh[29556], Fresh[29555], Fresh[29554], Fresh[29553], Fresh[29552], Fresh[29551], Fresh[29550], Fresh[29549], Fresh[29548], Fresh[29547], Fresh[29546], Fresh[29545], Fresh[29544], Fresh[29543], Fresh[29542], Fresh[29541], Fresh[29540], Fresh[29539], Fresh[29538], Fresh[29537], Fresh[29536], Fresh[29535], Fresh[29534], Fresh[29533], Fresh[29532], Fresh[29531], Fresh[29530], Fresh[29529], Fresh[29528], Fresh[29527], Fresh[29526], Fresh[29525], Fresh[29524], Fresh[29523], Fresh[29522], Fresh[29521], Fresh[29520], Fresh[29519], Fresh[29518], Fresh[29517], Fresh[29516], Fresh[29515], Fresh[29514], Fresh[29513], Fresh[29512], Fresh[29511], Fresh[29510], Fresh[29509], Fresh[29508], Fresh[29507], Fresh[29506], Fresh[29505], Fresh[29504], Fresh[29503], Fresh[29502], Fresh[29501], Fresh[29500], Fresh[29499], Fresh[29498], Fresh[29497], Fresh[29496], Fresh[29495], Fresh[29494], Fresh[29493], Fresh[29492], Fresh[29491], Fresh[29490], Fresh[29489], Fresh[29488], Fresh[29487], Fresh[29486], Fresh[29485], Fresh[29484], Fresh[29483], Fresh[29482], Fresh[29481], Fresh[29480], Fresh[29479], Fresh[29478], Fresh[29477], Fresh[29476], Fresh[29475], Fresh[29474], Fresh[29473], Fresh[29472], Fresh[29471], Fresh[29470], Fresh[29469], Fresh[29468], Fresh[29467], Fresh[29466], Fresh[29465], Fresh[29464], Fresh[29463], Fresh[29462], Fresh[29461], Fresh[29460], Fresh[29459], Fresh[29458], Fresh[29457], Fresh[29456], Fresh[29455], Fresh[29454], Fresh[29453], Fresh[29452], Fresh[29451], Fresh[29450], Fresh[29449], Fresh[29448], Fresh[29447], Fresh[29446], Fresh[29445], Fresh[29444], Fresh[29443], Fresh[29442], Fresh[29441], Fresh[29440], Fresh[29439], Fresh[29438], Fresh[29437], Fresh[29436], Fresh[29435], Fresh[29434], Fresh[29433], Fresh[29432], Fresh[29431], Fresh[29430], Fresh[29429], Fresh[29428], Fresh[29427], Fresh[29426], Fresh[29425], Fresh[29424], Fresh[29423], Fresh[29422], Fresh[29421], Fresh[29420], Fresh[29419], Fresh[29418], Fresh[29417], Fresh[29416], Fresh[29415], Fresh[29414], Fresh[29413], Fresh[29412], Fresh[29411], Fresh[29410], Fresh[29409], Fresh[29408], Fresh[29407], Fresh[29406], Fresh[29405], Fresh[29404], Fresh[29403], Fresh[29402], Fresh[29401], Fresh[29400], Fresh[29399], Fresh[29398], Fresh[29397], Fresh[29396], Fresh[29395], Fresh[29394], Fresh[29393], Fresh[29392], Fresh[29391], Fresh[29390], Fresh[29389], Fresh[29388], Fresh[29387], Fresh[29386], Fresh[29385], Fresh[29384], Fresh[29383], Fresh[29382], Fresh[29381], Fresh[29380], Fresh[29379], Fresh[29378], Fresh[29377], Fresh[29376], Fresh[29375], Fresh[29374], Fresh[29373], Fresh[29372], Fresh[29371], Fresh[29370], Fresh[29369], Fresh[29368], Fresh[29367], Fresh[29366], Fresh[29365], Fresh[29364], Fresh[29363], Fresh[29362], Fresh[29361], Fresh[29360], Fresh[29359], Fresh[29358], Fresh[29357], Fresh[29356], Fresh[29355], Fresh[29354], Fresh[29353], Fresh[29352], Fresh[29351], Fresh[29350], Fresh[29349], Fresh[29348], Fresh[29347], Fresh[29346], Fresh[29345], Fresh[29344], Fresh[29343], Fresh[29342], Fresh[29341], Fresh[29340], Fresh[29339], Fresh[29338], Fresh[29337], Fresh[29336], Fresh[29335], Fresh[29334], Fresh[29333], Fresh[29332], Fresh[29331], Fresh[29330], Fresh[29329], Fresh[29328], Fresh[29327], Fresh[29326], Fresh[29325], Fresh[29324], Fresh[29323], Fresh[29322], Fresh[29321], Fresh[29320], Fresh[29319], Fresh[29318], Fresh[29317], Fresh[29316], Fresh[29315], Fresh[29314], Fresh[29313], Fresh[29312], Fresh[29311], Fresh[29310], Fresh[29309], Fresh[29308], Fresh[29307], Fresh[29306], Fresh[29305], Fresh[29304], Fresh[29303], Fresh[29302], Fresh[29301], Fresh[29300], Fresh[29299], Fresh[29298], Fresh[29297], Fresh[29296], Fresh[29295], Fresh[29294], Fresh[29293], Fresh[29292], Fresh[29291], Fresh[29290], Fresh[29289], Fresh[29288], Fresh[29287], Fresh[29286], Fresh[29285], Fresh[29284], Fresh[29283], Fresh[29282], Fresh[29281], Fresh[29280], Fresh[29279], Fresh[29278], Fresh[29277], Fresh[29276], Fresh[29275], Fresh[29274], Fresh[29273], Fresh[29272], Fresh[29271], Fresh[29270], Fresh[29269], Fresh[29268], Fresh[29267], Fresh[29266], Fresh[29265], Fresh[29264], Fresh[29263], Fresh[29262], Fresh[29261], Fresh[29260], Fresh[29259], Fresh[29258], Fresh[29257], Fresh[29256], Fresh[29255], Fresh[29254], Fresh[29253], Fresh[29252], Fresh[29251], Fresh[29250], Fresh[29249], Fresh[29248], Fresh[29247], Fresh[29246], Fresh[29245], Fresh[29244], Fresh[29243], Fresh[29242], Fresh[29241], Fresh[29240], Fresh[29239], Fresh[29238], Fresh[29237], Fresh[29236], Fresh[29235], Fresh[29234], Fresh[29233], Fresh[29232], Fresh[29231], Fresh[29230], Fresh[29229], Fresh[29228], Fresh[29227], Fresh[29226], Fresh[29225], Fresh[29224], Fresh[29223], Fresh[29222], Fresh[29221], Fresh[29220], Fresh[29219], Fresh[29218], Fresh[29217], Fresh[29216], Fresh[29215], Fresh[29214], Fresh[29213], Fresh[29212], Fresh[29211], Fresh[29210], Fresh[29209], Fresh[29208], Fresh[29207], Fresh[29206], Fresh[29205], Fresh[29204], Fresh[29203], Fresh[29202], Fresh[29201], Fresh[29200], Fresh[29199], Fresh[29198], Fresh[29197], Fresh[29196], Fresh[29195], Fresh[29194], Fresh[29193], Fresh[29192], Fresh[29191], Fresh[29190], Fresh[29189], Fresh[29188], Fresh[29187], Fresh[29186], Fresh[29185], Fresh[29184], Fresh[29183], Fresh[29182], Fresh[29181], Fresh[29180], Fresh[29179], Fresh[29178], Fresh[29177], Fresh[29176], Fresh[29175], Fresh[29174], Fresh[29173], Fresh[29172], Fresh[29171], Fresh[29170], Fresh[29169], Fresh[29168], Fresh[29167], Fresh[29166], Fresh[29165], Fresh[29164], Fresh[29163], Fresh[29162], Fresh[29161], Fresh[29160], Fresh[29159], Fresh[29158], Fresh[29157], Fresh[29156], Fresh[29155], Fresh[29154], Fresh[29153], Fresh[29152], Fresh[29151], Fresh[29150], Fresh[29149], Fresh[29148], Fresh[29147], Fresh[29146], Fresh[29145], Fresh[29144], Fresh[29143], Fresh[29142], Fresh[29141], Fresh[29140], Fresh[29139], Fresh[29138], Fresh[29137], Fresh[29136], Fresh[29135], Fresh[29134], Fresh[29133], Fresh[29132], Fresh[29131], Fresh[29130], Fresh[29129], Fresh[29128], Fresh[29127], Fresh[29126], Fresh[29125], Fresh[29124], Fresh[29123], Fresh[29122], Fresh[29121], Fresh[29120], Fresh[29119], Fresh[29118], Fresh[29117], Fresh[29116], Fresh[29115], Fresh[29114], Fresh[29113], Fresh[29112], Fresh[29111], Fresh[29110], Fresh[29109], Fresh[29108], Fresh[29107], Fresh[29106], Fresh[29105], Fresh[29104], Fresh[29103], Fresh[29102], Fresh[29101], Fresh[29100], Fresh[29099], Fresh[29098], Fresh[29097], Fresh[29096], Fresh[29095], Fresh[29094], Fresh[29093], Fresh[29092], Fresh[29091], Fresh[29090], Fresh[29089], Fresh[29088], Fresh[29087], Fresh[29086], Fresh[29085], Fresh[29084], Fresh[29083], Fresh[29082], Fresh[29081], Fresh[29080], Fresh[29079], Fresh[29078], Fresh[29077], Fresh[29076], Fresh[29075], Fresh[29074], Fresh[29073], Fresh[29072], Fresh[29071], Fresh[29070], Fresh[29069], Fresh[29068], Fresh[29067], Fresh[29066], Fresh[29065], Fresh[29064], Fresh[29063], Fresh[29062], Fresh[29061], Fresh[29060], Fresh[29059], Fresh[29058], Fresh[29057], Fresh[29056], Fresh[29055], Fresh[29054], Fresh[29053], Fresh[29052], Fresh[29051], Fresh[29050], Fresh[29049], Fresh[29048], Fresh[29047], Fresh[29046], Fresh[29045], Fresh[29044], Fresh[29043], Fresh[29042], Fresh[29041], Fresh[29040], Fresh[29039], Fresh[29038], Fresh[29037], Fresh[29036], Fresh[29035], Fresh[29034], Fresh[29033], Fresh[29032], Fresh[29031], Fresh[29030], Fresh[29029], Fresh[29028], Fresh[29027], Fresh[29026], Fresh[29025], Fresh[29024], Fresh[29023], Fresh[29022], Fresh[29021], Fresh[29020], Fresh[29019], Fresh[29018], Fresh[29017], Fresh[29016], Fresh[29015], Fresh[29014], Fresh[29013], Fresh[29012], Fresh[29011], Fresh[29010], Fresh[29009], Fresh[29008], Fresh[29007], Fresh[29006], Fresh[29005], Fresh[29004], Fresh[29003], Fresh[29002], Fresh[29001], Fresh[29000], Fresh[28999], Fresh[28998], Fresh[28997], Fresh[28996], Fresh[28995], Fresh[28994], Fresh[28993], Fresh[28992], Fresh[28991], Fresh[28990], Fresh[28989], Fresh[28988], Fresh[28987], Fresh[28986], Fresh[28985], Fresh[28984], Fresh[28983], Fresh[28982], Fresh[28981], Fresh[28980], Fresh[28979], Fresh[28978], Fresh[28977], Fresh[28976], Fresh[28975], Fresh[28974], Fresh[28973], Fresh[28972], Fresh[28971], Fresh[28970], Fresh[28969], Fresh[28968], Fresh[28967], Fresh[28966], Fresh[28965], Fresh[28964], Fresh[28963], Fresh[28962], Fresh[28961], Fresh[28960], Fresh[28959], Fresh[28958], Fresh[28957], Fresh[28956], Fresh[28955], Fresh[28954], Fresh[28953], Fresh[28952], Fresh[28951], Fresh[28950], Fresh[28949], Fresh[28948], Fresh[28947], Fresh[28946], Fresh[28945], Fresh[28944], Fresh[28943], Fresh[28942], Fresh[28941], Fresh[28940], Fresh[28939], Fresh[28938], Fresh[28937], Fresh[28936], Fresh[28935], Fresh[28934], Fresh[28933], Fresh[28932], Fresh[28931], Fresh[28930], Fresh[28929], Fresh[28928], Fresh[28927], Fresh[28926], Fresh[28925], Fresh[28924], Fresh[28923], Fresh[28922], Fresh[28921], Fresh[28920], Fresh[28919], Fresh[28918], Fresh[28917], Fresh[28916], Fresh[28915], Fresh[28914], Fresh[28913], Fresh[28912], Fresh[28911], Fresh[28910], Fresh[28909], Fresh[28908], Fresh[28907], Fresh[28906], Fresh[28905], Fresh[28904], Fresh[28903], Fresh[28902], Fresh[28901], Fresh[28900], Fresh[28899], Fresh[28898], Fresh[28897], Fresh[28896], Fresh[28895], Fresh[28894], Fresh[28893], Fresh[28892], Fresh[28891], Fresh[28890], Fresh[28889], Fresh[28888], Fresh[28887], Fresh[28886], Fresh[28885], Fresh[28884], Fresh[28883], Fresh[28882], Fresh[28881], Fresh[28880], Fresh[28879], Fresh[28878], Fresh[28877], Fresh[28876], Fresh[28875], Fresh[28874], Fresh[28873], Fresh[28872], Fresh[28871], Fresh[28870], Fresh[28869], Fresh[28868], Fresh[28867], Fresh[28866], Fresh[28865], Fresh[28864], Fresh[28863], Fresh[28862], Fresh[28861], Fresh[28860], Fresh[28859], Fresh[28858], Fresh[28857], Fresh[28856], Fresh[28855], Fresh[28854], Fresh[28853], Fresh[28852], Fresh[28851], Fresh[28850], Fresh[28849], Fresh[28848], Fresh[28847], Fresh[28846], Fresh[28845], Fresh[28844], Fresh[28843], Fresh[28842], Fresh[28841], Fresh[28840], Fresh[28839], Fresh[28838], Fresh[28837], Fresh[28836], Fresh[28835], Fresh[28834], Fresh[28833], Fresh[28832], Fresh[28831], Fresh[28830], Fresh[28829], Fresh[28828], Fresh[28827], Fresh[28826], Fresh[28825], Fresh[28824], Fresh[28823], Fresh[28822], Fresh[28821], Fresh[28820], Fresh[28819], Fresh[28818], Fresh[28817], Fresh[28816], Fresh[28815], Fresh[28814], Fresh[28813], Fresh[28812], Fresh[28811], Fresh[28810], Fresh[28809], Fresh[28808], Fresh[28807], Fresh[28806], Fresh[28805], Fresh[28804], Fresh[28803], Fresh[28802], Fresh[28801], Fresh[28800], Fresh[28799], Fresh[28798], Fresh[28797], Fresh[28796], Fresh[28795], Fresh[28794], Fresh[28793], Fresh[28792], Fresh[28791], Fresh[28790], Fresh[28789], Fresh[28788], Fresh[28787], Fresh[28786], Fresh[28785], Fresh[28784], Fresh[28783], Fresh[28782], Fresh[28781], Fresh[28780], Fresh[28779], Fresh[28778], Fresh[28777], Fresh[28776], Fresh[28775], Fresh[28774], Fresh[28773], Fresh[28772], Fresh[28771], Fresh[28770], Fresh[28769], Fresh[28768], Fresh[28767], Fresh[28766], Fresh[28765], Fresh[28764], Fresh[28763], Fresh[28762], Fresh[28761], Fresh[28760], Fresh[28759], Fresh[28758], Fresh[28757], Fresh[28756], Fresh[28755], Fresh[28754], Fresh[28753], Fresh[28752], Fresh[28751], Fresh[28750], Fresh[28749], Fresh[28748], Fresh[28747], Fresh[28746], Fresh[28745], Fresh[28744], Fresh[28743], Fresh[28742], Fresh[28741], Fresh[28740], Fresh[28739], Fresh[28738], Fresh[28737], Fresh[28736], Fresh[28735], Fresh[28734], Fresh[28733], Fresh[28732], Fresh[28731], Fresh[28730], Fresh[28729], Fresh[28728], Fresh[28727], Fresh[28726], Fresh[28725], Fresh[28724], Fresh[28723], Fresh[28722], Fresh[28721], Fresh[28720], Fresh[28719], Fresh[28718], Fresh[28717], Fresh[28716], Fresh[28715], Fresh[28714], Fresh[28713], Fresh[28712], Fresh[28711], Fresh[28710], Fresh[28709], Fresh[28708], Fresh[28707], Fresh[28706], Fresh[28705], Fresh[28704], Fresh[28703], Fresh[28702], Fresh[28701], Fresh[28700], Fresh[28699], Fresh[28698], Fresh[28697], Fresh[28696], Fresh[28695], Fresh[28694], Fresh[28693], Fresh[28692], Fresh[28691], Fresh[28690], Fresh[28689], Fresh[28688], Fresh[28687], Fresh[28686], Fresh[28685], Fresh[28684], Fresh[28683], Fresh[28682], Fresh[28681], Fresh[28680], Fresh[28679], Fresh[28678], Fresh[28677], Fresh[28676], Fresh[28675], Fresh[28674], Fresh[28673], Fresh[28672], Fresh[28671], Fresh[28670], Fresh[28669], Fresh[28668], Fresh[28667], Fresh[28666], Fresh[28665], Fresh[28664], Fresh[28663], Fresh[28662], Fresh[28661], Fresh[28660], Fresh[28659], Fresh[28658], Fresh[28657], Fresh[28656], Fresh[28655], Fresh[28654], Fresh[28653], Fresh[28652], Fresh[28651], Fresh[28650], Fresh[28649], Fresh[28648], Fresh[28647], Fresh[28646], Fresh[28645], Fresh[28644], Fresh[28643], Fresh[28642], Fresh[28641], Fresh[28640], Fresh[28639], Fresh[28638], Fresh[28637], Fresh[28636], Fresh[28635], Fresh[28634], Fresh[28633], Fresh[28632], Fresh[28631], Fresh[28630], Fresh[28629], Fresh[28628], Fresh[28627], Fresh[28626], Fresh[28625], Fresh[28624], Fresh[28623], Fresh[28622], Fresh[28621], Fresh[28620], Fresh[28619], Fresh[28618], Fresh[28617], Fresh[28616], Fresh[28615], Fresh[28614], Fresh[28613], Fresh[28612], Fresh[28611], Fresh[28610], Fresh[28609], Fresh[28608], Fresh[28607], Fresh[28606], Fresh[28605], Fresh[28604], Fresh[28603], Fresh[28602], Fresh[28601], Fresh[28600], Fresh[28599], Fresh[28598], Fresh[28597], Fresh[28596], Fresh[28595], Fresh[28594], Fresh[28593], Fresh[28592], Fresh[28591], Fresh[28590], Fresh[28589], Fresh[28588], Fresh[28587], Fresh[28586], Fresh[28585], Fresh[28584], Fresh[28583], Fresh[28582], Fresh[28581], Fresh[28580], Fresh[28579], Fresh[28578], Fresh[28577], Fresh[28576], Fresh[28575], Fresh[28574], Fresh[28573], Fresh[28572], Fresh[28571], Fresh[28570], Fresh[28569], Fresh[28568], Fresh[28567], Fresh[28566], Fresh[28565], Fresh[28564], Fresh[28563], Fresh[28562], Fresh[28561], Fresh[28560], Fresh[28559], Fresh[28558], Fresh[28557], Fresh[28556], Fresh[28555], Fresh[28554], Fresh[28553], Fresh[28552], Fresh[28551], Fresh[28550], Fresh[28549], Fresh[28548], Fresh[28547], Fresh[28546], Fresh[28545], Fresh[28544], Fresh[28543], Fresh[28542], Fresh[28541], Fresh[28540], Fresh[28539], Fresh[28538], Fresh[28537], Fresh[28536], Fresh[28535], Fresh[28534], Fresh[28533], Fresh[28532], Fresh[28531], Fresh[28530], Fresh[28529], Fresh[28528], Fresh[28527], Fresh[28526], Fresh[28525], Fresh[28524], Fresh[28523], Fresh[28522], Fresh[28521], Fresh[28520], Fresh[28519], Fresh[28518], Fresh[28517], Fresh[28516], Fresh[28515], Fresh[28514], Fresh[28513], Fresh[28512], Fresh[28511], Fresh[28510], Fresh[28509], Fresh[28508], Fresh[28507], Fresh[28506], Fresh[28505], Fresh[28504], Fresh[28503], Fresh[28502], Fresh[28501], Fresh[28500], Fresh[28499], Fresh[28498], Fresh[28497], Fresh[28496], Fresh[28495], Fresh[28494], Fresh[28493], Fresh[28492], Fresh[28491], Fresh[28490], Fresh[28489], Fresh[28488], Fresh[28487], Fresh[28486], Fresh[28485], Fresh[28484], Fresh[28483], Fresh[28482], Fresh[28481], Fresh[28480], Fresh[28479], Fresh[28478], Fresh[28477], Fresh[28476], Fresh[28475], Fresh[28474], Fresh[28473], Fresh[28472], Fresh[28471], Fresh[28470], Fresh[28469], Fresh[28468], Fresh[28467], Fresh[28466], Fresh[28465], Fresh[28464], Fresh[28463], Fresh[28462], Fresh[28461], Fresh[28460], Fresh[28459], Fresh[28458], Fresh[28457], Fresh[28456], Fresh[28455], Fresh[28454], Fresh[28453], Fresh[28452], Fresh[28451], Fresh[28450], Fresh[28449], Fresh[28448], Fresh[28447], Fresh[28446], Fresh[28445], Fresh[28444], Fresh[28443], Fresh[28442], Fresh[28441], Fresh[28440], Fresh[28439], Fresh[28438], Fresh[28437], Fresh[28436], Fresh[28435], Fresh[28434], Fresh[28433], Fresh[28432], Fresh[28431], Fresh[28430], Fresh[28429], Fresh[28428], Fresh[28427], Fresh[28426], Fresh[28425], Fresh[28424], Fresh[28423], Fresh[28422], Fresh[28421], Fresh[28420], Fresh[28419], Fresh[28418], Fresh[28417], Fresh[28416], Fresh[28415], Fresh[28414], Fresh[28413], Fresh[28412], Fresh[28411], Fresh[28410], Fresh[28409], Fresh[28408], Fresh[28407], Fresh[28406], Fresh[28405], Fresh[28404], Fresh[28403], Fresh[28402], Fresh[28401], Fresh[28400], Fresh[28399], Fresh[28398], Fresh[28397], Fresh[28396], Fresh[28395], Fresh[28394], Fresh[28393], Fresh[28392], Fresh[28391], Fresh[28390], Fresh[28389], Fresh[28388], Fresh[28387], Fresh[28386], Fresh[28385], Fresh[28384], Fresh[28383], Fresh[28382], Fresh[28381], Fresh[28380], Fresh[28379], Fresh[28378], Fresh[28377], Fresh[28376], Fresh[28375], Fresh[28374], Fresh[28373], Fresh[28372], Fresh[28371], Fresh[28370], Fresh[28369], Fresh[28368], Fresh[28367], Fresh[28366], Fresh[28365], Fresh[28364], Fresh[28363], Fresh[28362], Fresh[28361], Fresh[28360], Fresh[28359], Fresh[28358], Fresh[28357], Fresh[28356], Fresh[28355], Fresh[28354], Fresh[28353], Fresh[28352], Fresh[28351], Fresh[28350], Fresh[28349], Fresh[28348], Fresh[28347], Fresh[28346], Fresh[28345], Fresh[28344], Fresh[28343], Fresh[28342], Fresh[28341], Fresh[28340], Fresh[28339], Fresh[28338], Fresh[28337], Fresh[28336], Fresh[28335], Fresh[28334], Fresh[28333], Fresh[28332], Fresh[28331], Fresh[28330], Fresh[28329], Fresh[28328], Fresh[28327], Fresh[28326], Fresh[28325], Fresh[28324], Fresh[28323], Fresh[28322], Fresh[28321], Fresh[28320], Fresh[28319], Fresh[28318], Fresh[28317], Fresh[28316], Fresh[28315], Fresh[28314], Fresh[28313], Fresh[28312], Fresh[28311], Fresh[28310], Fresh[28309], Fresh[28308], Fresh[28307], Fresh[28306], Fresh[28305], Fresh[28304], Fresh[28303], Fresh[28302], Fresh[28301], Fresh[28300], Fresh[28299], Fresh[28298], Fresh[28297], Fresh[28296], Fresh[28295], Fresh[28294], Fresh[28293], Fresh[28292], Fresh[28291], Fresh[28290], Fresh[28289], Fresh[28288], Fresh[28287], Fresh[28286], Fresh[28285], Fresh[28284], Fresh[28283], Fresh[28282], Fresh[28281], Fresh[28280], Fresh[28279], Fresh[28278], Fresh[28277], Fresh[28276], Fresh[28275], Fresh[28274], Fresh[28273], Fresh[28272], Fresh[28271], Fresh[28270], Fresh[28269], Fresh[28268], Fresh[28267], Fresh[28266], Fresh[28265], Fresh[28264], Fresh[28263], Fresh[28262], Fresh[28261], Fresh[28260], Fresh[28259], Fresh[28258], Fresh[28257], Fresh[28256], Fresh[28255], Fresh[28254], Fresh[28253], Fresh[28252], Fresh[28251], Fresh[28250], Fresh[28249], Fresh[28248], Fresh[28247], Fresh[28246], Fresh[28245], Fresh[28244], Fresh[28243], Fresh[28242], Fresh[28241], Fresh[28240], Fresh[28239], Fresh[28238], Fresh[28237], Fresh[28236], Fresh[28235], Fresh[28234], Fresh[28233], Fresh[28232], Fresh[28231], Fresh[28230], Fresh[28229], Fresh[28228], Fresh[28227], Fresh[28226], Fresh[28225], Fresh[28224], Fresh[28223], Fresh[28222], Fresh[28221], Fresh[28220], Fresh[28219], Fresh[28218], Fresh[28217], Fresh[28216], Fresh[28215], Fresh[28214], Fresh[28213], Fresh[28212], Fresh[28211], Fresh[28210], Fresh[28209], Fresh[28208], Fresh[28207], Fresh[28206], Fresh[28205], Fresh[28204], Fresh[28203], Fresh[28202], Fresh[28201], Fresh[28200], Fresh[28199], Fresh[28198], Fresh[28197], Fresh[28196], Fresh[28195], Fresh[28194], Fresh[28193], Fresh[28192], Fresh[28191], Fresh[28190], Fresh[28189], Fresh[28188], Fresh[28187], Fresh[28186], Fresh[28185], Fresh[28184], Fresh[28183], Fresh[28182], Fresh[28181], Fresh[28180], Fresh[28179], Fresh[28178], Fresh[28177], Fresh[28176], Fresh[28175], Fresh[28174], Fresh[28173], Fresh[28172], Fresh[28171], Fresh[28170], Fresh[28169], Fresh[28168], Fresh[28167], Fresh[28166], Fresh[28165], Fresh[28164], Fresh[28163], Fresh[28162], Fresh[28161], Fresh[28160], Fresh[28159], Fresh[28158], Fresh[28157], Fresh[28156], Fresh[28155], Fresh[28154], Fresh[28153], Fresh[28152], Fresh[28151], Fresh[28150], Fresh[28149], Fresh[28148], Fresh[28147], Fresh[28146], Fresh[28145], Fresh[28144], Fresh[28143], Fresh[28142], Fresh[28141], Fresh[28140], Fresh[28139], Fresh[28138], Fresh[28137], Fresh[28136], Fresh[28135], Fresh[28134], Fresh[28133], Fresh[28132], Fresh[28131], Fresh[28130], Fresh[28129], Fresh[28128], Fresh[28127], Fresh[28126], Fresh[28125], Fresh[28124], Fresh[28123], Fresh[28122], Fresh[28121], Fresh[28120], Fresh[28119], Fresh[28118], Fresh[28117], Fresh[28116], Fresh[28115], Fresh[28114], Fresh[28113], Fresh[28112], Fresh[28111], Fresh[28110], Fresh[28109], Fresh[28108], Fresh[28107], Fresh[28106], Fresh[28105], Fresh[28104], Fresh[28103], Fresh[28102], Fresh[28101], Fresh[28100], Fresh[28099], Fresh[28098], Fresh[28097], Fresh[28096], Fresh[28095], Fresh[28094], Fresh[28093], Fresh[28092], Fresh[28091], Fresh[28090], Fresh[28089], Fresh[28088], Fresh[28087], Fresh[28086], Fresh[28085], Fresh[28084], Fresh[28083], Fresh[28082], Fresh[28081], Fresh[28080], Fresh[28079], Fresh[28078], Fresh[28077], Fresh[28076], Fresh[28075], Fresh[28074], Fresh[28073], Fresh[28072], Fresh[28071], Fresh[28070], Fresh[28069], Fresh[28068], Fresh[28067], Fresh[28066], Fresh[28065], Fresh[28064], Fresh[28063], Fresh[28062], Fresh[28061], Fresh[28060], Fresh[28059], Fresh[28058], Fresh[28057], Fresh[28056], Fresh[28055], Fresh[28054], Fresh[28053], Fresh[28052], Fresh[28051], Fresh[28050], Fresh[28049], Fresh[28048], Fresh[28047], Fresh[28046], Fresh[28045], Fresh[28044], Fresh[28043], Fresh[28042], Fresh[28041], Fresh[28040], Fresh[28039], Fresh[28038], Fresh[28037], Fresh[28036], Fresh[28035], Fresh[28034], Fresh[28033], Fresh[28032], Fresh[28031], Fresh[28030], Fresh[28029], Fresh[28028], Fresh[28027], Fresh[28026], Fresh[28025], Fresh[28024], Fresh[28023], Fresh[28022], Fresh[28021], Fresh[28020], Fresh[28019], Fresh[28018], Fresh[28017], Fresh[28016], Fresh[28015], Fresh[28014], Fresh[28013], Fresh[28012], Fresh[28011], Fresh[28010], Fresh[28009], Fresh[28008], Fresh[28007], Fresh[28006], Fresh[28005], Fresh[28004], Fresh[28003], Fresh[28002], Fresh[28001], Fresh[28000], Fresh[27999], Fresh[27998], Fresh[27997], Fresh[27996], Fresh[27995], Fresh[27994], Fresh[27993], Fresh[27992], Fresh[27991], Fresh[27990], Fresh[27989], Fresh[27988], Fresh[27987], Fresh[27986], Fresh[27985], Fresh[27984], Fresh[27983], Fresh[27982], Fresh[27981], Fresh[27980], Fresh[27979], Fresh[27978], Fresh[27977], Fresh[27976], Fresh[27975], Fresh[27974], Fresh[27973], Fresh[27972], Fresh[27971], Fresh[27970], Fresh[27969], Fresh[27968], Fresh[27967], Fresh[27966], Fresh[27965], Fresh[27964], Fresh[27963], Fresh[27962], Fresh[27961], Fresh[27960], Fresh[27959], Fresh[27958], Fresh[27957], Fresh[27956], Fresh[27955], Fresh[27954], Fresh[27953], Fresh[27952], Fresh[27951], Fresh[27950], Fresh[27949], Fresh[27948], Fresh[27947], Fresh[27946], Fresh[27945], Fresh[27944], Fresh[27943], Fresh[27942], Fresh[27941], Fresh[27940], Fresh[27939], Fresh[27938], Fresh[27937], Fresh[27936], Fresh[27935], Fresh[27934], Fresh[27933], Fresh[27932], Fresh[27931], Fresh[27930], Fresh[27929], Fresh[27928], Fresh[27927], Fresh[27926], Fresh[27925], Fresh[27924], Fresh[27923], Fresh[27922], Fresh[27921], Fresh[27920], Fresh[27919], Fresh[27918], Fresh[27917], Fresh[27916], Fresh[27915], Fresh[27914], Fresh[27913], Fresh[27912], Fresh[27911], Fresh[27910], Fresh[27909], Fresh[27908], Fresh[27907], Fresh[27906], Fresh[27905], Fresh[27904], Fresh[27903], Fresh[27902], Fresh[27901], Fresh[27900], Fresh[27899], Fresh[27898], Fresh[27897], Fresh[27896], Fresh[27895], Fresh[27894], Fresh[27893], Fresh[27892], Fresh[27891], Fresh[27890], Fresh[27889], Fresh[27888], Fresh[27887], Fresh[27886], Fresh[27885], Fresh[27884], Fresh[27883], Fresh[27882], Fresh[27881], Fresh[27880], Fresh[27879], Fresh[27878], Fresh[27877], Fresh[27876], Fresh[27875], Fresh[27874], Fresh[27873], Fresh[27872], Fresh[27871], Fresh[27870], Fresh[27869], Fresh[27868], Fresh[27867], Fresh[27866], Fresh[27865], Fresh[27864], Fresh[27863], Fresh[27862], Fresh[27861], Fresh[27860], Fresh[27859], Fresh[27858], Fresh[27857], Fresh[27856], Fresh[27855], Fresh[27854], Fresh[27853], Fresh[27852], Fresh[27851], Fresh[27850], Fresh[27849], Fresh[27848], Fresh[27847], Fresh[27846], Fresh[27845], Fresh[27844], Fresh[27843], Fresh[27842], Fresh[27841], Fresh[27840], Fresh[27839], Fresh[27838], Fresh[27837], Fresh[27836], Fresh[27835], Fresh[27834], Fresh[27833], Fresh[27832], Fresh[27831], Fresh[27830], Fresh[27829], Fresh[27828], Fresh[27827], Fresh[27826], Fresh[27825], Fresh[27824], Fresh[27823], Fresh[27822], Fresh[27821], Fresh[27820], Fresh[27819], Fresh[27818], Fresh[27817], Fresh[27816], Fresh[27815], Fresh[27814], Fresh[27813], Fresh[27812], Fresh[27811], Fresh[27810], Fresh[27809], Fresh[27808], Fresh[27807], Fresh[27806], Fresh[27805], Fresh[27804], Fresh[27803], Fresh[27802], Fresh[27801], Fresh[27800], Fresh[27799], Fresh[27798], Fresh[27797], Fresh[27796], Fresh[27795], Fresh[27794], Fresh[27793], Fresh[27792], Fresh[27791], Fresh[27790], Fresh[27789], Fresh[27788], Fresh[27787], Fresh[27786], Fresh[27785], Fresh[27784], Fresh[27783], Fresh[27782], Fresh[27781], Fresh[27780], Fresh[27779], Fresh[27778], Fresh[27777], Fresh[27776], Fresh[27775], Fresh[27774], Fresh[27773], Fresh[27772], Fresh[27771], Fresh[27770], Fresh[27769], Fresh[27768], Fresh[27767], Fresh[27766], Fresh[27765], Fresh[27764], Fresh[27763], Fresh[27762], Fresh[27761], Fresh[27760], Fresh[27759], Fresh[27758], Fresh[27757], Fresh[27756], Fresh[27755], Fresh[27754], Fresh[27753], Fresh[27752], Fresh[27751], Fresh[27750], Fresh[27749], Fresh[27748], Fresh[27747], Fresh[27746], Fresh[27745], Fresh[27744], Fresh[27743], Fresh[27742], Fresh[27741], Fresh[27740], Fresh[27739], Fresh[27738], Fresh[27737], Fresh[27736], Fresh[27735], Fresh[27734], Fresh[27733], Fresh[27732], Fresh[27731], Fresh[27730], Fresh[27729], Fresh[27728], Fresh[27727], Fresh[27726], Fresh[27725], Fresh[27724], Fresh[27723], Fresh[27722], Fresh[27721], Fresh[27720], Fresh[27719], Fresh[27718], Fresh[27717], Fresh[27716], Fresh[27715], Fresh[27714], Fresh[27713], Fresh[27712], Fresh[27711], Fresh[27710], Fresh[27709], Fresh[27708], Fresh[27707], Fresh[27706], Fresh[27705], Fresh[27704], Fresh[27703], Fresh[27702], Fresh[27701], Fresh[27700], Fresh[27699], Fresh[27698], Fresh[27697], Fresh[27696], Fresh[27695], Fresh[27694], Fresh[27693], Fresh[27692], Fresh[27691], Fresh[27690], Fresh[27689], Fresh[27688], Fresh[27687], Fresh[27686], Fresh[27685], Fresh[27684], Fresh[27683], Fresh[27682], Fresh[27681], Fresh[27680], Fresh[27679], Fresh[27678], Fresh[27677], Fresh[27676], Fresh[27675], Fresh[27674], Fresh[27673], Fresh[27672], Fresh[27671], Fresh[27670], Fresh[27669], Fresh[27668], Fresh[27667], Fresh[27666], Fresh[27665], Fresh[27664], Fresh[27663], Fresh[27662], Fresh[27661], Fresh[27660], Fresh[27659], Fresh[27658], Fresh[27657], Fresh[27656], Fresh[27655], Fresh[27654], Fresh[27653], Fresh[27652], Fresh[27651], Fresh[27650], Fresh[27649], Fresh[27648], Fresh[27647], Fresh[27646], Fresh[27645], Fresh[27644], Fresh[27643], Fresh[27642], Fresh[27641], Fresh[27640], Fresh[27639], Fresh[27638], Fresh[27637], Fresh[27636], Fresh[27635], Fresh[27634], Fresh[27633], Fresh[27632], Fresh[27631], Fresh[27630], Fresh[27629], Fresh[27628], Fresh[27627], Fresh[27626], Fresh[27625], Fresh[27624], Fresh[27623], Fresh[27622], Fresh[27621], Fresh[27620], Fresh[27619], Fresh[27618], Fresh[27617], Fresh[27616], Fresh[27615], Fresh[27614], Fresh[27613], Fresh[27612], Fresh[27611], Fresh[27610], Fresh[27609], Fresh[27608], Fresh[27607], Fresh[27606], Fresh[27605], Fresh[27604], Fresh[27603], Fresh[27602], Fresh[27601], Fresh[27600], Fresh[27599], Fresh[27598], Fresh[27597], Fresh[27596], Fresh[27595], Fresh[27594], Fresh[27593], Fresh[27592], Fresh[27591], Fresh[27590], Fresh[27589], Fresh[27588], Fresh[27587], Fresh[27586], Fresh[27585], Fresh[27584], Fresh[27583], Fresh[27582], Fresh[27581], Fresh[27580], Fresh[27579], Fresh[27578], Fresh[27577], Fresh[27576], Fresh[27575], Fresh[27574], Fresh[27573], Fresh[27572], Fresh[27571], Fresh[27570], Fresh[27569], Fresh[27568], Fresh[27567], Fresh[27566], Fresh[27565], Fresh[27564], Fresh[27563], Fresh[27562], Fresh[27561], Fresh[27560], Fresh[27559], Fresh[27558], Fresh[27557], Fresh[27556], Fresh[27555], Fresh[27554], Fresh[27553], Fresh[27552], Fresh[27551], Fresh[27550], Fresh[27549], Fresh[27548], Fresh[27547], Fresh[27546], Fresh[27545], Fresh[27544], Fresh[27543], Fresh[27542], Fresh[27541], Fresh[27540], Fresh[27539], Fresh[27538], Fresh[27537], Fresh[27536], Fresh[27535], Fresh[27534], Fresh[27533], Fresh[27532], Fresh[27531], Fresh[27530], Fresh[27529], Fresh[27528], Fresh[27527], Fresh[27526], Fresh[27525], Fresh[27524], Fresh[27523], Fresh[27522], Fresh[27521], Fresh[27520], Fresh[27519], Fresh[27518], Fresh[27517], Fresh[27516], Fresh[27515], Fresh[27514], Fresh[27513], Fresh[27512], Fresh[27511], Fresh[27510], Fresh[27509], Fresh[27508], Fresh[27507], Fresh[27506], Fresh[27505], Fresh[27504], Fresh[27503], Fresh[27502], Fresh[27501], Fresh[27500], Fresh[27499], Fresh[27498], Fresh[27497], Fresh[27496], Fresh[27495], Fresh[27494], Fresh[27493], Fresh[27492], Fresh[27491], Fresh[27490], Fresh[27489], Fresh[27488], Fresh[27487], Fresh[27486], Fresh[27485], Fresh[27484], Fresh[27483], Fresh[27482], Fresh[27481], Fresh[27480], Fresh[27479], Fresh[27478], Fresh[27477], Fresh[27476], Fresh[27475], Fresh[27474], Fresh[27473], Fresh[27472], Fresh[27471], Fresh[27470], Fresh[27469], Fresh[27468], Fresh[27467], Fresh[27466], Fresh[27465], Fresh[27464], Fresh[27463], Fresh[27462], Fresh[27461], Fresh[27460], Fresh[27459], Fresh[27458], Fresh[27457], Fresh[27456], Fresh[27455], Fresh[27454], Fresh[27453], Fresh[27452], Fresh[27451], Fresh[27450], Fresh[27449], Fresh[27448], Fresh[27447], Fresh[27446], Fresh[27445], Fresh[27444], Fresh[27443], Fresh[27442], Fresh[27441], Fresh[27440], Fresh[27439], Fresh[27438], Fresh[27437], Fresh[27436], Fresh[27435], Fresh[27434], Fresh[27433], Fresh[27432], Fresh[27431], Fresh[27430], Fresh[27429], Fresh[27428], Fresh[27427], Fresh[27426], Fresh[27425], Fresh[27424], Fresh[27423], Fresh[27422], Fresh[27421], Fresh[27420], Fresh[27419], Fresh[27418], Fresh[27417], Fresh[27416], Fresh[27415], Fresh[27414], Fresh[27413], Fresh[27412], Fresh[27411], Fresh[27410], Fresh[27409], Fresh[27408], Fresh[27407], Fresh[27406], Fresh[27405], Fresh[27404], Fresh[27403], Fresh[27402], Fresh[27401], Fresh[27400], Fresh[27399], Fresh[27398], Fresh[27397], Fresh[27396], Fresh[27395], Fresh[27394], Fresh[27393], Fresh[27392], Fresh[27391], Fresh[27390], Fresh[27389], Fresh[27388], Fresh[27387], Fresh[27386], Fresh[27385], Fresh[27384], Fresh[27383], Fresh[27382], Fresh[27381], Fresh[27380], Fresh[27379], Fresh[27378], Fresh[27377], Fresh[27376], Fresh[27375], Fresh[27374], Fresh[27373], Fresh[27372], Fresh[27371], Fresh[27370], Fresh[27369], Fresh[27368], Fresh[27367], Fresh[27366], Fresh[27365], Fresh[27364], Fresh[27363], Fresh[27362], Fresh[27361], Fresh[27360], Fresh[27359], Fresh[27358], Fresh[27357], Fresh[27356], Fresh[27355], Fresh[27354], Fresh[27353], Fresh[27352], Fresh[27351], Fresh[27350], Fresh[27349], Fresh[27348], Fresh[27347], Fresh[27346], Fresh[27345], Fresh[27344], Fresh[27343], Fresh[27342], Fresh[27341], Fresh[27340], Fresh[27339], Fresh[27338], Fresh[27337], Fresh[27336], Fresh[27335], Fresh[27334], Fresh[27333], Fresh[27332], Fresh[27331], Fresh[27330], Fresh[27329], Fresh[27328], Fresh[27327], Fresh[27326], Fresh[27325], Fresh[27324], Fresh[27323], Fresh[27322], Fresh[27321], Fresh[27320], Fresh[27319], Fresh[27318], Fresh[27317], Fresh[27316], Fresh[27315], Fresh[27314], Fresh[27313], Fresh[27312], Fresh[27311], Fresh[27310], Fresh[27309], Fresh[27308], Fresh[27307], Fresh[27306], Fresh[27305], Fresh[27304], Fresh[27303], Fresh[27302], Fresh[27301], Fresh[27300], Fresh[27299], Fresh[27298], Fresh[27297], Fresh[27296], Fresh[27295], Fresh[27294], Fresh[27293], Fresh[27292], Fresh[27291], Fresh[27290], Fresh[27289], Fresh[27288], Fresh[27287], Fresh[27286], Fresh[27285], Fresh[27284], Fresh[27283], Fresh[27282], Fresh[27281], Fresh[27280], Fresh[27279], Fresh[27278], Fresh[27277], Fresh[27276], Fresh[27275], Fresh[27274], Fresh[27273], Fresh[27272], Fresh[27271], Fresh[27270], Fresh[27269], Fresh[27268], Fresh[27267], Fresh[27266], Fresh[27265], Fresh[27264], Fresh[27263], Fresh[27262], Fresh[27261], Fresh[27260], Fresh[27259], Fresh[27258], Fresh[27257], Fresh[27256], Fresh[27255], Fresh[27254], Fresh[27253], Fresh[27252], Fresh[27251], Fresh[27250], Fresh[27249], Fresh[27248], Fresh[27247], Fresh[27246], Fresh[27245], Fresh[27244], Fresh[27243], Fresh[27242], Fresh[27241], Fresh[27240], Fresh[27239], Fresh[27238], Fresh[27237], Fresh[27236], Fresh[27235], Fresh[27234], Fresh[27233], Fresh[27232], Fresh[27231], Fresh[27230], Fresh[27229], Fresh[27228], Fresh[27227], Fresh[27226], Fresh[27225], Fresh[27224], Fresh[27223], Fresh[27222], Fresh[27221], Fresh[27220], Fresh[27219], Fresh[27218], Fresh[27217], Fresh[27216], Fresh[27215], Fresh[27214], Fresh[27213], Fresh[27212], Fresh[27211], Fresh[27210], Fresh[27209], Fresh[27208], Fresh[27207], Fresh[27206], Fresh[27205], Fresh[27204], Fresh[27203], Fresh[27202], Fresh[27201], Fresh[27200], Fresh[27199], Fresh[27198], Fresh[27197], Fresh[27196], Fresh[27195], Fresh[27194], Fresh[27193], Fresh[27192], Fresh[27191], Fresh[27190], Fresh[27189], Fresh[27188], Fresh[27187], Fresh[27186], Fresh[27185], Fresh[27184], Fresh[27183], Fresh[27182], Fresh[27181], Fresh[27180], Fresh[27179], Fresh[27178], Fresh[27177], Fresh[27176], Fresh[27175], Fresh[27174], Fresh[27173], Fresh[27172], Fresh[27171], Fresh[27170], Fresh[27169], Fresh[27168], Fresh[27167], Fresh[27166], Fresh[27165], Fresh[27164], Fresh[27163], Fresh[27162], Fresh[27161], Fresh[27160], Fresh[27159], Fresh[27158], Fresh[27157], Fresh[27156], Fresh[27155], Fresh[27154], Fresh[27153], Fresh[27152], Fresh[27151], Fresh[27150], Fresh[27149], Fresh[27148], Fresh[27147], Fresh[27146], Fresh[27145], Fresh[27144], Fresh[27143], Fresh[27142], Fresh[27141], Fresh[27140], Fresh[27139], Fresh[27138], Fresh[27137], Fresh[27136], Fresh[27135], Fresh[27134], Fresh[27133], Fresh[27132], Fresh[27131], Fresh[27130], Fresh[27129], Fresh[27128], Fresh[27127], Fresh[27126], Fresh[27125], Fresh[27124], Fresh[27123], Fresh[27122], Fresh[27121], Fresh[27120], Fresh[27119], Fresh[27118], Fresh[27117], Fresh[27116], Fresh[27115], Fresh[27114], Fresh[27113], Fresh[27112], Fresh[27111], Fresh[27110], Fresh[27109], Fresh[27108], Fresh[27107], Fresh[27106], Fresh[27105], Fresh[27104], Fresh[27103], Fresh[27102], Fresh[27101], Fresh[27100], Fresh[27099], Fresh[27098], Fresh[27097], Fresh[27096], Fresh[27095], Fresh[27094], Fresh[27093], Fresh[27092], Fresh[27091], Fresh[27090], Fresh[27089], Fresh[27088], Fresh[27087], Fresh[27086], Fresh[27085], Fresh[27084], Fresh[27083], Fresh[27082], Fresh[27081], Fresh[27080], Fresh[27079], Fresh[27078], Fresh[27077], Fresh[27076], Fresh[27075], Fresh[27074], Fresh[27073], Fresh[27072], Fresh[27071], Fresh[27070], Fresh[27069], Fresh[27068], Fresh[27067], Fresh[27066], Fresh[27065], Fresh[27064], Fresh[27063], Fresh[27062], Fresh[27061], Fresh[27060], Fresh[27059], Fresh[27058], Fresh[27057], Fresh[27056], Fresh[27055], Fresh[27054], Fresh[27053], Fresh[27052], Fresh[27051], Fresh[27050], Fresh[27049], Fresh[27048], Fresh[27047], Fresh[27046], Fresh[27045], Fresh[27044], Fresh[27043], Fresh[27042], Fresh[27041], Fresh[27040], Fresh[27039], Fresh[27038], Fresh[27037], Fresh[27036], Fresh[27035], Fresh[27034], Fresh[27033], Fresh[27032], Fresh[27031], Fresh[27030], Fresh[27029], Fresh[27028], Fresh[27027], Fresh[27026], Fresh[27025], Fresh[27024], Fresh[27023], Fresh[27022], Fresh[27021], Fresh[27020], Fresh[27019], Fresh[27018], Fresh[27017], Fresh[27016], Fresh[27015], Fresh[27014], Fresh[27013], Fresh[27012], Fresh[27011], Fresh[27010], Fresh[27009], Fresh[27008], Fresh[27007], Fresh[27006], Fresh[27005], Fresh[27004], Fresh[27003], Fresh[27002], Fresh[27001], Fresh[27000], Fresh[26999], Fresh[26998], Fresh[26997], Fresh[26996], Fresh[26995], Fresh[26994], Fresh[26993], Fresh[26992], Fresh[26991], Fresh[26990], Fresh[26989], Fresh[26988], Fresh[26987], Fresh[26986], Fresh[26985], Fresh[26984], Fresh[26983], Fresh[26982], Fresh[26981], Fresh[26980], Fresh[26979], Fresh[26978], Fresh[26977], Fresh[26976], Fresh[26975], Fresh[26974], Fresh[26973], Fresh[26972], Fresh[26971], Fresh[26970], Fresh[26969], Fresh[26968], Fresh[26967], Fresh[26966], Fresh[26965], Fresh[26964], Fresh[26963], Fresh[26962], Fresh[26961], Fresh[26960], Fresh[26959], Fresh[26958], Fresh[26957], Fresh[26956], Fresh[26955], Fresh[26954], Fresh[26953], Fresh[26952], Fresh[26951], Fresh[26950], Fresh[26949], Fresh[26948], Fresh[26947], Fresh[26946], Fresh[26945], Fresh[26944], Fresh[26943], Fresh[26942], Fresh[26941], Fresh[26940], Fresh[26939], Fresh[26938], Fresh[26937], Fresh[26936], Fresh[26935], Fresh[26934], Fresh[26933], Fresh[26932], Fresh[26931], Fresh[26930], Fresh[26929], Fresh[26928], Fresh[26927], Fresh[26926], Fresh[26925], Fresh[26924], Fresh[26923], Fresh[26922], Fresh[26921], Fresh[26920], Fresh[26919], Fresh[26918], Fresh[26917], Fresh[26916], Fresh[26915], Fresh[26914], Fresh[26913], Fresh[26912], Fresh[26911], Fresh[26910], Fresh[26909], Fresh[26908], Fresh[26907], Fresh[26906], Fresh[26905], Fresh[26904], Fresh[26903], Fresh[26902], Fresh[26901], Fresh[26900], Fresh[26899], Fresh[26898], Fresh[26897], Fresh[26896], Fresh[26895], Fresh[26894], Fresh[26893], Fresh[26892], Fresh[26891], Fresh[26890], Fresh[26889], Fresh[26888], Fresh[26887], Fresh[26886], Fresh[26885], Fresh[26884], Fresh[26883], Fresh[26882], Fresh[26881], Fresh[26880], Fresh[26879], Fresh[26878], Fresh[26877], Fresh[26876], Fresh[26875], Fresh[26874], Fresh[26873], Fresh[26872], Fresh[26871], Fresh[26870], Fresh[26869], Fresh[26868], Fresh[26867], Fresh[26866], Fresh[26865], Fresh[26864], Fresh[26863], Fresh[26862], Fresh[26861], Fresh[26860], Fresh[26859], Fresh[26858], Fresh[26857], Fresh[26856], Fresh[26855], Fresh[26854], Fresh[26853], Fresh[26852], Fresh[26851], Fresh[26850], Fresh[26849], Fresh[26848], Fresh[26847], Fresh[26846], Fresh[26845], Fresh[26844], Fresh[26843], Fresh[26842], Fresh[26841], Fresh[26840], Fresh[26839], Fresh[26838], Fresh[26837], Fresh[26836], Fresh[26835], Fresh[26834], Fresh[26833], Fresh[26832], Fresh[26831], Fresh[26830], Fresh[26829], Fresh[26828], Fresh[26827], Fresh[26826], Fresh[26825], Fresh[26824], Fresh[26823], Fresh[26822], Fresh[26821], Fresh[26820], Fresh[26819], Fresh[26818], Fresh[26817], Fresh[26816], Fresh[26815], Fresh[26814], Fresh[26813], Fresh[26812], Fresh[26811], Fresh[26810], Fresh[26809], Fresh[26808], Fresh[26807], Fresh[26806], Fresh[26805], Fresh[26804], Fresh[26803], Fresh[26802], Fresh[26801], Fresh[26800], Fresh[26799], Fresh[26798], Fresh[26797], Fresh[26796], Fresh[26795], Fresh[26794], Fresh[26793], Fresh[26792], Fresh[26791], Fresh[26790], Fresh[26789], Fresh[26788], Fresh[26787], Fresh[26786], Fresh[26785], Fresh[26784], Fresh[26783], Fresh[26782], Fresh[26781], Fresh[26780], Fresh[26779], Fresh[26778], Fresh[26777], Fresh[26776], Fresh[26775], Fresh[26774], Fresh[26773], Fresh[26772], Fresh[26771], Fresh[26770], Fresh[26769], Fresh[26768], Fresh[26767], Fresh[26766], Fresh[26765], Fresh[26764], Fresh[26763], Fresh[26762], Fresh[26761], Fresh[26760], Fresh[26759], Fresh[26758], Fresh[26757], Fresh[26756], Fresh[26755], Fresh[26754], Fresh[26753], Fresh[26752], Fresh[26751], Fresh[26750], Fresh[26749], Fresh[26748], Fresh[26747], Fresh[26746], Fresh[26745], Fresh[26744], Fresh[26743], Fresh[26742], Fresh[26741], Fresh[26740], Fresh[26739], Fresh[26738], Fresh[26737], Fresh[26736], Fresh[26735], Fresh[26734], Fresh[26733], Fresh[26732], Fresh[26731], Fresh[26730], Fresh[26729], Fresh[26728], Fresh[26727], Fresh[26726], Fresh[26725], Fresh[26724], Fresh[26723], Fresh[26722], Fresh[26721], Fresh[26720], Fresh[26719], Fresh[26718], Fresh[26717], Fresh[26716], Fresh[26715], Fresh[26714], Fresh[26713], Fresh[26712], Fresh[26711], Fresh[26710], Fresh[26709], Fresh[26708], Fresh[26707], Fresh[26706], Fresh[26705], Fresh[26704], Fresh[26703], Fresh[26702], Fresh[26701], Fresh[26700], Fresh[26699], Fresh[26698], Fresh[26697], Fresh[26696], Fresh[26695], Fresh[26694], Fresh[26693], Fresh[26692], Fresh[26691], Fresh[26690], Fresh[26689], Fresh[26688], Fresh[26687], Fresh[26686], Fresh[26685], Fresh[26684], Fresh[26683], Fresh[26682], Fresh[26681], Fresh[26680], Fresh[26679], Fresh[26678], Fresh[26677], Fresh[26676], Fresh[26675], Fresh[26674], Fresh[26673], Fresh[26672], Fresh[26671], Fresh[26670], Fresh[26669], Fresh[26668], Fresh[26667], Fresh[26666], Fresh[26665], Fresh[26664], Fresh[26663], Fresh[26662], Fresh[26661], Fresh[26660], Fresh[26659], Fresh[26658], Fresh[26657], Fresh[26656], Fresh[26655], Fresh[26654], Fresh[26653], Fresh[26652], Fresh[26651], Fresh[26650], Fresh[26649], Fresh[26648], Fresh[26647], Fresh[26646], Fresh[26645], Fresh[26644], Fresh[26643], Fresh[26642], Fresh[26641], Fresh[26640], Fresh[26639], Fresh[26638], Fresh[26637], Fresh[26636], Fresh[26635], Fresh[26634], Fresh[26633], Fresh[26632], Fresh[26631], Fresh[26630], Fresh[26629], Fresh[26628], Fresh[26627], Fresh[26626], Fresh[26625], Fresh[26624], Fresh[26623], Fresh[26622], Fresh[26621], Fresh[26620], Fresh[26619], Fresh[26618], Fresh[26617], Fresh[26616], Fresh[26615], Fresh[26614], Fresh[26613], Fresh[26612], Fresh[26611], Fresh[26610], Fresh[26609], Fresh[26608], Fresh[26607], Fresh[26606], Fresh[26605], Fresh[26604], Fresh[26603], Fresh[26602], Fresh[26601], Fresh[26600], Fresh[26599], Fresh[26598], Fresh[26597], Fresh[26596], Fresh[26595], Fresh[26594], Fresh[26593], Fresh[26592], Fresh[26591], Fresh[26590], Fresh[26589], Fresh[26588], Fresh[26587], Fresh[26586], Fresh[26585], Fresh[26584], Fresh[26583], Fresh[26582], Fresh[26581], Fresh[26580], Fresh[26579], Fresh[26578], Fresh[26577], Fresh[26576], Fresh[26575], Fresh[26574], Fresh[26573], Fresh[26572], Fresh[26571], Fresh[26570], Fresh[26569], Fresh[26568], Fresh[26567], Fresh[26566], Fresh[26565], Fresh[26564], Fresh[26563], Fresh[26562], Fresh[26561], Fresh[26560], Fresh[26559], Fresh[26558], Fresh[26557], Fresh[26556], Fresh[26555], Fresh[26554], Fresh[26553], Fresh[26552], Fresh[26551], Fresh[26550], Fresh[26549], Fresh[26548], Fresh[26547], Fresh[26546], Fresh[26545], Fresh[26544], Fresh[26543], Fresh[26542], Fresh[26541], Fresh[26540], Fresh[26539], Fresh[26538], Fresh[26537], Fresh[26536], Fresh[26535], Fresh[26534], Fresh[26533], Fresh[26532], Fresh[26531], Fresh[26530], Fresh[26529], Fresh[26528], Fresh[26527], Fresh[26526], Fresh[26525], Fresh[26524], Fresh[26523], Fresh[26522], Fresh[26521], Fresh[26520], Fresh[26519], Fresh[26518], Fresh[26517], Fresh[26516], Fresh[26515], Fresh[26514], Fresh[26513], Fresh[26512], Fresh[26511], Fresh[26510], Fresh[26509], Fresh[26508], Fresh[26507], Fresh[26506], Fresh[26505], Fresh[26504], Fresh[26503], Fresh[26502], Fresh[26501], Fresh[26500], Fresh[26499], Fresh[26498], Fresh[26497], Fresh[26496], Fresh[26495], Fresh[26494], Fresh[26493], Fresh[26492], Fresh[26491], Fresh[26490], Fresh[26489], Fresh[26488], Fresh[26487], Fresh[26486], Fresh[26485], Fresh[26484], Fresh[26483], Fresh[26482], Fresh[26481], Fresh[26480], Fresh[26479], Fresh[26478], Fresh[26477], Fresh[26476], Fresh[26475], Fresh[26474], Fresh[26473], Fresh[26472], Fresh[26471], Fresh[26470], Fresh[26469], Fresh[26468], Fresh[26467], Fresh[26466], Fresh[26465], Fresh[26464], Fresh[26463], Fresh[26462], Fresh[26461], Fresh[26460], Fresh[26459], Fresh[26458], Fresh[26457], Fresh[26456], Fresh[26455], Fresh[26454], Fresh[26453], Fresh[26452], Fresh[26451], Fresh[26450], Fresh[26449], Fresh[26448], Fresh[26447], Fresh[26446], Fresh[26445], Fresh[26444], Fresh[26443], Fresh[26442], Fresh[26441], Fresh[26440], Fresh[26439], Fresh[26438], Fresh[26437], Fresh[26436], Fresh[26435], Fresh[26434], Fresh[26433], Fresh[26432], Fresh[26431], Fresh[26430], Fresh[26429], Fresh[26428], Fresh[26427], Fresh[26426], Fresh[26425], Fresh[26424], Fresh[26423], Fresh[26422], Fresh[26421], Fresh[26420], Fresh[26419], Fresh[26418], Fresh[26417], Fresh[26416], Fresh[26415], Fresh[26414], Fresh[26413], Fresh[26412], Fresh[26411], Fresh[26410], Fresh[26409], Fresh[26408], Fresh[26407], Fresh[26406], Fresh[26405], Fresh[26404], Fresh[26403], Fresh[26402], Fresh[26401], Fresh[26400], Fresh[26399], Fresh[26398], Fresh[26397], Fresh[26396], Fresh[26395], Fresh[26394], Fresh[26393], Fresh[26392], Fresh[26391], Fresh[26390], Fresh[26389], Fresh[26388], Fresh[26387], Fresh[26386], Fresh[26385], Fresh[26384], Fresh[26383], Fresh[26382], Fresh[26381], Fresh[26380], Fresh[26379], Fresh[26378], Fresh[26377], Fresh[26376], Fresh[26375], Fresh[26374], Fresh[26373], Fresh[26372], Fresh[26371], Fresh[26370], Fresh[26369], Fresh[26368], Fresh[26367], Fresh[26366], Fresh[26365], Fresh[26364], Fresh[26363], Fresh[26362], Fresh[26361], Fresh[26360], Fresh[26359], Fresh[26358], Fresh[26357], Fresh[26356], Fresh[26355], Fresh[26354], Fresh[26353], Fresh[26352], Fresh[26351], Fresh[26350], Fresh[26349], Fresh[26348], Fresh[26347], Fresh[26346], Fresh[26345], Fresh[26344], Fresh[26343], Fresh[26342], Fresh[26341], Fresh[26340], Fresh[26339], Fresh[26338], Fresh[26337], Fresh[26336], Fresh[26335], Fresh[26334], Fresh[26333], Fresh[26332], Fresh[26331], Fresh[26330], Fresh[26329], Fresh[26328], Fresh[26327], Fresh[26326], Fresh[26325], Fresh[26324], Fresh[26323], Fresh[26322], Fresh[26321], Fresh[26320], Fresh[26319], Fresh[26318], Fresh[26317], Fresh[26316], Fresh[26315], Fresh[26314], Fresh[26313], Fresh[26312], Fresh[26311], Fresh[26310], Fresh[26309], Fresh[26308], Fresh[26307], Fresh[26306], Fresh[26305], Fresh[26304], Fresh[26303], Fresh[26302], Fresh[26301], Fresh[26300], Fresh[26299], Fresh[26298], Fresh[26297], Fresh[26296], Fresh[26295], Fresh[26294], Fresh[26293], Fresh[26292], Fresh[26291], Fresh[26290], Fresh[26289], Fresh[26288], Fresh[26287], Fresh[26286], Fresh[26285], Fresh[26284], Fresh[26283], Fresh[26282], Fresh[26281], Fresh[26280], Fresh[26279], Fresh[26278], Fresh[26277], Fresh[26276], Fresh[26275], Fresh[26274], Fresh[26273], Fresh[26272], Fresh[26271], Fresh[26270], Fresh[26269], Fresh[26268], Fresh[26267], Fresh[26266], Fresh[26265], Fresh[26264], Fresh[26263], Fresh[26262], Fresh[26261], Fresh[26260], Fresh[26259], Fresh[26258], Fresh[26257], Fresh[26256], Fresh[26255], Fresh[26254], Fresh[26253], Fresh[26252], Fresh[26251], Fresh[26250], Fresh[26249], Fresh[26248], Fresh[26247], Fresh[26246], Fresh[26245], Fresh[26244], Fresh[26243], Fresh[26242], Fresh[26241], Fresh[26240], Fresh[26239], Fresh[26238], Fresh[26237], Fresh[26236], Fresh[26235], Fresh[26234], Fresh[26233], Fresh[26232], Fresh[26231], Fresh[26230], Fresh[26229], Fresh[26228], Fresh[26227], Fresh[26226], Fresh[26225], Fresh[26224], Fresh[26223], Fresh[26222], Fresh[26221], Fresh[26220], Fresh[26219], Fresh[26218], Fresh[26217], Fresh[26216], Fresh[26215], Fresh[26214], Fresh[26213], Fresh[26212], Fresh[26211], Fresh[26210], Fresh[26209], Fresh[26208], Fresh[26207], Fresh[26206], Fresh[26205], Fresh[26204], Fresh[26203], Fresh[26202], Fresh[26201], Fresh[26200], Fresh[26199], Fresh[26198], Fresh[26197], Fresh[26196], Fresh[26195], Fresh[26194], Fresh[26193], Fresh[26192], Fresh[26191], Fresh[26190], Fresh[26189], Fresh[26188], Fresh[26187], Fresh[26186], Fresh[26185], Fresh[26184], Fresh[26183], Fresh[26182], Fresh[26181], Fresh[26180], Fresh[26179], Fresh[26178], Fresh[26177], Fresh[26176], Fresh[26175], Fresh[26174], Fresh[26173], Fresh[26172], Fresh[26171], Fresh[26170], Fresh[26169], Fresh[26168], Fresh[26167], Fresh[26166], Fresh[26165], Fresh[26164], Fresh[26163], Fresh[26162], Fresh[26161], Fresh[26160], Fresh[26159], Fresh[26158], Fresh[26157], Fresh[26156], Fresh[26155], Fresh[26154], Fresh[26153], Fresh[26152], Fresh[26151], Fresh[26150], Fresh[26149], Fresh[26148], Fresh[26147], Fresh[26146], Fresh[26145], Fresh[26144], Fresh[26143], Fresh[26142], Fresh[26141], Fresh[26140], Fresh[26139], Fresh[26138], Fresh[26137], Fresh[26136], Fresh[26135], Fresh[26134], Fresh[26133], Fresh[26132], Fresh[26131], Fresh[26130], Fresh[26129], Fresh[26128], Fresh[26127], Fresh[26126], Fresh[26125], Fresh[26124], Fresh[26123], Fresh[26122], Fresh[26121], Fresh[26120], Fresh[26119], Fresh[26118], Fresh[26117], Fresh[26116], Fresh[26115], Fresh[26114], Fresh[26113], Fresh[26112], Fresh[26111], Fresh[26110], Fresh[26109], Fresh[26108], Fresh[26107], Fresh[26106], Fresh[26105], Fresh[26104], Fresh[26103], Fresh[26102], Fresh[26101], Fresh[26100], Fresh[26099], Fresh[26098], Fresh[26097], Fresh[26096], Fresh[26095], Fresh[26094], Fresh[26093], Fresh[26092], Fresh[26091], Fresh[26090], Fresh[26089], Fresh[26088], Fresh[26087], Fresh[26086], Fresh[26085], Fresh[26084], Fresh[26083], Fresh[26082], Fresh[26081], Fresh[26080], Fresh[26079], Fresh[26078], Fresh[26077], Fresh[26076], Fresh[26075], Fresh[26074], Fresh[26073], Fresh[26072], Fresh[26071], Fresh[26070], Fresh[26069], Fresh[26068], Fresh[26067], Fresh[26066], Fresh[26065], Fresh[26064], Fresh[26063], Fresh[26062], Fresh[26061], Fresh[26060], Fresh[26059], Fresh[26058], Fresh[26057], Fresh[26056], Fresh[26055], Fresh[26054], Fresh[26053], Fresh[26052], Fresh[26051], Fresh[26050], Fresh[26049], Fresh[26048], Fresh[26047], Fresh[26046], Fresh[26045], Fresh[26044], Fresh[26043], Fresh[26042], Fresh[26041], Fresh[26040], Fresh[26039], Fresh[26038], Fresh[26037], Fresh[26036], Fresh[26035], Fresh[26034], Fresh[26033], Fresh[26032], Fresh[26031], Fresh[26030], Fresh[26029], Fresh[26028], Fresh[26027], Fresh[26026], Fresh[26025], Fresh[26024], Fresh[26023], Fresh[26022], Fresh[26021], Fresh[26020], Fresh[26019], Fresh[26018], Fresh[26017], Fresh[26016], Fresh[26015], Fresh[26014], Fresh[26013], Fresh[26012], Fresh[26011], Fresh[26010], Fresh[26009], Fresh[26008], Fresh[26007], Fresh[26006], Fresh[26005], Fresh[26004], Fresh[26003], Fresh[26002], Fresh[26001], Fresh[26000], Fresh[25999], Fresh[25998], Fresh[25997], Fresh[25996], Fresh[25995], Fresh[25994], Fresh[25993], Fresh[25992], Fresh[25991], Fresh[25990], Fresh[25989], Fresh[25988], Fresh[25987], Fresh[25986], Fresh[25985], Fresh[25984], Fresh[25983], Fresh[25982], Fresh[25981], Fresh[25980], Fresh[25979], Fresh[25978], Fresh[25977], Fresh[25976], Fresh[25975], Fresh[25974], Fresh[25973], Fresh[25972], Fresh[25971], Fresh[25970], Fresh[25969], Fresh[25968], Fresh[25967], Fresh[25966], Fresh[25965], Fresh[25964], Fresh[25963], Fresh[25962], Fresh[25961], Fresh[25960], Fresh[25959], Fresh[25958], Fresh[25957], Fresh[25956], Fresh[25955], Fresh[25954], Fresh[25953], Fresh[25952], Fresh[25951], Fresh[25950], Fresh[25949], Fresh[25948], Fresh[25947], Fresh[25946], Fresh[25945], Fresh[25944], Fresh[25943], Fresh[25942], Fresh[25941], Fresh[25940], Fresh[25939], Fresh[25938], Fresh[25937], Fresh[25936], Fresh[25935], Fresh[25934], Fresh[25933], Fresh[25932], Fresh[25931], Fresh[25930], Fresh[25929], Fresh[25928], Fresh[25927], Fresh[25926], Fresh[25925], Fresh[25924], Fresh[25923], Fresh[25922], Fresh[25921], Fresh[25920], Fresh[25919], Fresh[25918], Fresh[25917], Fresh[25916], Fresh[25915], Fresh[25914], Fresh[25913], Fresh[25912], Fresh[25911], Fresh[25910], Fresh[25909], Fresh[25908], Fresh[25907], Fresh[25906], Fresh[25905], Fresh[25904], Fresh[25903], Fresh[25902], Fresh[25901], Fresh[25900], Fresh[25899], Fresh[25898], Fresh[25897], Fresh[25896], Fresh[25895], Fresh[25894], Fresh[25893], Fresh[25892], Fresh[25891], Fresh[25890], Fresh[25889], Fresh[25888], Fresh[25887], Fresh[25886], Fresh[25885], Fresh[25884], Fresh[25883], Fresh[25882], Fresh[25881], Fresh[25880], Fresh[25879], Fresh[25878], Fresh[25877], Fresh[25876], Fresh[25875], Fresh[25874], Fresh[25873], Fresh[25872], Fresh[25871], Fresh[25870], Fresh[25869], Fresh[25868], Fresh[25867], Fresh[25866], Fresh[25865], Fresh[25864], Fresh[25863], Fresh[25862], Fresh[25861], Fresh[25860], Fresh[25859], Fresh[25858], Fresh[25857], Fresh[25856], Fresh[25855], Fresh[25854], Fresh[25853], Fresh[25852], Fresh[25851], Fresh[25850], Fresh[25849], Fresh[25848], Fresh[25847], Fresh[25846], Fresh[25845], Fresh[25844], Fresh[25843], Fresh[25842], Fresh[25841], Fresh[25840], Fresh[25839], Fresh[25838], Fresh[25837], Fresh[25836], Fresh[25835], Fresh[25834], Fresh[25833], Fresh[25832], Fresh[25831], Fresh[25830], Fresh[25829], Fresh[25828], Fresh[25827], Fresh[25826], Fresh[25825], Fresh[25824], Fresh[25823], Fresh[25822], Fresh[25821], Fresh[25820], Fresh[25819], Fresh[25818], Fresh[25817], Fresh[25816], Fresh[25815], Fresh[25814], Fresh[25813], Fresh[25812], Fresh[25811], Fresh[25810], Fresh[25809], Fresh[25808], Fresh[25807], Fresh[25806], Fresh[25805], Fresh[25804], Fresh[25803], Fresh[25802], Fresh[25801], Fresh[25800], Fresh[25799], Fresh[25798], Fresh[25797], Fresh[25796], Fresh[25795], Fresh[25794], Fresh[25793], Fresh[25792], Fresh[25791], Fresh[25790], Fresh[25789], Fresh[25788], Fresh[25787], Fresh[25786], Fresh[25785], Fresh[25784], Fresh[25783], Fresh[25782], Fresh[25781], Fresh[25780], Fresh[25779], Fresh[25778], Fresh[25777], Fresh[25776], Fresh[25775], Fresh[25774], Fresh[25773], Fresh[25772], Fresh[25771], Fresh[25770], Fresh[25769], Fresh[25768], Fresh[25767], Fresh[25766], Fresh[25765], Fresh[25764], Fresh[25763], Fresh[25762], Fresh[25761], Fresh[25760], Fresh[25759], Fresh[25758], Fresh[25757], Fresh[25756], Fresh[25755], Fresh[25754], Fresh[25753], Fresh[25752], Fresh[25751], Fresh[25750], Fresh[25749], Fresh[25748], Fresh[25747], Fresh[25746], Fresh[25745], Fresh[25744], Fresh[25743], Fresh[25742], Fresh[25741], Fresh[25740], Fresh[25739], Fresh[25738], Fresh[25737], Fresh[25736], Fresh[25735], Fresh[25734], Fresh[25733], Fresh[25732], Fresh[25731], Fresh[25730], Fresh[25729], Fresh[25728], Fresh[25727], Fresh[25726], Fresh[25725], Fresh[25724], Fresh[25723], Fresh[25722], Fresh[25721], Fresh[25720], Fresh[25719], Fresh[25718], Fresh[25717], Fresh[25716], Fresh[25715], Fresh[25714], Fresh[25713], Fresh[25712], Fresh[25711], Fresh[25710], Fresh[25709], Fresh[25708], Fresh[25707], Fresh[25706], Fresh[25705], Fresh[25704], Fresh[25703], Fresh[25702], Fresh[25701], Fresh[25700], Fresh[25699], Fresh[25698], Fresh[25697], Fresh[25696], Fresh[25695], Fresh[25694], Fresh[25693], Fresh[25692], Fresh[25691], Fresh[25690], Fresh[25689], Fresh[25688], Fresh[25687], Fresh[25686], Fresh[25685], Fresh[25684], Fresh[25683], Fresh[25682], Fresh[25681], Fresh[25680], Fresh[25679], Fresh[25678], Fresh[25677], Fresh[25676], Fresh[25675], Fresh[25674], Fresh[25673], Fresh[25672], Fresh[25671], Fresh[25670], Fresh[25669], Fresh[25668], Fresh[25667], Fresh[25666], Fresh[25665], Fresh[25664], Fresh[25663], Fresh[25662], Fresh[25661], Fresh[25660], Fresh[25659], Fresh[25658], Fresh[25657], Fresh[25656], Fresh[25655], Fresh[25654], Fresh[25653], Fresh[25652], Fresh[25651], Fresh[25650], Fresh[25649], Fresh[25648], Fresh[25647], Fresh[25646], Fresh[25645], Fresh[25644], Fresh[25643], Fresh[25642], Fresh[25641], Fresh[25640], Fresh[25639], Fresh[25638], Fresh[25637], Fresh[25636], Fresh[25635], Fresh[25634], Fresh[25633], Fresh[25632], Fresh[25631], Fresh[25630], Fresh[25629], Fresh[25628], Fresh[25627], Fresh[25626], Fresh[25625], Fresh[25624], Fresh[25623], Fresh[25622], Fresh[25621], Fresh[25620], Fresh[25619], Fresh[25618], Fresh[25617], Fresh[25616], Fresh[25615], Fresh[25614], Fresh[25613], Fresh[25612], Fresh[25611], Fresh[25610], Fresh[25609], Fresh[25608], Fresh[25607], Fresh[25606], Fresh[25605], Fresh[25604], Fresh[25603], Fresh[25602], Fresh[25601], Fresh[25600], Fresh[25599], Fresh[25598], Fresh[25597], Fresh[25596], Fresh[25595], Fresh[25594], Fresh[25593], Fresh[25592], Fresh[25591], Fresh[25590], Fresh[25589], Fresh[25588], Fresh[25587], Fresh[25586], Fresh[25585], Fresh[25584], Fresh[25583], Fresh[25582], Fresh[25581], Fresh[25580], Fresh[25579], Fresh[25578], Fresh[25577], Fresh[25576], Fresh[25575], Fresh[25574], Fresh[25573], Fresh[25572], Fresh[25571], Fresh[25570], Fresh[25569], Fresh[25568], Fresh[25567], Fresh[25566], Fresh[25565], Fresh[25564], Fresh[25563], Fresh[25562], Fresh[25561], Fresh[25560], Fresh[25559], Fresh[25558], Fresh[25557], Fresh[25556], Fresh[25555], Fresh[25554], Fresh[25553], Fresh[25552], Fresh[25551], Fresh[25550], Fresh[25549], Fresh[25548], Fresh[25547], Fresh[25546], Fresh[25545], Fresh[25544], Fresh[25543], Fresh[25542], Fresh[25541], Fresh[25540], Fresh[25539], Fresh[25538], Fresh[25537], Fresh[25536], Fresh[25535], Fresh[25534], Fresh[25533], Fresh[25532], Fresh[25531], Fresh[25530], Fresh[25529], Fresh[25528], Fresh[25527], Fresh[25526], Fresh[25525], Fresh[25524], Fresh[25523], Fresh[25522], Fresh[25521], Fresh[25520], Fresh[25519], Fresh[25518], Fresh[25517], Fresh[25516], Fresh[25515], Fresh[25514], Fresh[25513], Fresh[25512], Fresh[25511], Fresh[25510], Fresh[25509], Fresh[25508], Fresh[25507], Fresh[25506], Fresh[25505], Fresh[25504], Fresh[25503], Fresh[25502], Fresh[25501], Fresh[25500], Fresh[25499], Fresh[25498], Fresh[25497], Fresh[25496], Fresh[25495], Fresh[25494], Fresh[25493], Fresh[25492], Fresh[25491], Fresh[25490], Fresh[25489], Fresh[25488], Fresh[25487], Fresh[25486], Fresh[25485], Fresh[25484], Fresh[25483], Fresh[25482], Fresh[25481], Fresh[25480], Fresh[25479], Fresh[25478], Fresh[25477], Fresh[25476], Fresh[25475], Fresh[25474], Fresh[25473], Fresh[25472], Fresh[25471], Fresh[25470], Fresh[25469], Fresh[25468], Fresh[25467], Fresh[25466], Fresh[25465], Fresh[25464], Fresh[25463], Fresh[25462], Fresh[25461], Fresh[25460], Fresh[25459], Fresh[25458], Fresh[25457], Fresh[25456], Fresh[25455], Fresh[25454], Fresh[25453], Fresh[25452], Fresh[25451], Fresh[25450], Fresh[25449], Fresh[25448], Fresh[25447], Fresh[25446], Fresh[25445], Fresh[25444], Fresh[25443], Fresh[25442], Fresh[25441], Fresh[25440], Fresh[25439], Fresh[25438], Fresh[25437], Fresh[25436], Fresh[25435], Fresh[25434], Fresh[25433], Fresh[25432], Fresh[25431], Fresh[25430], Fresh[25429], Fresh[25428], Fresh[25427], Fresh[25426], Fresh[25425], Fresh[25424], Fresh[25423], Fresh[25422], Fresh[25421], Fresh[25420], Fresh[25419], Fresh[25418], Fresh[25417], Fresh[25416], Fresh[25415], Fresh[25414], Fresh[25413], Fresh[25412], Fresh[25411], Fresh[25410], Fresh[25409], Fresh[25408], Fresh[25407], Fresh[25406], Fresh[25405], Fresh[25404], Fresh[25403], Fresh[25402], Fresh[25401], Fresh[25400], Fresh[25399], Fresh[25398], Fresh[25397], Fresh[25396], Fresh[25395], Fresh[25394], Fresh[25393], Fresh[25392], Fresh[25391], Fresh[25390], Fresh[25389], Fresh[25388], Fresh[25387], Fresh[25386], Fresh[25385], Fresh[25384], Fresh[25383], Fresh[25382], Fresh[25381], Fresh[25380], Fresh[25379], Fresh[25378], Fresh[25377], Fresh[25376], Fresh[25375], Fresh[25374], Fresh[25373], Fresh[25372], Fresh[25371], Fresh[25370], Fresh[25369], Fresh[25368], Fresh[25367], Fresh[25366], Fresh[25365], Fresh[25364], Fresh[25363], Fresh[25362], Fresh[25361], Fresh[25360], Fresh[25359], Fresh[25358], Fresh[25357], Fresh[25356], Fresh[25355], Fresh[25354], Fresh[25353], Fresh[25352], Fresh[25351], Fresh[25350], Fresh[25349], Fresh[25348], Fresh[25347], Fresh[25346], Fresh[25345], Fresh[25344], Fresh[25343], Fresh[25342], Fresh[25341], Fresh[25340], Fresh[25339], Fresh[25338], Fresh[25337], Fresh[25336], Fresh[25335], Fresh[25334], Fresh[25333], Fresh[25332], Fresh[25331], Fresh[25330], Fresh[25329], Fresh[25328], Fresh[25327], Fresh[25326], Fresh[25325], Fresh[25324], Fresh[25323], Fresh[25322], Fresh[25321], Fresh[25320], Fresh[25319], Fresh[25318], Fresh[25317], Fresh[25316], Fresh[25315], Fresh[25314], Fresh[25313], Fresh[25312], Fresh[25311], Fresh[25310], Fresh[25309], Fresh[25308], Fresh[25307], Fresh[25306], Fresh[25305], Fresh[25304], Fresh[25303], Fresh[25302], Fresh[25301], Fresh[25300], Fresh[25299], Fresh[25298], Fresh[25297], Fresh[25296], Fresh[25295], Fresh[25294], Fresh[25293], Fresh[25292], Fresh[25291], Fresh[25290], Fresh[25289], Fresh[25288], Fresh[25287], Fresh[25286], Fresh[25285], Fresh[25284], Fresh[25283], Fresh[25282], Fresh[25281], Fresh[25280], Fresh[25279], Fresh[25278], Fresh[25277], Fresh[25276], Fresh[25275], Fresh[25274], Fresh[25273], Fresh[25272], Fresh[25271], Fresh[25270], Fresh[25269], Fresh[25268], Fresh[25267], Fresh[25266], Fresh[25265], Fresh[25264], Fresh[25263], Fresh[25262], Fresh[25261], Fresh[25260], Fresh[25259], Fresh[25258], Fresh[25257], Fresh[25256], Fresh[25255], Fresh[25254], Fresh[25253], Fresh[25252], Fresh[25251], Fresh[25250], Fresh[25249], Fresh[25248], Fresh[25247], Fresh[25246], Fresh[25245], Fresh[25244], Fresh[25243], Fresh[25242], Fresh[25241], Fresh[25240], Fresh[25239], Fresh[25238], Fresh[25237], Fresh[25236], Fresh[25235], Fresh[25234], Fresh[25233], Fresh[25232], Fresh[25231], Fresh[25230], Fresh[25229], Fresh[25228], Fresh[25227], Fresh[25226], Fresh[25225], Fresh[25224], Fresh[25223], Fresh[25222], Fresh[25221], Fresh[25220], Fresh[25219], Fresh[25218], Fresh[25217], Fresh[25216], Fresh[25215], Fresh[25214], Fresh[25213], Fresh[25212], Fresh[25211], Fresh[25210], Fresh[25209], Fresh[25208], Fresh[25207], Fresh[25206], Fresh[25205], Fresh[25204], Fresh[25203], Fresh[25202], Fresh[25201], Fresh[25200], Fresh[25199], Fresh[25198], Fresh[25197], Fresh[25196], Fresh[25195], Fresh[25194], Fresh[25193], Fresh[25192], Fresh[25191], Fresh[25190], Fresh[25189], Fresh[25188], Fresh[25187], Fresh[25186], Fresh[25185], Fresh[25184], Fresh[25183], Fresh[25182], Fresh[25181], Fresh[25180], Fresh[25179], Fresh[25178], Fresh[25177], Fresh[25176], Fresh[25175], Fresh[25174], Fresh[25173], Fresh[25172], Fresh[25171], Fresh[25170], Fresh[25169], Fresh[25168], Fresh[25167], Fresh[25166], Fresh[25165], Fresh[25164], Fresh[25163], Fresh[25162], Fresh[25161], Fresh[25160], Fresh[25159], Fresh[25158], Fresh[25157], Fresh[25156], Fresh[25155], Fresh[25154], Fresh[25153], Fresh[25152], Fresh[25151], Fresh[25150], Fresh[25149], Fresh[25148], Fresh[25147], Fresh[25146], Fresh[25145], Fresh[25144], Fresh[25143], Fresh[25142], Fresh[25141], Fresh[25140], Fresh[25139], Fresh[25138], Fresh[25137], Fresh[25136], Fresh[25135], Fresh[25134], Fresh[25133], Fresh[25132], Fresh[25131], Fresh[25130], Fresh[25129], Fresh[25128], Fresh[25127], Fresh[25126], Fresh[25125], Fresh[25124], Fresh[25123], Fresh[25122], Fresh[25121], Fresh[25120], Fresh[25119], Fresh[25118], Fresh[25117], Fresh[25116], Fresh[25115], Fresh[25114], Fresh[25113], Fresh[25112], Fresh[25111], Fresh[25110], Fresh[25109], Fresh[25108], Fresh[25107], Fresh[25106], Fresh[25105], Fresh[25104], Fresh[25103], Fresh[25102], Fresh[25101], Fresh[25100], Fresh[25099], Fresh[25098], Fresh[25097], Fresh[25096], Fresh[25095], Fresh[25094], Fresh[25093], Fresh[25092], Fresh[25091], Fresh[25090], Fresh[25089], Fresh[25088], Fresh[25087], Fresh[25086], Fresh[25085], Fresh[25084], Fresh[25083], Fresh[25082], Fresh[25081], Fresh[25080], Fresh[25079], Fresh[25078], Fresh[25077], Fresh[25076], Fresh[25075], Fresh[25074], Fresh[25073], Fresh[25072], Fresh[25071], Fresh[25070], Fresh[25069], Fresh[25068], Fresh[25067], Fresh[25066], Fresh[25065], Fresh[25064], Fresh[25063], Fresh[25062], Fresh[25061], Fresh[25060], Fresh[25059], Fresh[25058], Fresh[25057], Fresh[25056], Fresh[25055], Fresh[25054], Fresh[25053], Fresh[25052], Fresh[25051], Fresh[25050], Fresh[25049], Fresh[25048], Fresh[25047], Fresh[25046], Fresh[25045], Fresh[25044], Fresh[25043], Fresh[25042], Fresh[25041], Fresh[25040], Fresh[25039], Fresh[25038], Fresh[25037], Fresh[25036], Fresh[25035], Fresh[25034], Fresh[25033], Fresh[25032], Fresh[25031], Fresh[25030], Fresh[25029], Fresh[25028], Fresh[25027], Fresh[25026], Fresh[25025], Fresh[25024], Fresh[25023], Fresh[25022], Fresh[25021], Fresh[25020], Fresh[25019], Fresh[25018], Fresh[25017], Fresh[25016], Fresh[25015], Fresh[25014], Fresh[25013], Fresh[25012], Fresh[25011], Fresh[25010], Fresh[25009], Fresh[25008], Fresh[25007], Fresh[25006], Fresh[25005], Fresh[25004], Fresh[25003], Fresh[25002], Fresh[25001], Fresh[25000], Fresh[24999], Fresh[24998], Fresh[24997], Fresh[24996], Fresh[24995], Fresh[24994], Fresh[24993], Fresh[24992], Fresh[24991], Fresh[24990], Fresh[24989], Fresh[24988], Fresh[24987], Fresh[24986], Fresh[24985], Fresh[24984], Fresh[24983], Fresh[24982], Fresh[24981], Fresh[24980], Fresh[24979], Fresh[24978], Fresh[24977], Fresh[24976], Fresh[24975], Fresh[24974], Fresh[24973], Fresh[24972], Fresh[24971], Fresh[24970], Fresh[24969], Fresh[24968], Fresh[24967], Fresh[24966], Fresh[24965], Fresh[24964], Fresh[24963], Fresh[24962], Fresh[24961], Fresh[24960], Fresh[24959], Fresh[24958], Fresh[24957], Fresh[24956], Fresh[24955], Fresh[24954], Fresh[24953], Fresh[24952], Fresh[24951], Fresh[24950], Fresh[24949], Fresh[24948], Fresh[24947], Fresh[24946], Fresh[24945], Fresh[24944], Fresh[24943], Fresh[24942], Fresh[24941], Fresh[24940], Fresh[24939], Fresh[24938], Fresh[24937], Fresh[24936], Fresh[24935], Fresh[24934], Fresh[24933], Fresh[24932], Fresh[24931], Fresh[24930], Fresh[24929], Fresh[24928], Fresh[24927], Fresh[24926], Fresh[24925], Fresh[24924], Fresh[24923], Fresh[24922], Fresh[24921], Fresh[24920], Fresh[24919], Fresh[24918], Fresh[24917], Fresh[24916], Fresh[24915], Fresh[24914], Fresh[24913], Fresh[24912], Fresh[24911], Fresh[24910], Fresh[24909], Fresh[24908], Fresh[24907], Fresh[24906], Fresh[24905], Fresh[24904], Fresh[24903], Fresh[24902], Fresh[24901], Fresh[24900], Fresh[24899], Fresh[24898], Fresh[24897], Fresh[24896], Fresh[24895], Fresh[24894], Fresh[24893], Fresh[24892], Fresh[24891], Fresh[24890], Fresh[24889], Fresh[24888], Fresh[24887], Fresh[24886], Fresh[24885], Fresh[24884], Fresh[24883], Fresh[24882], Fresh[24881], Fresh[24880], Fresh[24879], Fresh[24878], Fresh[24877], Fresh[24876], Fresh[24875], Fresh[24874], Fresh[24873], Fresh[24872], Fresh[24871], Fresh[24870], Fresh[24869], Fresh[24868], Fresh[24867], Fresh[24866], Fresh[24865], Fresh[24864], Fresh[24863], Fresh[24862], Fresh[24861], Fresh[24860], Fresh[24859], Fresh[24858], Fresh[24857], Fresh[24856], Fresh[24855], Fresh[24854], Fresh[24853], Fresh[24852], Fresh[24851], Fresh[24850], Fresh[24849], Fresh[24848], Fresh[24847], Fresh[24846], Fresh[24845], Fresh[24844], Fresh[24843], Fresh[24842], Fresh[24841], Fresh[24840], Fresh[24839], Fresh[24838], Fresh[24837], Fresh[24836], Fresh[24835], Fresh[24834], Fresh[24833], Fresh[24832], Fresh[24831], Fresh[24830], Fresh[24829], Fresh[24828], Fresh[24827], Fresh[24826], Fresh[24825], Fresh[24824], Fresh[24823], Fresh[24822], Fresh[24821], Fresh[24820], Fresh[24819], Fresh[24818], Fresh[24817], Fresh[24816], Fresh[24815], Fresh[24814], Fresh[24813], Fresh[24812], Fresh[24811], Fresh[24810], Fresh[24809], Fresh[24808], Fresh[24807], Fresh[24806], Fresh[24805], Fresh[24804], Fresh[24803], Fresh[24802], Fresh[24801], Fresh[24800], Fresh[24799], Fresh[24798], Fresh[24797], Fresh[24796], Fresh[24795], Fresh[24794], Fresh[24793], Fresh[24792], Fresh[24791], Fresh[24790], Fresh[24789], Fresh[24788], Fresh[24787], Fresh[24786], Fresh[24785], Fresh[24784], Fresh[24783], Fresh[24782], Fresh[24781], Fresh[24780], Fresh[24779], Fresh[24778], Fresh[24777], Fresh[24776], Fresh[24775], Fresh[24774], Fresh[24773], Fresh[24772], Fresh[24771], Fresh[24770], Fresh[24769], Fresh[24768], Fresh[24767], Fresh[24766], Fresh[24765], Fresh[24764], Fresh[24763], Fresh[24762], Fresh[24761], Fresh[24760], Fresh[24759], Fresh[24758], Fresh[24757], Fresh[24756], Fresh[24755], Fresh[24754], Fresh[24753], Fresh[24752], Fresh[24751], Fresh[24750], Fresh[24749], Fresh[24748], Fresh[24747], Fresh[24746], Fresh[24745], Fresh[24744], Fresh[24743], Fresh[24742], Fresh[24741], Fresh[24740], Fresh[24739], Fresh[24738], Fresh[24737], Fresh[24736], Fresh[24735], Fresh[24734], Fresh[24733], Fresh[24732], Fresh[24731], Fresh[24730], Fresh[24729], Fresh[24728], Fresh[24727], Fresh[24726], Fresh[24725], Fresh[24724], Fresh[24723], Fresh[24722], Fresh[24721], Fresh[24720], Fresh[24719], Fresh[24718], Fresh[24717], Fresh[24716], Fresh[24715], Fresh[24714], Fresh[24713], Fresh[24712], Fresh[24711], Fresh[24710], Fresh[24709], Fresh[24708], Fresh[24707], Fresh[24706], Fresh[24705], Fresh[24704], Fresh[24703], Fresh[24702], Fresh[24701], Fresh[24700], Fresh[24699], Fresh[24698], Fresh[24697], Fresh[24696], Fresh[24695], Fresh[24694], Fresh[24693], Fresh[24692], Fresh[24691], Fresh[24690], Fresh[24689], Fresh[24688], Fresh[24687], Fresh[24686], Fresh[24685], Fresh[24684], Fresh[24683], Fresh[24682], Fresh[24681], Fresh[24680], Fresh[24679], Fresh[24678], Fresh[24677], Fresh[24676], Fresh[24675], Fresh[24674], Fresh[24673], Fresh[24672], Fresh[24671], Fresh[24670], Fresh[24669], Fresh[24668], Fresh[24667], Fresh[24666], Fresh[24665], Fresh[24664], Fresh[24663], Fresh[24662], Fresh[24661], Fresh[24660], Fresh[24659], Fresh[24658], Fresh[24657], Fresh[24656], Fresh[24655], Fresh[24654], Fresh[24653], Fresh[24652], Fresh[24651], Fresh[24650], Fresh[24649], Fresh[24648], Fresh[24647], Fresh[24646], Fresh[24645], Fresh[24644], Fresh[24643], Fresh[24642], Fresh[24641], Fresh[24640], Fresh[24639], Fresh[24638], Fresh[24637], Fresh[24636], Fresh[24635], Fresh[24634], Fresh[24633], Fresh[24632], Fresh[24631], Fresh[24630], Fresh[24629], Fresh[24628], Fresh[24627], Fresh[24626], Fresh[24625], Fresh[24624], Fresh[24623], Fresh[24622], Fresh[24621], Fresh[24620], Fresh[24619], Fresh[24618], Fresh[24617], Fresh[24616], Fresh[24615], Fresh[24614], Fresh[24613], Fresh[24612], Fresh[24611], Fresh[24610], Fresh[24609], Fresh[24608], Fresh[24607], Fresh[24606], Fresh[24605], Fresh[24604], Fresh[24603], Fresh[24602], Fresh[24601], Fresh[24600], Fresh[24599], Fresh[24598], Fresh[24597], Fresh[24596], Fresh[24595], Fresh[24594], Fresh[24593], Fresh[24592], Fresh[24591], Fresh[24590], Fresh[24589], Fresh[24588], Fresh[24587], Fresh[24586], Fresh[24585], Fresh[24584], Fresh[24583], Fresh[24582], Fresh[24581], Fresh[24580], Fresh[24579], Fresh[24578], Fresh[24577], Fresh[24576], Fresh[24575], Fresh[24574], Fresh[24573], Fresh[24572], Fresh[24571], Fresh[24570], Fresh[24569], Fresh[24568], Fresh[24567], Fresh[24566], Fresh[24565], Fresh[24564], Fresh[24563], Fresh[24562], Fresh[24561], Fresh[24560], Fresh[24559], Fresh[24558], Fresh[24557], Fresh[24556], Fresh[24555], Fresh[24554], Fresh[24553], Fresh[24552], Fresh[24551], Fresh[24550], Fresh[24549], Fresh[24548], Fresh[24547], Fresh[24546], Fresh[24545], Fresh[24544], Fresh[24543], Fresh[24542], Fresh[24541], Fresh[24540], Fresh[24539], Fresh[24538], Fresh[24537], Fresh[24536], Fresh[24535], Fresh[24534], Fresh[24533], Fresh[24532], Fresh[24531], Fresh[24530], Fresh[24529], Fresh[24528], Fresh[24527], Fresh[24526], Fresh[24525], Fresh[24524], Fresh[24523], Fresh[24522], Fresh[24521], Fresh[24520], Fresh[24519], Fresh[24518], Fresh[24517], Fresh[24516], Fresh[24515], Fresh[24514], Fresh[24513], Fresh[24512], Fresh[24511], Fresh[24510], Fresh[24509], Fresh[24508], Fresh[24507], Fresh[24506], Fresh[24505], Fresh[24504], Fresh[24503], Fresh[24502], Fresh[24501], Fresh[24500], Fresh[24499], Fresh[24498], Fresh[24497], Fresh[24496], Fresh[24495], Fresh[24494], Fresh[24493], Fresh[24492], Fresh[24491], Fresh[24490], Fresh[24489], Fresh[24488], Fresh[24487], Fresh[24486], Fresh[24485], Fresh[24484], Fresh[24483], Fresh[24482], Fresh[24481], Fresh[24480], Fresh[24479], Fresh[24478], Fresh[24477], Fresh[24476], Fresh[24475], Fresh[24474], Fresh[24473], Fresh[24472], Fresh[24471], Fresh[24470], Fresh[24469], Fresh[24468], Fresh[24467], Fresh[24466], Fresh[24465], Fresh[24464], Fresh[24463], Fresh[24462], Fresh[24461], Fresh[24460], Fresh[24459], Fresh[24458], Fresh[24457], Fresh[24456], Fresh[24455], Fresh[24454], Fresh[24453], Fresh[24452], Fresh[24451], Fresh[24450], Fresh[24449], Fresh[24448], Fresh[24447], Fresh[24446], Fresh[24445], Fresh[24444], Fresh[24443], Fresh[24442], Fresh[24441], Fresh[24440], Fresh[24439], Fresh[24438], Fresh[24437], Fresh[24436], Fresh[24435], Fresh[24434], Fresh[24433], Fresh[24432], Fresh[24431], Fresh[24430], Fresh[24429], Fresh[24428], Fresh[24427], Fresh[24426], Fresh[24425], Fresh[24424], Fresh[24423], Fresh[24422], Fresh[24421], Fresh[24420], Fresh[24419], Fresh[24418], Fresh[24417], Fresh[24416], Fresh[24415], Fresh[24414], Fresh[24413], Fresh[24412], Fresh[24411], Fresh[24410], Fresh[24409], Fresh[24408], Fresh[24407], Fresh[24406], Fresh[24405], Fresh[24404], Fresh[24403], Fresh[24402], Fresh[24401], Fresh[24400], Fresh[24399], Fresh[24398], Fresh[24397], Fresh[24396], Fresh[24395], Fresh[24394], Fresh[24393], Fresh[24392], Fresh[24391], Fresh[24390], Fresh[24389], Fresh[24388], Fresh[24387], Fresh[24386], Fresh[24385], Fresh[24384], Fresh[24383], Fresh[24382], Fresh[24381], Fresh[24380], Fresh[24379], Fresh[24378], Fresh[24377], Fresh[24376], Fresh[24375], Fresh[24374], Fresh[24373], Fresh[24372], Fresh[24371], Fresh[24370], Fresh[24369], Fresh[24368], Fresh[24367], Fresh[24366], Fresh[24365], Fresh[24364], Fresh[24363], Fresh[24362], Fresh[24361], Fresh[24360], Fresh[24359], Fresh[24358], Fresh[24357], Fresh[24356], Fresh[24355], Fresh[24354], Fresh[24353], Fresh[24352], Fresh[24351], Fresh[24350], Fresh[24349], Fresh[24348], Fresh[24347], Fresh[24346], Fresh[24345], Fresh[24344], Fresh[24343], Fresh[24342], Fresh[24341], Fresh[24340], Fresh[24339], Fresh[24338], Fresh[24337], Fresh[24336], Fresh[24335], Fresh[24334], Fresh[24333], Fresh[24332], Fresh[24331], Fresh[24330], Fresh[24329], Fresh[24328], Fresh[24327], Fresh[24326], Fresh[24325], Fresh[24324], Fresh[24323], Fresh[24322], Fresh[24321], Fresh[24320], Fresh[24319], Fresh[24318], Fresh[24317], Fresh[24316], Fresh[24315], Fresh[24314], Fresh[24313], Fresh[24312], Fresh[24311], Fresh[24310], Fresh[24309], Fresh[24308], Fresh[24307], Fresh[24306], Fresh[24305], Fresh[24304], Fresh[24303], Fresh[24302], Fresh[24301], Fresh[24300], Fresh[24299], Fresh[24298], Fresh[24297], Fresh[24296], Fresh[24295], Fresh[24294], Fresh[24293], Fresh[24292], Fresh[24291], Fresh[24290], Fresh[24289], Fresh[24288], Fresh[24287], Fresh[24286], Fresh[24285], Fresh[24284], Fresh[24283], Fresh[24282], Fresh[24281], Fresh[24280], Fresh[24279], Fresh[24278], Fresh[24277], Fresh[24276], Fresh[24275], Fresh[24274], Fresh[24273], Fresh[24272], Fresh[24271], Fresh[24270], Fresh[24269], Fresh[24268], Fresh[24267], Fresh[24266], Fresh[24265], Fresh[24264], Fresh[24263], Fresh[24262], Fresh[24261], Fresh[24260], Fresh[24259], Fresh[24258], Fresh[24257], Fresh[24256], Fresh[24255], Fresh[24254], Fresh[24253], Fresh[24252], Fresh[24251], Fresh[24250], Fresh[24249], Fresh[24248], Fresh[24247], Fresh[24246], Fresh[24245], Fresh[24244], Fresh[24243], Fresh[24242], Fresh[24241], Fresh[24240], Fresh[24239], Fresh[24238], Fresh[24237], Fresh[24236], Fresh[24235], Fresh[24234], Fresh[24233], Fresh[24232], Fresh[24231], Fresh[24230], Fresh[24229], Fresh[24228], Fresh[24227], Fresh[24226], Fresh[24225], Fresh[24224], Fresh[24223], Fresh[24222], Fresh[24221], Fresh[24220], Fresh[24219], Fresh[24218], Fresh[24217], Fresh[24216], Fresh[24215], Fresh[24214], Fresh[24213], Fresh[24212], Fresh[24211], Fresh[24210], Fresh[24209], Fresh[24208], Fresh[24207], Fresh[24206], Fresh[24205], Fresh[24204], Fresh[24203], Fresh[24202], Fresh[24201], Fresh[24200], Fresh[24199], Fresh[24198], Fresh[24197], Fresh[24196], Fresh[24195], Fresh[24194], Fresh[24193], Fresh[24192], Fresh[24191], Fresh[24190], Fresh[24189], Fresh[24188], Fresh[24187], Fresh[24186], Fresh[24185], Fresh[24184], Fresh[24183], Fresh[24182], Fresh[24181], Fresh[24180], Fresh[24179], Fresh[24178], Fresh[24177], Fresh[24176], Fresh[24175], Fresh[24174], Fresh[24173], Fresh[24172], Fresh[24171], Fresh[24170], Fresh[24169], Fresh[24168], Fresh[24167], Fresh[24166], Fresh[24165], Fresh[24164], Fresh[24163], Fresh[24162], Fresh[24161], Fresh[24160], Fresh[24159], Fresh[24158], Fresh[24157], Fresh[24156], Fresh[24155], Fresh[24154], Fresh[24153], Fresh[24152], Fresh[24151], Fresh[24150], Fresh[24149], Fresh[24148], Fresh[24147], Fresh[24146], Fresh[24145], Fresh[24144], Fresh[24143], Fresh[24142], Fresh[24141], Fresh[24140], Fresh[24139], Fresh[24138], Fresh[24137], Fresh[24136], Fresh[24135], Fresh[24134], Fresh[24133], Fresh[24132], Fresh[24131], Fresh[24130], Fresh[24129], Fresh[24128], Fresh[24127], Fresh[24126], Fresh[24125], Fresh[24124], Fresh[24123], Fresh[24122], Fresh[24121], Fresh[24120], Fresh[24119], Fresh[24118], Fresh[24117], Fresh[24116], Fresh[24115], Fresh[24114], Fresh[24113], Fresh[24112], Fresh[24111], Fresh[24110], Fresh[24109], Fresh[24108], Fresh[24107], Fresh[24106], Fresh[24105], Fresh[24104], Fresh[24103], Fresh[24102], Fresh[24101], Fresh[24100], Fresh[24099], Fresh[24098], Fresh[24097], Fresh[24096], Fresh[24095], Fresh[24094], Fresh[24093], Fresh[24092], Fresh[24091], Fresh[24090], Fresh[24089], Fresh[24088], Fresh[24087], Fresh[24086], Fresh[24085], Fresh[24084], Fresh[24083], Fresh[24082], Fresh[24081], Fresh[24080], Fresh[24079], Fresh[24078], Fresh[24077], Fresh[24076], Fresh[24075], Fresh[24074], Fresh[24073], Fresh[24072], Fresh[24071], Fresh[24070], Fresh[24069], Fresh[24068], Fresh[24067], Fresh[24066], Fresh[24065], Fresh[24064], Fresh[24063], Fresh[24062], Fresh[24061], Fresh[24060], Fresh[24059], Fresh[24058], Fresh[24057], Fresh[24056], Fresh[24055], Fresh[24054], Fresh[24053], Fresh[24052], Fresh[24051], Fresh[24050], Fresh[24049], Fresh[24048], Fresh[24047], Fresh[24046], Fresh[24045], Fresh[24044], Fresh[24043], Fresh[24042], Fresh[24041], Fresh[24040], Fresh[24039], Fresh[24038], Fresh[24037], Fresh[24036], Fresh[24035], Fresh[24034], Fresh[24033], Fresh[24032], Fresh[24031], Fresh[24030], Fresh[24029], Fresh[24028], Fresh[24027], Fresh[24026], Fresh[24025], Fresh[24024], Fresh[24023], Fresh[24022], Fresh[24021], Fresh[24020], Fresh[24019], Fresh[24018], Fresh[24017], Fresh[24016], Fresh[24015], Fresh[24014], Fresh[24013], Fresh[24012], Fresh[24011], Fresh[24010], Fresh[24009], Fresh[24008], Fresh[24007], Fresh[24006], Fresh[24005], Fresh[24004], Fresh[24003], Fresh[24002], Fresh[24001], Fresh[24000], Fresh[23999], Fresh[23998], Fresh[23997], Fresh[23996], Fresh[23995], Fresh[23994], Fresh[23993], Fresh[23992], Fresh[23991], Fresh[23990], Fresh[23989], Fresh[23988], Fresh[23987], Fresh[23986], Fresh[23985], Fresh[23984], Fresh[23983], Fresh[23982], Fresh[23981], Fresh[23980], Fresh[23979], Fresh[23978], Fresh[23977], Fresh[23976], Fresh[23975], Fresh[23974], Fresh[23973], Fresh[23972], Fresh[23971], Fresh[23970], Fresh[23969], Fresh[23968], Fresh[23967], Fresh[23966], Fresh[23965], Fresh[23964], Fresh[23963], Fresh[23962], Fresh[23961], Fresh[23960], Fresh[23959], Fresh[23958], Fresh[23957], Fresh[23956], Fresh[23955], Fresh[23954], Fresh[23953], Fresh[23952], Fresh[23951], Fresh[23950], Fresh[23949], Fresh[23948], Fresh[23947], Fresh[23946], Fresh[23945], Fresh[23944], Fresh[23943], Fresh[23942], Fresh[23941], Fresh[23940], Fresh[23939], Fresh[23938], Fresh[23937], Fresh[23936], Fresh[23935], Fresh[23934], Fresh[23933], Fresh[23932], Fresh[23931], Fresh[23930], Fresh[23929], Fresh[23928], Fresh[23927], Fresh[23926], Fresh[23925], Fresh[23924], Fresh[23923], Fresh[23922], Fresh[23921], Fresh[23920], Fresh[23919], Fresh[23918], Fresh[23917], Fresh[23916], Fresh[23915], Fresh[23914], Fresh[23913], Fresh[23912], Fresh[23911], Fresh[23910], Fresh[23909], Fresh[23908], Fresh[23907], Fresh[23906], Fresh[23905], Fresh[23904], Fresh[23903], Fresh[23902], Fresh[23901], Fresh[23900], Fresh[23899], Fresh[23898], Fresh[23897], Fresh[23896], Fresh[23895], Fresh[23894], Fresh[23893], Fresh[23892], Fresh[23891], Fresh[23890], Fresh[23889], Fresh[23888], Fresh[23887], Fresh[23886], Fresh[23885], Fresh[23884], Fresh[23883], Fresh[23882], Fresh[23881], Fresh[23880], Fresh[23879], Fresh[23878], Fresh[23877], Fresh[23876], Fresh[23875], Fresh[23874], Fresh[23873], Fresh[23872], Fresh[23871], Fresh[23870], Fresh[23869], Fresh[23868], Fresh[23867], Fresh[23866], Fresh[23865], Fresh[23864], Fresh[23863], Fresh[23862], Fresh[23861], Fresh[23860], Fresh[23859], Fresh[23858], Fresh[23857], Fresh[23856], Fresh[23855], Fresh[23854], Fresh[23853], Fresh[23852], Fresh[23851], Fresh[23850], Fresh[23849], Fresh[23848], Fresh[23847], Fresh[23846], Fresh[23845], Fresh[23844], Fresh[23843], Fresh[23842], Fresh[23841], Fresh[23840], Fresh[23839], Fresh[23838], Fresh[23837], Fresh[23836], Fresh[23835], Fresh[23834], Fresh[23833], Fresh[23832], Fresh[23831], Fresh[23830], Fresh[23829], Fresh[23828], Fresh[23827], Fresh[23826], Fresh[23825], Fresh[23824], Fresh[23823], Fresh[23822], Fresh[23821], Fresh[23820], Fresh[23819], Fresh[23818], Fresh[23817], Fresh[23816], Fresh[23815], Fresh[23814], Fresh[23813], Fresh[23812], Fresh[23811], Fresh[23810], Fresh[23809], Fresh[23808], Fresh[23807], Fresh[23806], Fresh[23805], Fresh[23804], Fresh[23803], Fresh[23802], Fresh[23801], Fresh[23800], Fresh[23799], Fresh[23798], Fresh[23797], Fresh[23796], Fresh[23795], Fresh[23794], Fresh[23793], Fresh[23792], Fresh[23791], Fresh[23790], Fresh[23789], Fresh[23788], Fresh[23787], Fresh[23786], Fresh[23785], Fresh[23784], Fresh[23783], Fresh[23782], Fresh[23781], Fresh[23780], Fresh[23779], Fresh[23778], Fresh[23777], Fresh[23776], Fresh[23775], Fresh[23774], Fresh[23773], Fresh[23772], Fresh[23771], Fresh[23770], Fresh[23769], Fresh[23768], Fresh[23767], Fresh[23766], Fresh[23765], Fresh[23764], Fresh[23763], Fresh[23762], Fresh[23761], Fresh[23760], Fresh[23759], Fresh[23758], Fresh[23757], Fresh[23756], Fresh[23755], Fresh[23754], Fresh[23753], Fresh[23752], Fresh[23751], Fresh[23750], Fresh[23749], Fresh[23748], Fresh[23747], Fresh[23746], Fresh[23745], Fresh[23744], Fresh[23743], Fresh[23742], Fresh[23741], Fresh[23740], Fresh[23739], Fresh[23738], Fresh[23737], Fresh[23736], Fresh[23735], Fresh[23734], Fresh[23733], Fresh[23732], Fresh[23731], Fresh[23730], Fresh[23729], Fresh[23728], Fresh[23727], Fresh[23726], Fresh[23725], Fresh[23724], Fresh[23723], Fresh[23722], Fresh[23721], Fresh[23720], Fresh[23719], Fresh[23718], Fresh[23717], Fresh[23716], Fresh[23715], Fresh[23714], Fresh[23713], Fresh[23712], Fresh[23711], Fresh[23710], Fresh[23709], Fresh[23708], Fresh[23707], Fresh[23706], Fresh[23705], Fresh[23704], Fresh[23703], Fresh[23702], Fresh[23701], Fresh[23700], Fresh[23699], Fresh[23698], Fresh[23697], Fresh[23696], Fresh[23695], Fresh[23694], Fresh[23693], Fresh[23692], Fresh[23691], Fresh[23690], Fresh[23689], Fresh[23688], Fresh[23687], Fresh[23686], Fresh[23685], Fresh[23684], Fresh[23683], Fresh[23682], Fresh[23681], Fresh[23680], Fresh[23679], Fresh[23678], Fresh[23677], Fresh[23676], Fresh[23675], Fresh[23674], Fresh[23673], Fresh[23672], Fresh[23671], Fresh[23670], Fresh[23669], Fresh[23668], Fresh[23667], Fresh[23666], Fresh[23665], Fresh[23664], Fresh[23663], Fresh[23662], Fresh[23661], Fresh[23660], Fresh[23659], Fresh[23658], Fresh[23657], Fresh[23656], Fresh[23655], Fresh[23654], Fresh[23653], Fresh[23652], Fresh[23651], Fresh[23650], Fresh[23649], Fresh[23648], Fresh[23647], Fresh[23646], Fresh[23645], Fresh[23644], Fresh[23643], Fresh[23642], Fresh[23641], Fresh[23640], Fresh[23639], Fresh[23638], Fresh[23637], Fresh[23636], Fresh[23635], Fresh[23634], Fresh[23633], Fresh[23632], Fresh[23631], Fresh[23630], Fresh[23629], Fresh[23628], Fresh[23627], Fresh[23626], Fresh[23625], Fresh[23624], Fresh[23623], Fresh[23622], Fresh[23621], Fresh[23620], Fresh[23619], Fresh[23618], Fresh[23617], Fresh[23616], Fresh[23615], Fresh[23614], Fresh[23613], Fresh[23612], Fresh[23611], Fresh[23610], Fresh[23609], Fresh[23608], Fresh[23607], Fresh[23606], Fresh[23605], Fresh[23604], Fresh[23603], Fresh[23602], Fresh[23601], Fresh[23600], Fresh[23599], Fresh[23598], Fresh[23597], Fresh[23596], Fresh[23595], Fresh[23594], Fresh[23593], Fresh[23592], Fresh[23591], Fresh[23590], Fresh[23589], Fresh[23588], Fresh[23587], Fresh[23586], Fresh[23585], Fresh[23584], Fresh[23583], Fresh[23582], Fresh[23581], Fresh[23580], Fresh[23579], Fresh[23578], Fresh[23577], Fresh[23576], Fresh[23575], Fresh[23574], Fresh[23573], Fresh[23572], Fresh[23571], Fresh[23570], Fresh[23569], Fresh[23568], Fresh[23567], Fresh[23566], Fresh[23565], Fresh[23564], Fresh[23563], Fresh[23562], Fresh[23561], Fresh[23560], Fresh[23559], Fresh[23558], Fresh[23557], Fresh[23556], Fresh[23555], Fresh[23554], Fresh[23553], Fresh[23552], Fresh[23551], Fresh[23550], Fresh[23549], Fresh[23548], Fresh[23547], Fresh[23546], Fresh[23545], Fresh[23544], Fresh[23543], Fresh[23542], Fresh[23541], Fresh[23540], Fresh[23539], Fresh[23538], Fresh[23537], Fresh[23536], Fresh[23535], Fresh[23534], Fresh[23533], Fresh[23532], Fresh[23531], Fresh[23530], Fresh[23529], Fresh[23528], Fresh[23527], Fresh[23526], Fresh[23525], Fresh[23524], Fresh[23523], Fresh[23522], Fresh[23521], Fresh[23520], Fresh[23519], Fresh[23518], Fresh[23517], Fresh[23516], Fresh[23515], Fresh[23514], Fresh[23513], Fresh[23512], Fresh[23511], Fresh[23510], Fresh[23509], Fresh[23508], Fresh[23507], Fresh[23506], Fresh[23505], Fresh[23504], Fresh[23503], Fresh[23502], Fresh[23501], Fresh[23500], Fresh[23499], Fresh[23498], Fresh[23497], Fresh[23496], Fresh[23495], Fresh[23494], Fresh[23493], Fresh[23492], Fresh[23491], Fresh[23490], Fresh[23489], Fresh[23488], Fresh[23487], Fresh[23486], Fresh[23485], Fresh[23484], Fresh[23483], Fresh[23482], Fresh[23481], Fresh[23480], Fresh[23479], Fresh[23478], Fresh[23477], Fresh[23476], Fresh[23475], Fresh[23474], Fresh[23473], Fresh[23472], Fresh[23471], Fresh[23470], Fresh[23469], Fresh[23468], Fresh[23467], Fresh[23466], Fresh[23465], Fresh[23464], Fresh[23463], Fresh[23462], Fresh[23461], Fresh[23460], Fresh[23459], Fresh[23458], Fresh[23457], Fresh[23456], Fresh[23455], Fresh[23454], Fresh[23453], Fresh[23452], Fresh[23451], Fresh[23450], Fresh[23449], Fresh[23448], Fresh[23447], Fresh[23446], Fresh[23445], Fresh[23444], Fresh[23443], Fresh[23442], Fresh[23441], Fresh[23440], Fresh[23439], Fresh[23438], Fresh[23437], Fresh[23436], Fresh[23435], Fresh[23434], Fresh[23433], Fresh[23432], Fresh[23431], Fresh[23430], Fresh[23429], Fresh[23428], Fresh[23427], Fresh[23426], Fresh[23425], Fresh[23424], Fresh[23423], Fresh[23422], Fresh[23421], Fresh[23420], Fresh[23419], Fresh[23418], Fresh[23417], Fresh[23416], Fresh[23415], Fresh[23414], Fresh[23413], Fresh[23412], Fresh[23411], Fresh[23410], Fresh[23409], Fresh[23408], Fresh[23407], Fresh[23406], Fresh[23405], Fresh[23404], Fresh[23403], Fresh[23402], Fresh[23401], Fresh[23400], Fresh[23399], Fresh[23398], Fresh[23397], Fresh[23396], Fresh[23395], Fresh[23394], Fresh[23393], Fresh[23392], Fresh[23391], Fresh[23390], Fresh[23389], Fresh[23388], Fresh[23387], Fresh[23386], Fresh[23385], Fresh[23384], Fresh[23383], Fresh[23382], Fresh[23381], Fresh[23380], Fresh[23379], Fresh[23378], Fresh[23377], Fresh[23376], Fresh[23375], Fresh[23374], Fresh[23373], Fresh[23372], Fresh[23371], Fresh[23370], Fresh[23369], Fresh[23368], Fresh[23367], Fresh[23366], Fresh[23365], Fresh[23364], Fresh[23363], Fresh[23362], Fresh[23361], Fresh[23360], Fresh[23359], Fresh[23358], Fresh[23357], Fresh[23356], Fresh[23355], Fresh[23354], Fresh[23353], Fresh[23352], Fresh[23351], Fresh[23350], Fresh[23349], Fresh[23348], Fresh[23347], Fresh[23346], Fresh[23345], Fresh[23344], Fresh[23343], Fresh[23342], Fresh[23341], Fresh[23340], Fresh[23339], Fresh[23338], Fresh[23337], Fresh[23336], Fresh[23335], Fresh[23334], Fresh[23333], Fresh[23332], Fresh[23331], Fresh[23330], Fresh[23329], Fresh[23328], Fresh[23327], Fresh[23326], Fresh[23325], Fresh[23324], Fresh[23323], Fresh[23322], Fresh[23321], Fresh[23320], Fresh[23319], Fresh[23318], Fresh[23317], Fresh[23316], Fresh[23315], Fresh[23314], Fresh[23313], Fresh[23312], Fresh[23311], Fresh[23310], Fresh[23309], Fresh[23308], Fresh[23307], Fresh[23306], Fresh[23305], Fresh[23304], Fresh[23303], Fresh[23302], Fresh[23301], Fresh[23300], Fresh[23299], Fresh[23298], Fresh[23297], Fresh[23296], Fresh[23295], Fresh[23294], Fresh[23293], Fresh[23292], Fresh[23291], Fresh[23290], Fresh[23289], Fresh[23288], Fresh[23287], Fresh[23286], Fresh[23285], Fresh[23284], Fresh[23283], Fresh[23282], Fresh[23281], Fresh[23280], Fresh[23279], Fresh[23278], Fresh[23277], Fresh[23276], Fresh[23275], Fresh[23274], Fresh[23273], Fresh[23272], Fresh[23271], Fresh[23270], Fresh[23269], Fresh[23268], Fresh[23267], Fresh[23266], Fresh[23265], Fresh[23264], Fresh[23263], Fresh[23262], Fresh[23261], Fresh[23260], Fresh[23259], Fresh[23258], Fresh[23257], Fresh[23256], Fresh[23255], Fresh[23254], Fresh[23253], Fresh[23252], Fresh[23251], Fresh[23250], Fresh[23249], Fresh[23248], Fresh[23247], Fresh[23246], Fresh[23245], Fresh[23244], Fresh[23243], Fresh[23242], Fresh[23241], Fresh[23240], Fresh[23239], Fresh[23238], Fresh[23237], Fresh[23236], Fresh[23235], Fresh[23234], Fresh[23233], Fresh[23232], Fresh[23231], Fresh[23230], Fresh[23229], Fresh[23228], Fresh[23227], Fresh[23226], Fresh[23225], Fresh[23224], Fresh[23223], Fresh[23222], Fresh[23221], Fresh[23220], Fresh[23219], Fresh[23218], Fresh[23217], Fresh[23216], Fresh[23215], Fresh[23214], Fresh[23213], Fresh[23212], Fresh[23211], Fresh[23210], Fresh[23209], Fresh[23208], Fresh[23207], Fresh[23206], Fresh[23205], Fresh[23204], Fresh[23203], Fresh[23202], Fresh[23201], Fresh[23200], Fresh[23199], Fresh[23198], Fresh[23197], Fresh[23196], Fresh[23195], Fresh[23194], Fresh[23193], Fresh[23192], Fresh[23191], Fresh[23190], Fresh[23189], Fresh[23188], Fresh[23187], Fresh[23186], Fresh[23185], Fresh[23184], Fresh[23183], Fresh[23182], Fresh[23181], Fresh[23180], Fresh[23179], Fresh[23178], Fresh[23177], Fresh[23176], Fresh[23175], Fresh[23174], Fresh[23173], Fresh[23172], Fresh[23171], Fresh[23170], Fresh[23169], Fresh[23168], Fresh[23167], Fresh[23166], Fresh[23165], Fresh[23164], Fresh[23163], Fresh[23162], Fresh[23161], Fresh[23160], Fresh[23159], Fresh[23158], Fresh[23157], Fresh[23156], Fresh[23155], Fresh[23154], Fresh[23153], Fresh[23152], Fresh[23151], Fresh[23150], Fresh[23149], Fresh[23148], Fresh[23147], Fresh[23146], Fresh[23145], Fresh[23144], Fresh[23143], Fresh[23142], Fresh[23141], Fresh[23140], Fresh[23139], Fresh[23138], Fresh[23137], Fresh[23136], Fresh[23135], Fresh[23134], Fresh[23133], Fresh[23132], Fresh[23131], Fresh[23130], Fresh[23129], Fresh[23128], Fresh[23127], Fresh[23126], Fresh[23125], Fresh[23124], Fresh[23123], Fresh[23122], Fresh[23121], Fresh[23120], Fresh[23119], Fresh[23118], Fresh[23117], Fresh[23116], Fresh[23115], Fresh[23114], Fresh[23113], Fresh[23112], Fresh[23111], Fresh[23110], Fresh[23109], Fresh[23108], Fresh[23107], Fresh[23106], Fresh[23105], Fresh[23104], Fresh[23103], Fresh[23102], Fresh[23101], Fresh[23100], Fresh[23099], Fresh[23098], Fresh[23097], Fresh[23096], Fresh[23095], Fresh[23094], Fresh[23093], Fresh[23092], Fresh[23091], Fresh[23090], Fresh[23089], Fresh[23088], Fresh[23087], Fresh[23086], Fresh[23085], Fresh[23084], Fresh[23083], Fresh[23082], Fresh[23081], Fresh[23080], Fresh[23079], Fresh[23078], Fresh[23077], Fresh[23076], Fresh[23075], Fresh[23074], Fresh[23073], Fresh[23072], Fresh[23071], Fresh[23070], Fresh[23069], Fresh[23068], Fresh[23067], Fresh[23066], Fresh[23065], Fresh[23064], Fresh[23063], Fresh[23062], Fresh[23061], Fresh[23060], Fresh[23059], Fresh[23058], Fresh[23057], Fresh[23056], Fresh[23055], Fresh[23054], Fresh[23053], Fresh[23052], Fresh[23051], Fresh[23050], Fresh[23049], Fresh[23048], Fresh[23047], Fresh[23046], Fresh[23045], Fresh[23044], Fresh[23043], Fresh[23042], Fresh[23041], Fresh[23040], Fresh[23039], Fresh[23038], Fresh[23037], Fresh[23036], Fresh[23035], Fresh[23034], Fresh[23033], Fresh[23032], Fresh[23031], Fresh[23030], Fresh[23029], Fresh[23028], Fresh[23027], Fresh[23026], Fresh[23025], Fresh[23024], Fresh[23023], Fresh[23022], Fresh[23021], Fresh[23020], Fresh[23019], Fresh[23018], Fresh[23017], Fresh[23016], Fresh[23015], Fresh[23014], Fresh[23013], Fresh[23012], Fresh[23011], Fresh[23010], Fresh[23009], Fresh[23008], Fresh[23007], Fresh[23006], Fresh[23005], Fresh[23004], Fresh[23003], Fresh[23002], Fresh[23001], Fresh[23000], Fresh[22999], Fresh[22998], Fresh[22997], Fresh[22996], Fresh[22995], Fresh[22994], Fresh[22993], Fresh[22992], Fresh[22991], Fresh[22990], Fresh[22989], Fresh[22988], Fresh[22987], Fresh[22986], Fresh[22985], Fresh[22984], Fresh[22983], Fresh[22982], Fresh[22981], Fresh[22980], Fresh[22979], Fresh[22978], Fresh[22977], Fresh[22976], Fresh[22975], Fresh[22974], Fresh[22973], Fresh[22972], Fresh[22971], Fresh[22970], Fresh[22969], Fresh[22968], Fresh[22967], Fresh[22966], Fresh[22965], Fresh[22964], Fresh[22963], Fresh[22962], Fresh[22961], Fresh[22960], Fresh[22959], Fresh[22958], Fresh[22957], Fresh[22956], Fresh[22955], Fresh[22954], Fresh[22953], Fresh[22952], Fresh[22951], Fresh[22950], Fresh[22949], Fresh[22948], Fresh[22947], Fresh[22946], Fresh[22945], Fresh[22944], Fresh[22943], Fresh[22942], Fresh[22941], Fresh[22940], Fresh[22939], Fresh[22938], Fresh[22937], Fresh[22936], Fresh[22935], Fresh[22934], Fresh[22933], Fresh[22932], Fresh[22931], Fresh[22930], Fresh[22929], Fresh[22928], Fresh[22927], Fresh[22926], Fresh[22925], Fresh[22924], Fresh[22923], Fresh[22922], Fresh[22921], Fresh[22920], Fresh[22919], Fresh[22918], Fresh[22917], Fresh[22916], Fresh[22915], Fresh[22914], Fresh[22913], Fresh[22912], Fresh[22911], Fresh[22910], Fresh[22909], Fresh[22908], Fresh[22907], Fresh[22906], Fresh[22905], Fresh[22904], Fresh[22903], Fresh[22902], Fresh[22901], Fresh[22900], Fresh[22899], Fresh[22898], Fresh[22897], Fresh[22896], Fresh[22895], Fresh[22894], Fresh[22893], Fresh[22892], Fresh[22891], Fresh[22890], Fresh[22889], Fresh[22888], Fresh[22887], Fresh[22886], Fresh[22885], Fresh[22884], Fresh[22883], Fresh[22882], Fresh[22881], Fresh[22880], Fresh[22879], Fresh[22878], Fresh[22877], Fresh[22876], Fresh[22875], Fresh[22874], Fresh[22873], Fresh[22872], Fresh[22871], Fresh[22870], Fresh[22869], Fresh[22868], Fresh[22867], Fresh[22866], Fresh[22865], Fresh[22864], Fresh[22863], Fresh[22862], Fresh[22861], Fresh[22860], Fresh[22859], Fresh[22858], Fresh[22857], Fresh[22856], Fresh[22855], Fresh[22854], Fresh[22853], Fresh[22852], Fresh[22851], Fresh[22850], Fresh[22849], Fresh[22848], Fresh[22847], Fresh[22846], Fresh[22845], Fresh[22844], Fresh[22843], Fresh[22842], Fresh[22841], Fresh[22840], Fresh[22839], Fresh[22838], Fresh[22837], Fresh[22836], Fresh[22835], Fresh[22834], Fresh[22833], Fresh[22832], Fresh[22831], Fresh[22830], Fresh[22829], Fresh[22828], Fresh[22827], Fresh[22826], Fresh[22825], Fresh[22824], Fresh[22823], Fresh[22822], Fresh[22821], Fresh[22820], Fresh[22819], Fresh[22818], Fresh[22817], Fresh[22816], Fresh[22815], Fresh[22814], Fresh[22813], Fresh[22812], Fresh[22811], Fresh[22810], Fresh[22809], Fresh[22808], Fresh[22807], Fresh[22806], Fresh[22805], Fresh[22804], Fresh[22803], Fresh[22802], Fresh[22801], Fresh[22800], Fresh[22799], Fresh[22798], Fresh[22797], Fresh[22796], Fresh[22795], Fresh[22794], Fresh[22793], Fresh[22792], Fresh[22791], Fresh[22790], Fresh[22789], Fresh[22788], Fresh[22787], Fresh[22786], Fresh[22785], Fresh[22784], Fresh[22783], Fresh[22782], Fresh[22781], Fresh[22780], Fresh[22779], Fresh[22778], Fresh[22777], Fresh[22776], Fresh[22775], Fresh[22774], Fresh[22773], Fresh[22772], Fresh[22771], Fresh[22770], Fresh[22769], Fresh[22768], Fresh[22767], Fresh[22766], Fresh[22765], Fresh[22764], Fresh[22763], Fresh[22762], Fresh[22761], Fresh[22760], Fresh[22759], Fresh[22758], Fresh[22757], Fresh[22756], Fresh[22755], Fresh[22754], Fresh[22753], Fresh[22752], Fresh[22751], Fresh[22750], Fresh[22749], Fresh[22748], Fresh[22747], Fresh[22746], Fresh[22745], Fresh[22744], Fresh[22743], Fresh[22742], Fresh[22741], Fresh[22740], Fresh[22739], Fresh[22738], Fresh[22737], Fresh[22736], Fresh[22735], Fresh[22734], Fresh[22733], Fresh[22732], Fresh[22731], Fresh[22730], Fresh[22729], Fresh[22728], Fresh[22727], Fresh[22726], Fresh[22725], Fresh[22724], Fresh[22723], Fresh[22722], Fresh[22721], Fresh[22720], Fresh[22719], Fresh[22718], Fresh[22717], Fresh[22716], Fresh[22715], Fresh[22714], Fresh[22713], Fresh[22712], Fresh[22711], Fresh[22710], Fresh[22709], Fresh[22708], Fresh[22707], Fresh[22706], Fresh[22705], Fresh[22704], Fresh[22703], Fresh[22702], Fresh[22701], Fresh[22700], Fresh[22699], Fresh[22698], Fresh[22697], Fresh[22696], Fresh[22695], Fresh[22694], Fresh[22693], Fresh[22692], Fresh[22691], Fresh[22690], Fresh[22689], Fresh[22688], Fresh[22687], Fresh[22686], Fresh[22685], Fresh[22684], Fresh[22683], Fresh[22682], Fresh[22681], Fresh[22680], Fresh[22679], Fresh[22678], Fresh[22677], Fresh[22676], Fresh[22675], Fresh[22674], Fresh[22673], Fresh[22672], Fresh[22671], Fresh[22670], Fresh[22669], Fresh[22668], Fresh[22667], Fresh[22666], Fresh[22665], Fresh[22664], Fresh[22663], Fresh[22662], Fresh[22661], Fresh[22660], Fresh[22659], Fresh[22658], Fresh[22657], Fresh[22656], Fresh[22655], Fresh[22654], Fresh[22653], Fresh[22652], Fresh[22651], Fresh[22650], Fresh[22649], Fresh[22648], Fresh[22647], Fresh[22646], Fresh[22645], Fresh[22644], Fresh[22643], Fresh[22642], Fresh[22641], Fresh[22640], Fresh[22639], Fresh[22638], Fresh[22637], Fresh[22636], Fresh[22635], Fresh[22634], Fresh[22633], Fresh[22632], Fresh[22631], Fresh[22630], Fresh[22629], Fresh[22628], Fresh[22627], Fresh[22626], Fresh[22625], Fresh[22624], Fresh[22623], Fresh[22622], Fresh[22621], Fresh[22620], Fresh[22619], Fresh[22618], Fresh[22617], Fresh[22616], Fresh[22615], Fresh[22614], Fresh[22613], Fresh[22612], Fresh[22611], Fresh[22610], Fresh[22609], Fresh[22608], Fresh[22607], Fresh[22606], Fresh[22605], Fresh[22604], Fresh[22603], Fresh[22602], Fresh[22601], Fresh[22600], Fresh[22599], Fresh[22598], Fresh[22597], Fresh[22596], Fresh[22595], Fresh[22594], Fresh[22593], Fresh[22592], Fresh[22591], Fresh[22590], Fresh[22589], Fresh[22588], Fresh[22587], Fresh[22586], Fresh[22585], Fresh[22584], Fresh[22583], Fresh[22582], Fresh[22581], Fresh[22580], Fresh[22579], Fresh[22578], Fresh[22577], Fresh[22576], Fresh[22575], Fresh[22574], Fresh[22573], Fresh[22572], Fresh[22571], Fresh[22570], Fresh[22569], Fresh[22568], Fresh[22567], Fresh[22566], Fresh[22565], Fresh[22564], Fresh[22563], Fresh[22562], Fresh[22561], Fresh[22560], Fresh[22559], Fresh[22558], Fresh[22557], Fresh[22556], Fresh[22555], Fresh[22554], Fresh[22553], Fresh[22552], Fresh[22551], Fresh[22550], Fresh[22549], Fresh[22548], Fresh[22547], Fresh[22546], Fresh[22545], Fresh[22544], Fresh[22543], Fresh[22542], Fresh[22541], Fresh[22540], Fresh[22539], Fresh[22538], Fresh[22537], Fresh[22536], Fresh[22535], Fresh[22534], Fresh[22533], Fresh[22532], Fresh[22531], Fresh[22530], Fresh[22529], Fresh[22528], Fresh[22527], Fresh[22526], Fresh[22525], Fresh[22524], Fresh[22523], Fresh[22522], Fresh[22521], Fresh[22520], Fresh[22519], Fresh[22518], Fresh[22517], Fresh[22516], Fresh[22515], Fresh[22514], Fresh[22513], Fresh[22512], Fresh[22511], Fresh[22510], Fresh[22509], Fresh[22508], Fresh[22507], Fresh[22506], Fresh[22505], Fresh[22504], Fresh[22503], Fresh[22502], Fresh[22501], Fresh[22500], Fresh[22499], Fresh[22498], Fresh[22497], Fresh[22496], Fresh[22495], Fresh[22494], Fresh[22493], Fresh[22492], Fresh[22491], Fresh[22490], Fresh[22489], Fresh[22488], Fresh[22487], Fresh[22486], Fresh[22485], Fresh[22484], Fresh[22483], Fresh[22482], Fresh[22481], Fresh[22480], Fresh[22479], Fresh[22478], Fresh[22477], Fresh[22476], Fresh[22475], Fresh[22474], Fresh[22473], Fresh[22472], Fresh[22471], Fresh[22470], Fresh[22469], Fresh[22468], Fresh[22467], Fresh[22466], Fresh[22465], Fresh[22464], Fresh[22463], Fresh[22462], Fresh[22461], Fresh[22460], Fresh[22459], Fresh[22458], Fresh[22457], Fresh[22456], Fresh[22455], Fresh[22454], Fresh[22453], Fresh[22452], Fresh[22451], Fresh[22450], Fresh[22449], Fresh[22448], Fresh[22447], Fresh[22446], Fresh[22445], Fresh[22444], Fresh[22443], Fresh[22442], Fresh[22441], Fresh[22440], Fresh[22439], Fresh[22438], Fresh[22437], Fresh[22436], Fresh[22435], Fresh[22434], Fresh[22433], Fresh[22432], Fresh[22431], Fresh[22430], Fresh[22429], Fresh[22428], Fresh[22427], Fresh[22426], Fresh[22425], Fresh[22424], Fresh[22423], Fresh[22422], Fresh[22421], Fresh[22420], Fresh[22419], Fresh[22418], Fresh[22417], Fresh[22416], Fresh[22415], Fresh[22414], Fresh[22413], Fresh[22412], Fresh[22411], Fresh[22410], Fresh[22409], Fresh[22408], Fresh[22407], Fresh[22406], Fresh[22405], Fresh[22404], Fresh[22403], Fresh[22402], Fresh[22401], Fresh[22400], Fresh[22399], Fresh[22398], Fresh[22397], Fresh[22396], Fresh[22395], Fresh[22394], Fresh[22393], Fresh[22392], Fresh[22391], Fresh[22390], Fresh[22389], Fresh[22388], Fresh[22387], Fresh[22386], Fresh[22385], Fresh[22384], Fresh[22383], Fresh[22382], Fresh[22381], Fresh[22380], Fresh[22379], Fresh[22378], Fresh[22377], Fresh[22376], Fresh[22375], Fresh[22374], Fresh[22373], Fresh[22372], Fresh[22371], Fresh[22370], Fresh[22369], Fresh[22368], Fresh[22367], Fresh[22366], Fresh[22365], Fresh[22364], Fresh[22363], Fresh[22362], Fresh[22361], Fresh[22360], Fresh[22359], Fresh[22358], Fresh[22357], Fresh[22356], Fresh[22355], Fresh[22354], Fresh[22353], Fresh[22352], Fresh[22351], Fresh[22350], Fresh[22349], Fresh[22348], Fresh[22347], Fresh[22346], Fresh[22345], Fresh[22344], Fresh[22343], Fresh[22342], Fresh[22341], Fresh[22340], Fresh[22339], Fresh[22338], Fresh[22337], Fresh[22336], Fresh[22335], Fresh[22334], Fresh[22333], Fresh[22332], Fresh[22331], Fresh[22330], Fresh[22329], Fresh[22328], Fresh[22327], Fresh[22326], Fresh[22325], Fresh[22324], Fresh[22323], Fresh[22322], Fresh[22321], Fresh[22320], Fresh[22319], Fresh[22318], Fresh[22317], Fresh[22316], Fresh[22315], Fresh[22314], Fresh[22313], Fresh[22312], Fresh[22311], Fresh[22310], Fresh[22309], Fresh[22308], Fresh[22307], Fresh[22306], Fresh[22305], Fresh[22304], Fresh[22303], Fresh[22302], Fresh[22301], Fresh[22300], Fresh[22299], Fresh[22298], Fresh[22297], Fresh[22296], Fresh[22295], Fresh[22294], Fresh[22293], Fresh[22292], Fresh[22291], Fresh[22290], Fresh[22289], Fresh[22288], Fresh[22287], Fresh[22286], Fresh[22285], Fresh[22284], Fresh[22283], Fresh[22282], Fresh[22281], Fresh[22280], Fresh[22279], Fresh[22278], Fresh[22277], Fresh[22276], Fresh[22275], Fresh[22274], Fresh[22273], Fresh[22272], Fresh[22271], Fresh[22270], Fresh[22269], Fresh[22268], Fresh[22267], Fresh[22266], Fresh[22265], Fresh[22264], Fresh[22263], Fresh[22262], Fresh[22261], Fresh[22260], Fresh[22259], Fresh[22258], Fresh[22257], Fresh[22256], Fresh[22255], Fresh[22254], Fresh[22253], Fresh[22252], Fresh[22251], Fresh[22250], Fresh[22249], Fresh[22248], Fresh[22247], Fresh[22246], Fresh[22245], Fresh[22244], Fresh[22243], Fresh[22242], Fresh[22241], Fresh[22240], Fresh[22239], Fresh[22238], Fresh[22237], Fresh[22236], Fresh[22235], Fresh[22234], Fresh[22233], Fresh[22232], Fresh[22231], Fresh[22230], Fresh[22229], Fresh[22228], Fresh[22227], Fresh[22226], Fresh[22225], Fresh[22224], Fresh[22223], Fresh[22222], Fresh[22221], Fresh[22220], Fresh[22219], Fresh[22218], Fresh[22217], Fresh[22216], Fresh[22215], Fresh[22214], Fresh[22213], Fresh[22212], Fresh[22211], Fresh[22210], Fresh[22209], Fresh[22208], Fresh[22207], Fresh[22206], Fresh[22205], Fresh[22204], Fresh[22203], Fresh[22202], Fresh[22201], Fresh[22200], Fresh[22199], Fresh[22198], Fresh[22197], Fresh[22196], Fresh[22195], Fresh[22194], Fresh[22193], Fresh[22192], Fresh[22191], Fresh[22190], Fresh[22189], Fresh[22188], Fresh[22187], Fresh[22186], Fresh[22185], Fresh[22184], Fresh[22183], Fresh[22182], Fresh[22181], Fresh[22180], Fresh[22179], Fresh[22178], Fresh[22177], Fresh[22176], Fresh[22175], Fresh[22174], Fresh[22173], Fresh[22172], Fresh[22171], Fresh[22170], Fresh[22169], Fresh[22168], Fresh[22167], Fresh[22166], Fresh[22165], Fresh[22164], Fresh[22163], Fresh[22162], Fresh[22161], Fresh[22160], Fresh[22159], Fresh[22158], Fresh[22157], Fresh[22156], Fresh[22155], Fresh[22154], Fresh[22153], Fresh[22152], Fresh[22151], Fresh[22150], Fresh[22149], Fresh[22148], Fresh[22147], Fresh[22146], Fresh[22145], Fresh[22144], Fresh[22143], Fresh[22142], Fresh[22141], Fresh[22140], Fresh[22139], Fresh[22138], Fresh[22137], Fresh[22136], Fresh[22135], Fresh[22134], Fresh[22133], Fresh[22132], Fresh[22131], Fresh[22130], Fresh[22129], Fresh[22128], Fresh[22127], Fresh[22126], Fresh[22125], Fresh[22124], Fresh[22123], Fresh[22122], Fresh[22121], Fresh[22120], Fresh[22119], Fresh[22118], Fresh[22117], Fresh[22116], Fresh[22115], Fresh[22114], Fresh[22113], Fresh[22112], Fresh[22111], Fresh[22110], Fresh[22109], Fresh[22108], Fresh[22107], Fresh[22106], Fresh[22105], Fresh[22104], Fresh[22103], Fresh[22102], Fresh[22101], Fresh[22100], Fresh[22099], Fresh[22098], Fresh[22097], Fresh[22096], Fresh[22095], Fresh[22094], Fresh[22093], Fresh[22092], Fresh[22091], Fresh[22090], Fresh[22089], Fresh[22088], Fresh[22087], Fresh[22086], Fresh[22085], Fresh[22084], Fresh[22083], Fresh[22082], Fresh[22081], Fresh[22080], Fresh[22079], Fresh[22078], Fresh[22077], Fresh[22076], Fresh[22075], Fresh[22074], Fresh[22073], Fresh[22072], Fresh[22071], Fresh[22070], Fresh[22069], Fresh[22068], Fresh[22067], Fresh[22066], Fresh[22065], Fresh[22064], Fresh[22063], Fresh[22062], Fresh[22061], Fresh[22060], Fresh[22059], Fresh[22058], Fresh[22057], Fresh[22056], Fresh[22055], Fresh[22054], Fresh[22053], Fresh[22052], Fresh[22051], Fresh[22050], Fresh[22049], Fresh[22048], Fresh[22047], Fresh[22046], Fresh[22045], Fresh[22044], Fresh[22043], Fresh[22042], Fresh[22041], Fresh[22040], Fresh[22039], Fresh[22038], Fresh[22037], Fresh[22036], Fresh[22035], Fresh[22034], Fresh[22033], Fresh[22032], Fresh[22031], Fresh[22030], Fresh[22029], Fresh[22028], Fresh[22027], Fresh[22026], Fresh[22025], Fresh[22024], Fresh[22023], Fresh[22022], Fresh[22021], Fresh[22020], Fresh[22019], Fresh[22018], Fresh[22017], Fresh[22016], Fresh[22015], Fresh[22014], Fresh[22013], Fresh[22012], Fresh[22011], Fresh[22010], Fresh[22009], Fresh[22008], Fresh[22007], Fresh[22006], Fresh[22005], Fresh[22004], Fresh[22003], Fresh[22002], Fresh[22001], Fresh[22000], Fresh[21999], Fresh[21998], Fresh[21997], Fresh[21996], Fresh[21995], Fresh[21994], Fresh[21993], Fresh[21992], Fresh[21991], Fresh[21990], Fresh[21989], Fresh[21988], Fresh[21987], Fresh[21986], Fresh[21985], Fresh[21984], Fresh[21983], Fresh[21982], Fresh[21981], Fresh[21980], Fresh[21979], Fresh[21978], Fresh[21977], Fresh[21976], Fresh[21975], Fresh[21974], Fresh[21973], Fresh[21972], Fresh[21971], Fresh[21970], Fresh[21969], Fresh[21968], Fresh[21967], Fresh[21966], Fresh[21965], Fresh[21964], Fresh[21963], Fresh[21962], Fresh[21961], Fresh[21960], Fresh[21959], Fresh[21958], Fresh[21957], Fresh[21956], Fresh[21955], Fresh[21954], Fresh[21953], Fresh[21952], Fresh[21951], Fresh[21950], Fresh[21949], Fresh[21948], Fresh[21947], Fresh[21946], Fresh[21945], Fresh[21944], Fresh[21943], Fresh[21942], Fresh[21941], Fresh[21940], Fresh[21939], Fresh[21938], Fresh[21937], Fresh[21936], Fresh[21935], Fresh[21934], Fresh[21933], Fresh[21932], Fresh[21931], Fresh[21930], Fresh[21929], Fresh[21928], Fresh[21927], Fresh[21926], Fresh[21925], Fresh[21924], Fresh[21923], Fresh[21922], Fresh[21921], Fresh[21920], Fresh[21919], Fresh[21918], Fresh[21917], Fresh[21916], Fresh[21915], Fresh[21914], Fresh[21913], Fresh[21912], Fresh[21911], Fresh[21910], Fresh[21909], Fresh[21908], Fresh[21907], Fresh[21906], Fresh[21905], Fresh[21904], Fresh[21903], Fresh[21902], Fresh[21901], Fresh[21900], Fresh[21899], Fresh[21898], Fresh[21897], Fresh[21896], Fresh[21895], Fresh[21894], Fresh[21893], Fresh[21892], Fresh[21891], Fresh[21890], Fresh[21889], Fresh[21888], Fresh[21887], Fresh[21886], Fresh[21885], Fresh[21884], Fresh[21883], Fresh[21882], Fresh[21881], Fresh[21880], Fresh[21879], Fresh[21878], Fresh[21877], Fresh[21876], Fresh[21875], Fresh[21874], Fresh[21873], Fresh[21872], Fresh[21871], Fresh[21870], Fresh[21869], Fresh[21868], Fresh[21867], Fresh[21866], Fresh[21865], Fresh[21864], Fresh[21863], Fresh[21862], Fresh[21861], Fresh[21860], Fresh[21859], Fresh[21858], Fresh[21857], Fresh[21856], Fresh[21855], Fresh[21854], Fresh[21853], Fresh[21852], Fresh[21851], Fresh[21850], Fresh[21849], Fresh[21848], Fresh[21847], Fresh[21846], Fresh[21845], Fresh[21844], Fresh[21843], Fresh[21842], Fresh[21841], Fresh[21840], Fresh[21839], Fresh[21838], Fresh[21837], Fresh[21836], Fresh[21835], Fresh[21834], Fresh[21833], Fresh[21832], Fresh[21831], Fresh[21830], Fresh[21829], Fresh[21828], Fresh[21827], Fresh[21826], Fresh[21825], Fresh[21824], Fresh[21823], Fresh[21822], Fresh[21821], Fresh[21820], Fresh[21819], Fresh[21818], Fresh[21817], Fresh[21816], Fresh[21815], Fresh[21814], Fresh[21813], Fresh[21812], Fresh[21811], Fresh[21810], Fresh[21809], Fresh[21808], Fresh[21807], Fresh[21806], Fresh[21805], Fresh[21804], Fresh[21803], Fresh[21802], Fresh[21801], Fresh[21800], Fresh[21799], Fresh[21798], Fresh[21797], Fresh[21796], Fresh[21795], Fresh[21794], Fresh[21793], Fresh[21792], Fresh[21791], Fresh[21790], Fresh[21789], Fresh[21788], Fresh[21787], Fresh[21786], Fresh[21785], Fresh[21784], Fresh[21783], Fresh[21782], Fresh[21781], Fresh[21780], Fresh[21779], Fresh[21778], Fresh[21777], Fresh[21776], Fresh[21775], Fresh[21774], Fresh[21773], Fresh[21772], Fresh[21771], Fresh[21770], Fresh[21769], Fresh[21768], Fresh[21767], Fresh[21766], Fresh[21765], Fresh[21764], Fresh[21763], Fresh[21762], Fresh[21761], Fresh[21760], Fresh[21759], Fresh[21758], Fresh[21757], Fresh[21756], Fresh[21755], Fresh[21754], Fresh[21753], Fresh[21752], Fresh[21751], Fresh[21750], Fresh[21749], Fresh[21748], Fresh[21747], Fresh[21746], Fresh[21745], Fresh[21744], Fresh[21743], Fresh[21742], Fresh[21741], Fresh[21740], Fresh[21739], Fresh[21738], Fresh[21737], Fresh[21736], Fresh[21735], Fresh[21734], Fresh[21733], Fresh[21732], Fresh[21731], Fresh[21730], Fresh[21729], Fresh[21728], Fresh[21727], Fresh[21726], Fresh[21725], Fresh[21724], Fresh[21723], Fresh[21722], Fresh[21721], Fresh[21720], Fresh[21719], Fresh[21718], Fresh[21717], Fresh[21716], Fresh[21715], Fresh[21714], Fresh[21713], Fresh[21712], Fresh[21711], Fresh[21710], Fresh[21709], Fresh[21708], Fresh[21707], Fresh[21706], Fresh[21705], Fresh[21704], Fresh[21703], Fresh[21702], Fresh[21701], Fresh[21700], Fresh[21699], Fresh[21698], Fresh[21697], Fresh[21696], Fresh[21695], Fresh[21694], Fresh[21693], Fresh[21692], Fresh[21691], Fresh[21690], Fresh[21689], Fresh[21688], Fresh[21687], Fresh[21686], Fresh[21685], Fresh[21684], Fresh[21683], Fresh[21682], Fresh[21681], Fresh[21680], Fresh[21679], Fresh[21678], Fresh[21677], Fresh[21676], Fresh[21675], Fresh[21674], Fresh[21673], Fresh[21672], Fresh[21671], Fresh[21670], Fresh[21669], Fresh[21668], Fresh[21667], Fresh[21666], Fresh[21665], Fresh[21664], Fresh[21663], Fresh[21662], Fresh[21661], Fresh[21660], Fresh[21659], Fresh[21658], Fresh[21657], Fresh[21656], Fresh[21655], Fresh[21654], Fresh[21653], Fresh[21652], Fresh[21651], Fresh[21650], Fresh[21649], Fresh[21648], Fresh[21647], Fresh[21646], Fresh[21645], Fresh[21644], Fresh[21643], Fresh[21642], Fresh[21641], Fresh[21640], Fresh[21639], Fresh[21638], Fresh[21637], Fresh[21636], Fresh[21635], Fresh[21634], Fresh[21633], Fresh[21632], Fresh[21631], Fresh[21630], Fresh[21629], Fresh[21628], Fresh[21627], Fresh[21626], Fresh[21625], Fresh[21624], Fresh[21623], Fresh[21622], Fresh[21621], Fresh[21620], Fresh[21619], Fresh[21618], Fresh[21617], Fresh[21616], Fresh[21615], Fresh[21614], Fresh[21613], Fresh[21612], Fresh[21611], Fresh[21610], Fresh[21609], Fresh[21608], Fresh[21607], Fresh[21606], Fresh[21605], Fresh[21604], Fresh[21603], Fresh[21602], Fresh[21601], Fresh[21600], Fresh[21599], Fresh[21598], Fresh[21597], Fresh[21596], Fresh[21595], Fresh[21594], Fresh[21593], Fresh[21592], Fresh[21591], Fresh[21590], Fresh[21589], Fresh[21588], Fresh[21587], Fresh[21586], Fresh[21585], Fresh[21584], Fresh[21583], Fresh[21582], Fresh[21581], Fresh[21580], Fresh[21579], Fresh[21578], Fresh[21577], Fresh[21576], Fresh[21575], Fresh[21574], Fresh[21573], Fresh[21572], Fresh[21571], Fresh[21570], Fresh[21569], Fresh[21568], Fresh[21567], Fresh[21566], Fresh[21565], Fresh[21564], Fresh[21563], Fresh[21562], Fresh[21561], Fresh[21560], Fresh[21559], Fresh[21558], Fresh[21557], Fresh[21556], Fresh[21555], Fresh[21554], Fresh[21553], Fresh[21552], Fresh[21551], Fresh[21550], Fresh[21549], Fresh[21548], Fresh[21547], Fresh[21546], Fresh[21545], Fresh[21544], Fresh[21543], Fresh[21542], Fresh[21541], Fresh[21540], Fresh[21539], Fresh[21538], Fresh[21537], Fresh[21536], Fresh[21535], Fresh[21534], Fresh[21533], Fresh[21532], Fresh[21531], Fresh[21530], Fresh[21529], Fresh[21528], Fresh[21527], Fresh[21526], Fresh[21525], Fresh[21524], Fresh[21523], Fresh[21522], Fresh[21521], Fresh[21520], Fresh[21519], Fresh[21518], Fresh[21517], Fresh[21516], Fresh[21515], Fresh[21514], Fresh[21513], Fresh[21512], Fresh[21511], Fresh[21510], Fresh[21509], Fresh[21508], Fresh[21507], Fresh[21506], Fresh[21505], Fresh[21504], Fresh[21503], Fresh[21502], Fresh[21501], Fresh[21500], Fresh[21499], Fresh[21498], Fresh[21497], Fresh[21496], Fresh[21495], Fresh[21494], Fresh[21493], Fresh[21492], Fresh[21491], Fresh[21490], Fresh[21489], Fresh[21488], Fresh[21487], Fresh[21486], Fresh[21485], Fresh[21484], Fresh[21483], Fresh[21482], Fresh[21481], Fresh[21480], Fresh[21479], Fresh[21478], Fresh[21477], Fresh[21476], Fresh[21475], Fresh[21474], Fresh[21473], Fresh[21472], Fresh[21471], Fresh[21470], Fresh[21469], Fresh[21468], Fresh[21467], Fresh[21466], Fresh[21465], Fresh[21464], Fresh[21463], Fresh[21462], Fresh[21461], Fresh[21460], Fresh[21459], Fresh[21458], Fresh[21457], Fresh[21456], Fresh[21455], Fresh[21454], Fresh[21453], Fresh[21452], Fresh[21451], Fresh[21450], Fresh[21449], Fresh[21448], Fresh[21447], Fresh[21446], Fresh[21445], Fresh[21444], Fresh[21443], Fresh[21442], Fresh[21441], Fresh[21440], Fresh[21439], Fresh[21438], Fresh[21437], Fresh[21436], Fresh[21435], Fresh[21434], Fresh[21433], Fresh[21432], Fresh[21431], Fresh[21430], Fresh[21429], Fresh[21428], Fresh[21427], Fresh[21426], Fresh[21425], Fresh[21424], Fresh[21423], Fresh[21422], Fresh[21421], Fresh[21420], Fresh[21419], Fresh[21418], Fresh[21417], Fresh[21416], Fresh[21415], Fresh[21414], Fresh[21413], Fresh[21412], Fresh[21411], Fresh[21410], Fresh[21409], Fresh[21408], Fresh[21407], Fresh[21406], Fresh[21405], Fresh[21404], Fresh[21403], Fresh[21402], Fresh[21401], Fresh[21400], Fresh[21399], Fresh[21398], Fresh[21397], Fresh[21396], Fresh[21395], Fresh[21394], Fresh[21393], Fresh[21392], Fresh[21391], Fresh[21390], Fresh[21389], Fresh[21388], Fresh[21387], Fresh[21386], Fresh[21385], Fresh[21384], Fresh[21383], Fresh[21382], Fresh[21381], Fresh[21380], Fresh[21379], Fresh[21378], Fresh[21377], Fresh[21376], Fresh[21375], Fresh[21374], Fresh[21373], Fresh[21372], Fresh[21371], Fresh[21370], Fresh[21369], Fresh[21368], Fresh[21367], Fresh[21366], Fresh[21365], Fresh[21364], Fresh[21363], Fresh[21362], Fresh[21361], Fresh[21360], Fresh[21359], Fresh[21358], Fresh[21357], Fresh[21356], Fresh[21355], Fresh[21354], Fresh[21353], Fresh[21352], Fresh[21351], Fresh[21350], Fresh[21349], Fresh[21348], Fresh[21347], Fresh[21346], Fresh[21345], Fresh[21344], Fresh[21343], Fresh[21342], Fresh[21341], Fresh[21340], Fresh[21339], Fresh[21338], Fresh[21337], Fresh[21336], Fresh[21335], Fresh[21334], Fresh[21333], Fresh[21332], Fresh[21331], Fresh[21330], Fresh[21329], Fresh[21328], Fresh[21327], Fresh[21326], Fresh[21325], Fresh[21324], Fresh[21323], Fresh[21322], Fresh[21321], Fresh[21320], Fresh[21319], Fresh[21318], Fresh[21317], Fresh[21316], Fresh[21315], Fresh[21314], Fresh[21313], Fresh[21312], Fresh[21311], Fresh[21310], Fresh[21309], Fresh[21308], Fresh[21307], Fresh[21306], Fresh[21305], Fresh[21304], Fresh[21303], Fresh[21302], Fresh[21301], Fresh[21300], Fresh[21299], Fresh[21298], Fresh[21297], Fresh[21296], Fresh[21295], Fresh[21294], Fresh[21293], Fresh[21292], Fresh[21291], Fresh[21290], Fresh[21289], Fresh[21288], Fresh[21287], Fresh[21286], Fresh[21285], Fresh[21284], Fresh[21283], Fresh[21282], Fresh[21281], Fresh[21280], Fresh[21279], Fresh[21278], Fresh[21277], Fresh[21276], Fresh[21275], Fresh[21274], Fresh[21273], Fresh[21272], Fresh[21271], Fresh[21270], Fresh[21269], Fresh[21268], Fresh[21267], Fresh[21266], Fresh[21265], Fresh[21264], Fresh[21263], Fresh[21262], Fresh[21261], Fresh[21260], Fresh[21259], Fresh[21258], Fresh[21257], Fresh[21256], Fresh[21255], Fresh[21254], Fresh[21253], Fresh[21252], Fresh[21251], Fresh[21250], Fresh[21249], Fresh[21248], Fresh[21247], Fresh[21246], Fresh[21245], Fresh[21244], Fresh[21243], Fresh[21242], Fresh[21241], Fresh[21240], Fresh[21239], Fresh[21238], Fresh[21237], Fresh[21236], Fresh[21235], Fresh[21234], Fresh[21233], Fresh[21232], Fresh[21231], Fresh[21230], Fresh[21229], Fresh[21228], Fresh[21227], Fresh[21226], Fresh[21225], Fresh[21224], Fresh[21223], Fresh[21222], Fresh[21221], Fresh[21220], Fresh[21219], Fresh[21218], Fresh[21217], Fresh[21216], Fresh[21215], Fresh[21214], Fresh[21213], Fresh[21212], Fresh[21211], Fresh[21210], Fresh[21209], Fresh[21208], Fresh[21207], Fresh[21206], Fresh[21205], Fresh[21204], Fresh[21203], Fresh[21202], Fresh[21201], Fresh[21200], Fresh[21199], Fresh[21198], Fresh[21197], Fresh[21196], Fresh[21195], Fresh[21194], Fresh[21193], Fresh[21192], Fresh[21191], Fresh[21190], Fresh[21189], Fresh[21188], Fresh[21187], Fresh[21186], Fresh[21185], Fresh[21184], Fresh[21183], Fresh[21182], Fresh[21181], Fresh[21180], Fresh[21179], Fresh[21178], Fresh[21177], Fresh[21176], Fresh[21175], Fresh[21174], Fresh[21173], Fresh[21172], Fresh[21171], Fresh[21170], Fresh[21169], Fresh[21168], Fresh[21167], Fresh[21166], Fresh[21165], Fresh[21164], Fresh[21163], Fresh[21162], Fresh[21161], Fresh[21160], Fresh[21159], Fresh[21158], Fresh[21157], Fresh[21156], Fresh[21155], Fresh[21154], Fresh[21153], Fresh[21152], Fresh[21151], Fresh[21150], Fresh[21149], Fresh[21148], Fresh[21147], Fresh[21146], Fresh[21145], Fresh[21144], Fresh[21143], Fresh[21142], Fresh[21141], Fresh[21140], Fresh[21139], Fresh[21138], Fresh[21137], Fresh[21136], Fresh[21135], Fresh[21134], Fresh[21133], Fresh[21132], Fresh[21131], Fresh[21130], Fresh[21129], Fresh[21128], Fresh[21127], Fresh[21126], Fresh[21125], Fresh[21124], Fresh[21123], Fresh[21122], Fresh[21121], Fresh[21120], Fresh[21119], Fresh[21118], Fresh[21117], Fresh[21116], Fresh[21115], Fresh[21114], Fresh[21113], Fresh[21112], Fresh[21111], Fresh[21110], Fresh[21109], Fresh[21108], Fresh[21107], Fresh[21106], Fresh[21105], Fresh[21104], Fresh[21103], Fresh[21102], Fresh[21101], Fresh[21100], Fresh[21099], Fresh[21098], Fresh[21097], Fresh[21096], Fresh[21095], Fresh[21094], Fresh[21093], Fresh[21092], Fresh[21091], Fresh[21090], Fresh[21089], Fresh[21088], Fresh[21087], Fresh[21086], Fresh[21085], Fresh[21084], Fresh[21083], Fresh[21082], Fresh[21081], Fresh[21080], Fresh[21079], Fresh[21078], Fresh[21077], Fresh[21076], Fresh[21075], Fresh[21074], Fresh[21073], Fresh[21072], Fresh[21071], Fresh[21070], Fresh[21069], Fresh[21068], Fresh[21067], Fresh[21066], Fresh[21065], Fresh[21064], Fresh[21063], Fresh[21062], Fresh[21061], Fresh[21060], Fresh[21059], Fresh[21058], Fresh[21057], Fresh[21056], Fresh[21055], Fresh[21054], Fresh[21053], Fresh[21052], Fresh[21051], Fresh[21050], Fresh[21049], Fresh[21048], Fresh[21047], Fresh[21046], Fresh[21045], Fresh[21044], Fresh[21043], Fresh[21042], Fresh[21041], Fresh[21040], Fresh[21039], Fresh[21038], Fresh[21037], Fresh[21036], Fresh[21035], Fresh[21034], Fresh[21033], Fresh[21032], Fresh[21031], Fresh[21030], Fresh[21029], Fresh[21028], Fresh[21027], Fresh[21026], Fresh[21025], Fresh[21024], Fresh[21023], Fresh[21022], Fresh[21021], Fresh[21020], Fresh[21019], Fresh[21018], Fresh[21017], Fresh[21016], Fresh[21015], Fresh[21014], Fresh[21013], Fresh[21012], Fresh[21011], Fresh[21010], Fresh[21009], Fresh[21008], Fresh[21007], Fresh[21006], Fresh[21005], Fresh[21004], Fresh[21003], Fresh[21002], Fresh[21001], Fresh[21000], Fresh[20999], Fresh[20998], Fresh[20997], Fresh[20996], Fresh[20995], Fresh[20994], Fresh[20993], Fresh[20992], Fresh[20991], Fresh[20990], Fresh[20989], Fresh[20988], Fresh[20987], Fresh[20986], Fresh[20985], Fresh[20984], Fresh[20983], Fresh[20982], Fresh[20981], Fresh[20980], Fresh[20979], Fresh[20978], Fresh[20977], Fresh[20976], Fresh[20975], Fresh[20974], Fresh[20973], Fresh[20972], Fresh[20971], Fresh[20970], Fresh[20969], Fresh[20968], Fresh[20967], Fresh[20966], Fresh[20965], Fresh[20964], Fresh[20963], Fresh[20962], Fresh[20961], Fresh[20960], Fresh[20959], Fresh[20958], Fresh[20957], Fresh[20956], Fresh[20955], Fresh[20954], Fresh[20953], Fresh[20952], Fresh[20951], Fresh[20950], Fresh[20949], Fresh[20948], Fresh[20947], Fresh[20946], Fresh[20945], Fresh[20944], Fresh[20943], Fresh[20942], Fresh[20941], Fresh[20940], Fresh[20939], Fresh[20938], Fresh[20937], Fresh[20936], Fresh[20935], Fresh[20934], Fresh[20933], Fresh[20932], Fresh[20931], Fresh[20930], Fresh[20929], Fresh[20928], Fresh[20927], Fresh[20926], Fresh[20925], Fresh[20924], Fresh[20923], Fresh[20922], Fresh[20921], Fresh[20920], Fresh[20919], Fresh[20918], Fresh[20917], Fresh[20916], Fresh[20915], Fresh[20914], Fresh[20913], Fresh[20912], Fresh[20911], Fresh[20910], Fresh[20909], Fresh[20908], Fresh[20907], Fresh[20906], Fresh[20905], Fresh[20904], Fresh[20903], Fresh[20902], Fresh[20901], Fresh[20900], Fresh[20899], Fresh[20898], Fresh[20897], Fresh[20896], Fresh[20895], Fresh[20894], Fresh[20893], Fresh[20892], Fresh[20891], Fresh[20890], Fresh[20889], Fresh[20888], Fresh[20887], Fresh[20886], Fresh[20885], Fresh[20884], Fresh[20883], Fresh[20882], Fresh[20881], Fresh[20880], Fresh[20879], Fresh[20878], Fresh[20877], Fresh[20876], Fresh[20875], Fresh[20874], Fresh[20873], Fresh[20872], Fresh[20871], Fresh[20870], Fresh[20869], Fresh[20868], Fresh[20867], Fresh[20866], Fresh[20865], Fresh[20864], Fresh[20863], Fresh[20862], Fresh[20861], Fresh[20860], Fresh[20859], Fresh[20858], Fresh[20857], Fresh[20856], Fresh[20855], Fresh[20854], Fresh[20853], Fresh[20852], Fresh[20851], Fresh[20850], Fresh[20849], Fresh[20848], Fresh[20847], Fresh[20846], Fresh[20845], Fresh[20844], Fresh[20843], Fresh[20842], Fresh[20841], Fresh[20840], Fresh[20839], Fresh[20838], Fresh[20837], Fresh[20836], Fresh[20835], Fresh[20834], Fresh[20833], Fresh[20832], Fresh[20831], Fresh[20830], Fresh[20829], Fresh[20828], Fresh[20827], Fresh[20826], Fresh[20825], Fresh[20824], Fresh[20823], Fresh[20822], Fresh[20821], Fresh[20820], Fresh[20819], Fresh[20818], Fresh[20817], Fresh[20816], Fresh[20815], Fresh[20814], Fresh[20813], Fresh[20812], Fresh[20811], Fresh[20810], Fresh[20809], Fresh[20808], Fresh[20807], Fresh[20806], Fresh[20805], Fresh[20804], Fresh[20803], Fresh[20802], Fresh[20801], Fresh[20800], Fresh[20799], Fresh[20798], Fresh[20797], Fresh[20796], Fresh[20795], Fresh[20794], Fresh[20793], Fresh[20792], Fresh[20791], Fresh[20790], Fresh[20789], Fresh[20788], Fresh[20787], Fresh[20786], Fresh[20785], Fresh[20784], Fresh[20783], Fresh[20782], Fresh[20781], Fresh[20780], Fresh[20779], Fresh[20778], Fresh[20777], Fresh[20776], Fresh[20775], Fresh[20774], Fresh[20773], Fresh[20772], Fresh[20771], Fresh[20770], Fresh[20769], Fresh[20768], Fresh[20767], Fresh[20766], Fresh[20765], Fresh[20764], Fresh[20763], Fresh[20762], Fresh[20761], Fresh[20760], Fresh[20759], Fresh[20758], Fresh[20757], Fresh[20756], Fresh[20755], Fresh[20754], Fresh[20753], Fresh[20752], Fresh[20751], Fresh[20750], Fresh[20749], Fresh[20748], Fresh[20747], Fresh[20746], Fresh[20745], Fresh[20744], Fresh[20743], Fresh[20742], Fresh[20741], Fresh[20740], Fresh[20739], Fresh[20738], Fresh[20737], Fresh[20736], Fresh[20735], Fresh[20734], Fresh[20733], Fresh[20732], Fresh[20731], Fresh[20730], Fresh[20729], Fresh[20728], Fresh[20727], Fresh[20726], Fresh[20725], Fresh[20724], Fresh[20723], Fresh[20722], Fresh[20721], Fresh[20720], Fresh[20719], Fresh[20718], Fresh[20717], Fresh[20716], Fresh[20715], Fresh[20714], Fresh[20713], Fresh[20712], Fresh[20711], Fresh[20710], Fresh[20709], Fresh[20708], Fresh[20707], Fresh[20706], Fresh[20705], Fresh[20704], Fresh[20703], Fresh[20702], Fresh[20701], Fresh[20700], Fresh[20699], Fresh[20698], Fresh[20697], Fresh[20696], Fresh[20695], Fresh[20694], Fresh[20693], Fresh[20692], Fresh[20691], Fresh[20690], Fresh[20689], Fresh[20688], Fresh[20687], Fresh[20686], Fresh[20685], Fresh[20684], Fresh[20683], Fresh[20682], Fresh[20681], Fresh[20680], Fresh[20679], Fresh[20678], Fresh[20677], Fresh[20676], Fresh[20675], Fresh[20674], Fresh[20673], Fresh[20672], Fresh[20671], Fresh[20670], Fresh[20669], Fresh[20668], Fresh[20667], Fresh[20666], Fresh[20665], Fresh[20664], Fresh[20663], Fresh[20662], Fresh[20661], Fresh[20660], Fresh[20659], Fresh[20658], Fresh[20657], Fresh[20656], Fresh[20655], Fresh[20654], Fresh[20653], Fresh[20652], Fresh[20651], Fresh[20650], Fresh[20649], Fresh[20648], Fresh[20647], Fresh[20646], Fresh[20645], Fresh[20644], Fresh[20643], Fresh[20642], Fresh[20641], Fresh[20640], Fresh[20639], Fresh[20638], Fresh[20637], Fresh[20636], Fresh[20635], Fresh[20634], Fresh[20633], Fresh[20632], Fresh[20631], Fresh[20630], Fresh[20629], Fresh[20628], Fresh[20627], Fresh[20626], Fresh[20625], Fresh[20624], Fresh[20623], Fresh[20622], Fresh[20621], Fresh[20620], Fresh[20619], Fresh[20618], Fresh[20617], Fresh[20616], Fresh[20615], Fresh[20614], Fresh[20613], Fresh[20612], Fresh[20611], Fresh[20610], Fresh[20609], Fresh[20608], Fresh[20607], Fresh[20606], Fresh[20605], Fresh[20604], Fresh[20603], Fresh[20602], Fresh[20601], Fresh[20600], Fresh[20599], Fresh[20598], Fresh[20597], Fresh[20596], Fresh[20595], Fresh[20594], Fresh[20593], Fresh[20592], Fresh[20591], Fresh[20590], Fresh[20589], Fresh[20588], Fresh[20587], Fresh[20586], Fresh[20585], Fresh[20584], Fresh[20583], Fresh[20582], Fresh[20581], Fresh[20580], Fresh[20579], Fresh[20578], Fresh[20577], Fresh[20576], Fresh[20575], Fresh[20574], Fresh[20573], Fresh[20572], Fresh[20571], Fresh[20570], Fresh[20569], Fresh[20568], Fresh[20567], Fresh[20566], Fresh[20565], Fresh[20564], Fresh[20563], Fresh[20562], Fresh[20561], Fresh[20560], Fresh[20559], Fresh[20558], Fresh[20557], Fresh[20556], Fresh[20555], Fresh[20554], Fresh[20553], Fresh[20552], Fresh[20551], Fresh[20550], Fresh[20549], Fresh[20548], Fresh[20547], Fresh[20546], Fresh[20545], Fresh[20544], Fresh[20543], Fresh[20542], Fresh[20541], Fresh[20540], Fresh[20539], Fresh[20538], Fresh[20537], Fresh[20536], Fresh[20535], Fresh[20534], Fresh[20533], Fresh[20532], Fresh[20531], Fresh[20530], Fresh[20529], Fresh[20528], Fresh[20527], Fresh[20526], Fresh[20525], Fresh[20524], Fresh[20523], Fresh[20522], Fresh[20521], Fresh[20520], Fresh[20519], Fresh[20518], Fresh[20517], Fresh[20516], Fresh[20515], Fresh[20514], Fresh[20513], Fresh[20512], Fresh[20511], Fresh[20510], Fresh[20509], Fresh[20508], Fresh[20507], Fresh[20506], Fresh[20505], Fresh[20504], Fresh[20503], Fresh[20502], Fresh[20501], Fresh[20500], Fresh[20499], Fresh[20498], Fresh[20497], Fresh[20496], Fresh[20495], Fresh[20494], Fresh[20493], Fresh[20492], Fresh[20491], Fresh[20490], Fresh[20489], Fresh[20488], Fresh[20487], Fresh[20486], Fresh[20485], Fresh[20484], Fresh[20483], Fresh[20482], Fresh[20481], Fresh[20480], Fresh[20479], Fresh[20478], Fresh[20477], Fresh[20476], Fresh[20475], Fresh[20474], Fresh[20473], Fresh[20472], Fresh[20471], Fresh[20470], Fresh[20469], Fresh[20468], Fresh[20467], Fresh[20466], Fresh[20465], Fresh[20464], Fresh[20463], Fresh[20462], Fresh[20461], Fresh[20460], Fresh[20459], Fresh[20458], Fresh[20457], Fresh[20456], Fresh[20455], Fresh[20454], Fresh[20453], Fresh[20452], Fresh[20451], Fresh[20450], Fresh[20449], Fresh[20448], Fresh[20447], Fresh[20446], Fresh[20445], Fresh[20444], Fresh[20443], Fresh[20442], Fresh[20441], Fresh[20440], Fresh[20439], Fresh[20438], Fresh[20437], Fresh[20436], Fresh[20435], Fresh[20434], Fresh[20433], Fresh[20432], Fresh[20431], Fresh[20430], Fresh[20429], Fresh[20428], Fresh[20427], Fresh[20426], Fresh[20425], Fresh[20424], Fresh[20423], Fresh[20422], Fresh[20421], Fresh[20420], Fresh[20419], Fresh[20418], Fresh[20417], Fresh[20416], Fresh[20415], Fresh[20414], Fresh[20413], Fresh[20412], Fresh[20411], Fresh[20410], Fresh[20409], Fresh[20408], Fresh[20407], Fresh[20406], Fresh[20405], Fresh[20404], Fresh[20403], Fresh[20402], Fresh[20401], Fresh[20400], Fresh[20399], Fresh[20398], Fresh[20397], Fresh[20396], Fresh[20395], Fresh[20394], Fresh[20393], Fresh[20392], Fresh[20391], Fresh[20390], Fresh[20389], Fresh[20388], Fresh[20387], Fresh[20386], Fresh[20385], Fresh[20384], Fresh[20383], Fresh[20382], Fresh[20381], Fresh[20380], Fresh[20379], Fresh[20378], Fresh[20377], Fresh[20376], Fresh[20375], Fresh[20374], Fresh[20373], Fresh[20372], Fresh[20371], Fresh[20370], Fresh[20369], Fresh[20368], Fresh[20367], Fresh[20366], Fresh[20365], Fresh[20364], Fresh[20363], Fresh[20362], Fresh[20361], Fresh[20360], Fresh[20359], Fresh[20358], Fresh[20357], Fresh[20356], Fresh[20355], Fresh[20354], Fresh[20353], Fresh[20352], Fresh[20351], Fresh[20350], Fresh[20349], Fresh[20348], Fresh[20347], Fresh[20346], Fresh[20345], Fresh[20344], Fresh[20343], Fresh[20342], Fresh[20341], Fresh[20340], Fresh[20339], Fresh[20338], Fresh[20337], Fresh[20336], Fresh[20335], Fresh[20334], Fresh[20333], Fresh[20332], Fresh[20331], Fresh[20330], Fresh[20329], Fresh[20328], Fresh[20327], Fresh[20326], Fresh[20325], Fresh[20324], Fresh[20323], Fresh[20322], Fresh[20321], Fresh[20320], Fresh[20319], Fresh[20318], Fresh[20317], Fresh[20316], Fresh[20315], Fresh[20314], Fresh[20313], Fresh[20312], Fresh[20311], Fresh[20310], Fresh[20309], Fresh[20308], Fresh[20307], Fresh[20306], Fresh[20305], Fresh[20304], Fresh[20303], Fresh[20302], Fresh[20301], Fresh[20300], Fresh[20299], Fresh[20298], Fresh[20297], Fresh[20296], Fresh[20295], Fresh[20294], Fresh[20293], Fresh[20292], Fresh[20291], Fresh[20290], Fresh[20289], Fresh[20288], Fresh[20287], Fresh[20286], Fresh[20285], Fresh[20284], Fresh[20283], Fresh[20282], Fresh[20281], Fresh[20280], Fresh[20279], Fresh[20278], Fresh[20277], Fresh[20276], Fresh[20275], Fresh[20274], Fresh[20273], Fresh[20272], Fresh[20271], Fresh[20270], Fresh[20269], Fresh[20268], Fresh[20267], Fresh[20266], Fresh[20265], Fresh[20264], Fresh[20263], Fresh[20262], Fresh[20261], Fresh[20260], Fresh[20259], Fresh[20258], Fresh[20257], Fresh[20256], Fresh[20255], Fresh[20254], Fresh[20253], Fresh[20252], Fresh[20251], Fresh[20250], Fresh[20249], Fresh[20248], Fresh[20247], Fresh[20246], Fresh[20245], Fresh[20244], Fresh[20243], Fresh[20242], Fresh[20241], Fresh[20240], Fresh[20239], Fresh[20238], Fresh[20237], Fresh[20236], Fresh[20235], Fresh[20234], Fresh[20233], Fresh[20232], Fresh[20231], Fresh[20230], Fresh[20229], Fresh[20228], Fresh[20227], Fresh[20226], Fresh[20225], Fresh[20224], Fresh[20223], Fresh[20222], Fresh[20221], Fresh[20220], Fresh[20219], Fresh[20218], Fresh[20217], Fresh[20216], Fresh[20215], Fresh[20214], Fresh[20213], Fresh[20212], Fresh[20211], Fresh[20210], Fresh[20209], Fresh[20208], Fresh[20207], Fresh[20206], Fresh[20205], Fresh[20204], Fresh[20203], Fresh[20202], Fresh[20201], Fresh[20200], Fresh[20199], Fresh[20198], Fresh[20197], Fresh[20196], Fresh[20195], Fresh[20194], Fresh[20193], Fresh[20192], Fresh[20191], Fresh[20190], Fresh[20189], Fresh[20188], Fresh[20187], Fresh[20186], Fresh[20185], Fresh[20184], Fresh[20183], Fresh[20182], Fresh[20181], Fresh[20180], Fresh[20179], Fresh[20178], Fresh[20177], Fresh[20176], Fresh[20175], Fresh[20174], Fresh[20173], Fresh[20172], Fresh[20171], Fresh[20170], Fresh[20169], Fresh[20168], Fresh[20167], Fresh[20166], Fresh[20165], Fresh[20164], Fresh[20163], Fresh[20162], Fresh[20161], Fresh[20160], Fresh[20159], Fresh[20158], Fresh[20157], Fresh[20156], Fresh[20155], Fresh[20154], Fresh[20153], Fresh[20152], Fresh[20151], Fresh[20150], Fresh[20149], Fresh[20148], Fresh[20147], Fresh[20146], Fresh[20145], Fresh[20144], Fresh[20143], Fresh[20142], Fresh[20141], Fresh[20140], Fresh[20139], Fresh[20138], Fresh[20137], Fresh[20136], Fresh[20135], Fresh[20134], Fresh[20133], Fresh[20132], Fresh[20131], Fresh[20130], Fresh[20129], Fresh[20128], Fresh[20127], Fresh[20126], Fresh[20125], Fresh[20124], Fresh[20123], Fresh[20122], Fresh[20121], Fresh[20120], Fresh[20119], Fresh[20118], Fresh[20117], Fresh[20116], Fresh[20115], Fresh[20114], Fresh[20113], Fresh[20112], Fresh[20111], Fresh[20110], Fresh[20109], Fresh[20108], Fresh[20107], Fresh[20106], Fresh[20105], Fresh[20104], Fresh[20103], Fresh[20102], Fresh[20101], Fresh[20100], Fresh[20099], Fresh[20098], Fresh[20097], Fresh[20096], Fresh[20095], Fresh[20094], Fresh[20093], Fresh[20092], Fresh[20091], Fresh[20090], Fresh[20089], Fresh[20088], Fresh[20087], Fresh[20086], Fresh[20085], Fresh[20084], Fresh[20083], Fresh[20082], Fresh[20081], Fresh[20080], Fresh[20079], Fresh[20078], Fresh[20077], Fresh[20076], Fresh[20075], Fresh[20074], Fresh[20073], Fresh[20072], Fresh[20071], Fresh[20070], Fresh[20069], Fresh[20068], Fresh[20067], Fresh[20066], Fresh[20065], Fresh[20064], Fresh[20063], Fresh[20062], Fresh[20061], Fresh[20060], Fresh[20059], Fresh[20058], Fresh[20057], Fresh[20056], Fresh[20055], Fresh[20054], Fresh[20053], Fresh[20052], Fresh[20051], Fresh[20050], Fresh[20049], Fresh[20048], Fresh[20047], Fresh[20046], Fresh[20045], Fresh[20044], Fresh[20043], Fresh[20042], Fresh[20041], Fresh[20040], Fresh[20039], Fresh[20038], Fresh[20037], Fresh[20036], Fresh[20035], Fresh[20034], Fresh[20033], Fresh[20032], Fresh[20031], Fresh[20030], Fresh[20029], Fresh[20028], Fresh[20027], Fresh[20026], Fresh[20025], Fresh[20024], Fresh[20023], Fresh[20022], Fresh[20021], Fresh[20020], Fresh[20019], Fresh[20018], Fresh[20017], Fresh[20016], Fresh[20015], Fresh[20014], Fresh[20013], Fresh[20012], Fresh[20011], Fresh[20010], Fresh[20009], Fresh[20008], Fresh[20007], Fresh[20006], Fresh[20005], Fresh[20004], Fresh[20003], Fresh[20002], Fresh[20001], Fresh[20000], Fresh[19999], Fresh[19998], Fresh[19997], Fresh[19996], Fresh[19995], Fresh[19994], Fresh[19993], Fresh[19992], Fresh[19991], Fresh[19990], Fresh[19989], Fresh[19988], Fresh[19987], Fresh[19986], Fresh[19985], Fresh[19984], Fresh[19983], Fresh[19982], Fresh[19981], Fresh[19980], Fresh[19979], Fresh[19978], Fresh[19977], Fresh[19976], Fresh[19975], Fresh[19974], Fresh[19973], Fresh[19972], Fresh[19971], Fresh[19970], Fresh[19969], Fresh[19968], Fresh[19967], Fresh[19966], Fresh[19965], Fresh[19964], Fresh[19963], Fresh[19962], Fresh[19961], Fresh[19960], Fresh[19959], Fresh[19958], Fresh[19957], Fresh[19956], Fresh[19955], Fresh[19954], Fresh[19953], Fresh[19952], Fresh[19951], Fresh[19950], Fresh[19949], Fresh[19948], Fresh[19947], Fresh[19946], Fresh[19945], Fresh[19944], Fresh[19943], Fresh[19942], Fresh[19941], Fresh[19940], Fresh[19939], Fresh[19938], Fresh[19937], Fresh[19936], Fresh[19935], Fresh[19934], Fresh[19933], Fresh[19932], Fresh[19931], Fresh[19930], Fresh[19929], Fresh[19928], Fresh[19927], Fresh[19926], Fresh[19925], Fresh[19924], Fresh[19923], Fresh[19922], Fresh[19921], Fresh[19920], Fresh[19919], Fresh[19918], Fresh[19917], Fresh[19916], Fresh[19915], Fresh[19914], Fresh[19913], Fresh[19912], Fresh[19911], Fresh[19910], Fresh[19909], Fresh[19908], Fresh[19907], Fresh[19906], Fresh[19905], Fresh[19904], Fresh[19903], Fresh[19902], Fresh[19901], Fresh[19900], Fresh[19899], Fresh[19898], Fresh[19897], Fresh[19896], Fresh[19895], Fresh[19894], Fresh[19893], Fresh[19892], Fresh[19891], Fresh[19890], Fresh[19889], Fresh[19888], Fresh[19887], Fresh[19886], Fresh[19885], Fresh[19884], Fresh[19883], Fresh[19882], Fresh[19881], Fresh[19880], Fresh[19879], Fresh[19878], Fresh[19877], Fresh[19876], Fresh[19875], Fresh[19874], Fresh[19873], Fresh[19872], Fresh[19871], Fresh[19870], Fresh[19869], Fresh[19868], Fresh[19867], Fresh[19866], Fresh[19865], Fresh[19864], Fresh[19863], Fresh[19862], Fresh[19861], Fresh[19860], Fresh[19859], Fresh[19858], Fresh[19857], Fresh[19856], Fresh[19855], Fresh[19854], Fresh[19853], Fresh[19852], Fresh[19851], Fresh[19850], Fresh[19849], Fresh[19848], Fresh[19847], Fresh[19846], Fresh[19845], Fresh[19844], Fresh[19843], Fresh[19842], Fresh[19841], Fresh[19840], Fresh[19839], Fresh[19838], Fresh[19837], Fresh[19836], Fresh[19835], Fresh[19834], Fresh[19833], Fresh[19832], Fresh[19831], Fresh[19830], Fresh[19829], Fresh[19828], Fresh[19827], Fresh[19826], Fresh[19825], Fresh[19824], Fresh[19823], Fresh[19822], Fresh[19821], Fresh[19820], Fresh[19819], Fresh[19818], Fresh[19817], Fresh[19816], Fresh[19815], Fresh[19814], Fresh[19813], Fresh[19812], Fresh[19811], Fresh[19810], Fresh[19809], Fresh[19808], Fresh[19807], Fresh[19806], Fresh[19805], Fresh[19804], Fresh[19803], Fresh[19802], Fresh[19801], Fresh[19800], Fresh[19799], Fresh[19798], Fresh[19797], Fresh[19796], Fresh[19795], Fresh[19794], Fresh[19793], Fresh[19792], Fresh[19791], Fresh[19790], Fresh[19789], Fresh[19788], Fresh[19787], Fresh[19786], Fresh[19785], Fresh[19784], Fresh[19783], Fresh[19782], Fresh[19781], Fresh[19780], Fresh[19779], Fresh[19778], Fresh[19777], Fresh[19776], Fresh[19775], Fresh[19774], Fresh[19773], Fresh[19772], Fresh[19771], Fresh[19770], Fresh[19769], Fresh[19768], Fresh[19767], Fresh[19766], Fresh[19765], Fresh[19764], Fresh[19763], Fresh[19762], Fresh[19761], Fresh[19760], Fresh[19759], Fresh[19758], Fresh[19757], Fresh[19756], Fresh[19755], Fresh[19754], Fresh[19753], Fresh[19752], Fresh[19751], Fresh[19750], Fresh[19749], Fresh[19748], Fresh[19747], Fresh[19746], Fresh[19745], Fresh[19744], Fresh[19743], Fresh[19742], Fresh[19741], Fresh[19740], Fresh[19739], Fresh[19738], Fresh[19737], Fresh[19736], Fresh[19735], Fresh[19734], Fresh[19733], Fresh[19732], Fresh[19731], Fresh[19730], Fresh[19729], Fresh[19728], Fresh[19727], Fresh[19726], Fresh[19725], Fresh[19724], Fresh[19723], Fresh[19722], Fresh[19721], Fresh[19720], Fresh[19719], Fresh[19718], Fresh[19717], Fresh[19716], Fresh[19715], Fresh[19714], Fresh[19713], Fresh[19712], Fresh[19711], Fresh[19710], Fresh[19709], Fresh[19708], Fresh[19707], Fresh[19706], Fresh[19705], Fresh[19704], Fresh[19703], Fresh[19702], Fresh[19701], Fresh[19700], Fresh[19699], Fresh[19698], Fresh[19697], Fresh[19696], Fresh[19695], Fresh[19694], Fresh[19693], Fresh[19692], Fresh[19691], Fresh[19690], Fresh[19689], Fresh[19688], Fresh[19687], Fresh[19686], Fresh[19685], Fresh[19684], Fresh[19683], Fresh[19682], Fresh[19681], Fresh[19680], Fresh[19679], Fresh[19678], Fresh[19677], Fresh[19676], Fresh[19675], Fresh[19674], Fresh[19673], Fresh[19672], Fresh[19671], Fresh[19670], Fresh[19669], Fresh[19668], Fresh[19667], Fresh[19666], Fresh[19665], Fresh[19664], Fresh[19663], Fresh[19662], Fresh[19661], Fresh[19660], Fresh[19659], Fresh[19658], Fresh[19657], Fresh[19656], Fresh[19655], Fresh[19654], Fresh[19653], Fresh[19652], Fresh[19651], Fresh[19650], Fresh[19649], Fresh[19648], Fresh[19647], Fresh[19646], Fresh[19645], Fresh[19644], Fresh[19643], Fresh[19642], Fresh[19641], Fresh[19640], Fresh[19639], Fresh[19638], Fresh[19637], Fresh[19636], Fresh[19635], Fresh[19634], Fresh[19633], Fresh[19632], Fresh[19631], Fresh[19630], Fresh[19629], Fresh[19628], Fresh[19627], Fresh[19626], Fresh[19625], Fresh[19624], Fresh[19623], Fresh[19622], Fresh[19621], Fresh[19620], Fresh[19619], Fresh[19618], Fresh[19617], Fresh[19616], Fresh[19615], Fresh[19614], Fresh[19613], Fresh[19612], Fresh[19611], Fresh[19610], Fresh[19609], Fresh[19608], Fresh[19607], Fresh[19606], Fresh[19605], Fresh[19604], Fresh[19603], Fresh[19602], Fresh[19601], Fresh[19600], Fresh[19599], Fresh[19598], Fresh[19597], Fresh[19596], Fresh[19595], Fresh[19594], Fresh[19593], Fresh[19592], Fresh[19591], Fresh[19590], Fresh[19589], Fresh[19588], Fresh[19587], Fresh[19586], Fresh[19585], Fresh[19584], Fresh[19583], Fresh[19582], Fresh[19581], Fresh[19580], Fresh[19579], Fresh[19578], Fresh[19577], Fresh[19576], Fresh[19575], Fresh[19574], Fresh[19573], Fresh[19572], Fresh[19571], Fresh[19570], Fresh[19569], Fresh[19568], Fresh[19567], Fresh[19566], Fresh[19565], Fresh[19564], Fresh[19563], Fresh[19562], Fresh[19561], Fresh[19560], Fresh[19559], Fresh[19558], Fresh[19557], Fresh[19556], Fresh[19555], Fresh[19554], Fresh[19553], Fresh[19552], Fresh[19551], Fresh[19550], Fresh[19549], Fresh[19548], Fresh[19547], Fresh[19546], Fresh[19545], Fresh[19544], Fresh[19543], Fresh[19542], Fresh[19541], Fresh[19540], Fresh[19539], Fresh[19538], Fresh[19537], Fresh[19536], Fresh[19535], Fresh[19534], Fresh[19533], Fresh[19532], Fresh[19531], Fresh[19530], Fresh[19529], Fresh[19528], Fresh[19527], Fresh[19526], Fresh[19525], Fresh[19524], Fresh[19523], Fresh[19522], Fresh[19521], Fresh[19520], Fresh[19519], Fresh[19518], Fresh[19517], Fresh[19516], Fresh[19515], Fresh[19514], Fresh[19513], Fresh[19512], Fresh[19511], Fresh[19510], Fresh[19509], Fresh[19508], Fresh[19507], Fresh[19506], Fresh[19505], Fresh[19504], Fresh[19503], Fresh[19502], Fresh[19501], Fresh[19500], Fresh[19499], Fresh[19498], Fresh[19497], Fresh[19496], Fresh[19495], Fresh[19494], Fresh[19493], Fresh[19492], Fresh[19491], Fresh[19490], Fresh[19489], Fresh[19488], Fresh[19487], Fresh[19486], Fresh[19485], Fresh[19484], Fresh[19483], Fresh[19482], Fresh[19481], Fresh[19480], Fresh[19479], Fresh[19478], Fresh[19477], Fresh[19476], Fresh[19475], Fresh[19474], Fresh[19473], Fresh[19472], Fresh[19471], Fresh[19470], Fresh[19469], Fresh[19468], Fresh[19467], Fresh[19466], Fresh[19465], Fresh[19464], Fresh[19463], Fresh[19462], Fresh[19461], Fresh[19460], Fresh[19459], Fresh[19458], Fresh[19457], Fresh[19456], Fresh[19455], Fresh[19454], Fresh[19453], Fresh[19452], Fresh[19451], Fresh[19450], Fresh[19449], Fresh[19448], Fresh[19447], Fresh[19446], Fresh[19445], Fresh[19444], Fresh[19443], Fresh[19442], Fresh[19441], Fresh[19440], Fresh[19439], Fresh[19438], Fresh[19437], Fresh[19436], Fresh[19435], Fresh[19434], Fresh[19433], Fresh[19432], Fresh[19431], Fresh[19430], Fresh[19429], Fresh[19428], Fresh[19427], Fresh[19426], Fresh[19425], Fresh[19424], Fresh[19423], Fresh[19422], Fresh[19421], Fresh[19420], Fresh[19419], Fresh[19418], Fresh[19417], Fresh[19416], Fresh[19415], Fresh[19414], Fresh[19413], Fresh[19412], Fresh[19411], Fresh[19410], Fresh[19409], Fresh[19408], Fresh[19407], Fresh[19406], Fresh[19405], Fresh[19404], Fresh[19403], Fresh[19402], Fresh[19401], Fresh[19400], Fresh[19399], Fresh[19398], Fresh[19397], Fresh[19396], Fresh[19395], Fresh[19394], Fresh[19393], Fresh[19392], Fresh[19391], Fresh[19390], Fresh[19389], Fresh[19388], Fresh[19387], Fresh[19386], Fresh[19385], Fresh[19384], Fresh[19383], Fresh[19382], Fresh[19381], Fresh[19380], Fresh[19379], Fresh[19378], Fresh[19377], Fresh[19376], Fresh[19375], Fresh[19374], Fresh[19373], Fresh[19372], Fresh[19371], Fresh[19370], Fresh[19369], Fresh[19368], Fresh[19367], Fresh[19366], Fresh[19365], Fresh[19364], Fresh[19363], Fresh[19362], Fresh[19361], Fresh[19360], Fresh[19359], Fresh[19358], Fresh[19357], Fresh[19356], Fresh[19355], Fresh[19354], Fresh[19353], Fresh[19352], Fresh[19351], Fresh[19350], Fresh[19349], Fresh[19348], Fresh[19347], Fresh[19346], Fresh[19345], Fresh[19344], Fresh[19343], Fresh[19342], Fresh[19341], Fresh[19340], Fresh[19339], Fresh[19338], Fresh[19337], Fresh[19336], Fresh[19335], Fresh[19334], Fresh[19333], Fresh[19332], Fresh[19331], Fresh[19330], Fresh[19329], Fresh[19328], Fresh[19327], Fresh[19326], Fresh[19325], Fresh[19324], Fresh[19323], Fresh[19322], Fresh[19321], Fresh[19320], Fresh[19319], Fresh[19318], Fresh[19317], Fresh[19316], Fresh[19315], Fresh[19314], Fresh[19313], Fresh[19312], Fresh[19311], Fresh[19310], Fresh[19309], Fresh[19308], Fresh[19307], Fresh[19306], Fresh[19305], Fresh[19304], Fresh[19303], Fresh[19302], Fresh[19301], Fresh[19300], Fresh[19299], Fresh[19298], Fresh[19297], Fresh[19296], Fresh[19295], Fresh[19294], Fresh[19293], Fresh[19292], Fresh[19291], Fresh[19290], Fresh[19289], Fresh[19288], Fresh[19287], Fresh[19286], Fresh[19285], Fresh[19284], Fresh[19283], Fresh[19282], Fresh[19281], Fresh[19280], Fresh[19279], Fresh[19278], Fresh[19277], Fresh[19276], Fresh[19275], Fresh[19274], Fresh[19273], Fresh[19272], Fresh[19271], Fresh[19270], Fresh[19269], Fresh[19268], Fresh[19267], Fresh[19266], Fresh[19265], Fresh[19264], Fresh[19263], Fresh[19262], Fresh[19261], Fresh[19260], Fresh[19259], Fresh[19258], Fresh[19257], Fresh[19256], Fresh[19255], Fresh[19254], Fresh[19253], Fresh[19252], Fresh[19251], Fresh[19250], Fresh[19249], Fresh[19248], Fresh[19247], Fresh[19246], Fresh[19245], Fresh[19244], Fresh[19243], Fresh[19242], Fresh[19241], Fresh[19240], Fresh[19239], Fresh[19238], Fresh[19237], Fresh[19236], Fresh[19235], Fresh[19234], Fresh[19233], Fresh[19232], Fresh[19231], Fresh[19230], Fresh[19229], Fresh[19228], Fresh[19227], Fresh[19226], Fresh[19225], Fresh[19224], Fresh[19223], Fresh[19222], Fresh[19221], Fresh[19220], Fresh[19219], Fresh[19218], Fresh[19217], Fresh[19216], Fresh[19215], Fresh[19214], Fresh[19213], Fresh[19212], Fresh[19211], Fresh[19210], Fresh[19209], Fresh[19208], Fresh[19207], Fresh[19206], Fresh[19205], Fresh[19204], Fresh[19203], Fresh[19202], Fresh[19201], Fresh[19200], Fresh[19199], Fresh[19198], Fresh[19197], Fresh[19196], Fresh[19195], Fresh[19194], Fresh[19193], Fresh[19192], Fresh[19191], Fresh[19190], Fresh[19189], Fresh[19188], Fresh[19187], Fresh[19186], Fresh[19185], Fresh[19184], Fresh[19183], Fresh[19182], Fresh[19181], Fresh[19180], Fresh[19179], Fresh[19178], Fresh[19177], Fresh[19176], Fresh[19175], Fresh[19174], Fresh[19173], Fresh[19172], Fresh[19171], Fresh[19170], Fresh[19169], Fresh[19168], Fresh[19167], Fresh[19166], Fresh[19165], Fresh[19164], Fresh[19163], Fresh[19162], Fresh[19161], Fresh[19160], Fresh[19159], Fresh[19158], Fresh[19157], Fresh[19156], Fresh[19155], Fresh[19154], Fresh[19153], Fresh[19152], Fresh[19151], Fresh[19150], Fresh[19149], Fresh[19148], Fresh[19147], Fresh[19146], Fresh[19145], Fresh[19144], Fresh[19143], Fresh[19142], Fresh[19141], Fresh[19140], Fresh[19139], Fresh[19138], Fresh[19137], Fresh[19136], Fresh[19135], Fresh[19134], Fresh[19133], Fresh[19132], Fresh[19131], Fresh[19130], Fresh[19129], Fresh[19128], Fresh[19127], Fresh[19126], Fresh[19125], Fresh[19124], Fresh[19123], Fresh[19122], Fresh[19121], Fresh[19120], Fresh[19119], Fresh[19118], Fresh[19117], Fresh[19116], Fresh[19115], Fresh[19114], Fresh[19113], Fresh[19112], Fresh[19111], Fresh[19110], Fresh[19109], Fresh[19108], Fresh[19107], Fresh[19106], Fresh[19105], Fresh[19104], Fresh[19103], Fresh[19102], Fresh[19101], Fresh[19100], Fresh[19099], Fresh[19098], Fresh[19097], Fresh[19096], Fresh[19095], Fresh[19094], Fresh[19093], Fresh[19092], Fresh[19091], Fresh[19090], Fresh[19089], Fresh[19088], Fresh[19087], Fresh[19086], Fresh[19085], Fresh[19084], Fresh[19083], Fresh[19082], Fresh[19081], Fresh[19080], Fresh[19079], Fresh[19078], Fresh[19077], Fresh[19076], Fresh[19075], Fresh[19074], Fresh[19073], Fresh[19072], Fresh[19071], Fresh[19070], Fresh[19069], Fresh[19068], Fresh[19067], Fresh[19066], Fresh[19065], Fresh[19064], Fresh[19063], Fresh[19062], Fresh[19061], Fresh[19060], Fresh[19059], Fresh[19058], Fresh[19057], Fresh[19056], Fresh[19055], Fresh[19054], Fresh[19053], Fresh[19052], Fresh[19051], Fresh[19050], Fresh[19049], Fresh[19048], Fresh[19047], Fresh[19046], Fresh[19045], Fresh[19044], Fresh[19043], Fresh[19042], Fresh[19041], Fresh[19040], Fresh[19039], Fresh[19038], Fresh[19037], Fresh[19036], Fresh[19035], Fresh[19034], Fresh[19033], Fresh[19032], Fresh[19031], Fresh[19030], Fresh[19029], Fresh[19028], Fresh[19027], Fresh[19026], Fresh[19025], Fresh[19024], Fresh[19023], Fresh[19022], Fresh[19021], Fresh[19020], Fresh[19019], Fresh[19018], Fresh[19017], Fresh[19016], Fresh[19015], Fresh[19014], Fresh[19013], Fresh[19012], Fresh[19011], Fresh[19010], Fresh[19009], Fresh[19008], Fresh[19007], Fresh[19006], Fresh[19005], Fresh[19004], Fresh[19003], Fresh[19002], Fresh[19001], Fresh[19000], Fresh[18999], Fresh[18998], Fresh[18997], Fresh[18996], Fresh[18995], Fresh[18994], Fresh[18993], Fresh[18992], Fresh[18991], Fresh[18990], Fresh[18989], Fresh[18988], Fresh[18987], Fresh[18986], Fresh[18985], Fresh[18984], Fresh[18983], Fresh[18982], Fresh[18981], Fresh[18980], Fresh[18979], Fresh[18978], Fresh[18977], Fresh[18976], Fresh[18975], Fresh[18974], Fresh[18973], Fresh[18972], Fresh[18971], Fresh[18970], Fresh[18969], Fresh[18968], Fresh[18967], Fresh[18966], Fresh[18965], Fresh[18964], Fresh[18963], Fresh[18962], Fresh[18961], Fresh[18960], Fresh[18959], Fresh[18958], Fresh[18957], Fresh[18956], Fresh[18955], Fresh[18954], Fresh[18953], Fresh[18952], Fresh[18951], Fresh[18950], Fresh[18949], Fresh[18948], Fresh[18947], Fresh[18946], Fresh[18945], Fresh[18944], Fresh[18943], Fresh[18942], Fresh[18941], Fresh[18940], Fresh[18939], Fresh[18938], Fresh[18937], Fresh[18936], Fresh[18935], Fresh[18934], Fresh[18933], Fresh[18932], Fresh[18931], Fresh[18930], Fresh[18929], Fresh[18928], Fresh[18927], Fresh[18926], Fresh[18925], Fresh[18924], Fresh[18923], Fresh[18922], Fresh[18921], Fresh[18920], Fresh[18919], Fresh[18918], Fresh[18917], Fresh[18916], Fresh[18915], Fresh[18914], Fresh[18913], Fresh[18912], Fresh[18911], Fresh[18910], Fresh[18909], Fresh[18908], Fresh[18907], Fresh[18906], Fresh[18905], Fresh[18904], Fresh[18903], Fresh[18902], Fresh[18901], Fresh[18900], Fresh[18899], Fresh[18898], Fresh[18897], Fresh[18896], Fresh[18895], Fresh[18894], Fresh[18893], Fresh[18892], Fresh[18891], Fresh[18890], Fresh[18889], Fresh[18888], Fresh[18887], Fresh[18886], Fresh[18885], Fresh[18884], Fresh[18883], Fresh[18882], Fresh[18881], Fresh[18880], Fresh[18879], Fresh[18878], Fresh[18877], Fresh[18876], Fresh[18875], Fresh[18874], Fresh[18873], Fresh[18872], Fresh[18871], Fresh[18870], Fresh[18869], Fresh[18868], Fresh[18867], Fresh[18866], Fresh[18865], Fresh[18864], Fresh[18863], Fresh[18862], Fresh[18861], Fresh[18860], Fresh[18859], Fresh[18858], Fresh[18857], Fresh[18856], Fresh[18855], Fresh[18854], Fresh[18853], Fresh[18852], Fresh[18851], Fresh[18850], Fresh[18849], Fresh[18848], Fresh[18847], Fresh[18846], Fresh[18845], Fresh[18844], Fresh[18843], Fresh[18842], Fresh[18841], Fresh[18840], Fresh[18839], Fresh[18838], Fresh[18837], Fresh[18836], Fresh[18835], Fresh[18834], Fresh[18833], Fresh[18832], Fresh[18831], Fresh[18830], Fresh[18829], Fresh[18828], Fresh[18827], Fresh[18826], Fresh[18825], Fresh[18824], Fresh[18823], Fresh[18822], Fresh[18821], Fresh[18820], Fresh[18819], Fresh[18818], Fresh[18817], Fresh[18816], Fresh[18815], Fresh[18814], Fresh[18813], Fresh[18812], Fresh[18811], Fresh[18810], Fresh[18809], Fresh[18808], Fresh[18807], Fresh[18806], Fresh[18805], Fresh[18804], Fresh[18803], Fresh[18802], Fresh[18801], Fresh[18800], Fresh[18799], Fresh[18798], Fresh[18797], Fresh[18796], Fresh[18795], Fresh[18794], Fresh[18793], Fresh[18792], Fresh[18791], Fresh[18790], Fresh[18789], Fresh[18788], Fresh[18787], Fresh[18786], Fresh[18785], Fresh[18784], Fresh[18783], Fresh[18782], Fresh[18781], Fresh[18780], Fresh[18779], Fresh[18778], Fresh[18777], Fresh[18776], Fresh[18775], Fresh[18774], Fresh[18773], Fresh[18772], Fresh[18771], Fresh[18770], Fresh[18769], Fresh[18768], Fresh[18767], Fresh[18766], Fresh[18765], Fresh[18764], Fresh[18763], Fresh[18762], Fresh[18761], Fresh[18760], Fresh[18759], Fresh[18758], Fresh[18757], Fresh[18756], Fresh[18755], Fresh[18754], Fresh[18753], Fresh[18752], Fresh[18751], Fresh[18750], Fresh[18749], Fresh[18748], Fresh[18747], Fresh[18746], Fresh[18745], Fresh[18744], Fresh[18743], Fresh[18742], Fresh[18741], Fresh[18740], Fresh[18739], Fresh[18738], Fresh[18737], Fresh[18736], Fresh[18735], Fresh[18734], Fresh[18733], Fresh[18732], Fresh[18731], Fresh[18730], Fresh[18729], Fresh[18728], Fresh[18727], Fresh[18726], Fresh[18725], Fresh[18724], Fresh[18723], Fresh[18722], Fresh[18721], Fresh[18720], Fresh[18719], Fresh[18718], Fresh[18717], Fresh[18716], Fresh[18715], Fresh[18714], Fresh[18713], Fresh[18712], Fresh[18711], Fresh[18710], Fresh[18709], Fresh[18708], Fresh[18707], Fresh[18706], Fresh[18705], Fresh[18704], Fresh[18703], Fresh[18702], Fresh[18701], Fresh[18700], Fresh[18699], Fresh[18698], Fresh[18697], Fresh[18696], Fresh[18695], Fresh[18694], Fresh[18693], Fresh[18692], Fresh[18691], Fresh[18690], Fresh[18689], Fresh[18688], Fresh[18687], Fresh[18686], Fresh[18685], Fresh[18684], Fresh[18683], Fresh[18682], Fresh[18681], Fresh[18680], Fresh[18679], Fresh[18678], Fresh[18677], Fresh[18676], Fresh[18675], Fresh[18674], Fresh[18673], Fresh[18672], Fresh[18671], Fresh[18670], Fresh[18669], Fresh[18668], Fresh[18667], Fresh[18666], Fresh[18665], Fresh[18664], Fresh[18663], Fresh[18662], Fresh[18661], Fresh[18660], Fresh[18659], Fresh[18658], Fresh[18657], Fresh[18656], Fresh[18655], Fresh[18654], Fresh[18653], Fresh[18652], Fresh[18651], Fresh[18650], Fresh[18649], Fresh[18648], Fresh[18647], Fresh[18646], Fresh[18645], Fresh[18644], Fresh[18643], Fresh[18642], Fresh[18641], Fresh[18640], Fresh[18639], Fresh[18638], Fresh[18637], Fresh[18636], Fresh[18635], Fresh[18634], Fresh[18633], Fresh[18632], Fresh[18631], Fresh[18630], Fresh[18629], Fresh[18628], Fresh[18627], Fresh[18626], Fresh[18625], Fresh[18624], Fresh[18623], Fresh[18622], Fresh[18621], Fresh[18620], Fresh[18619], Fresh[18618], Fresh[18617], Fresh[18616], Fresh[18615], Fresh[18614], Fresh[18613], Fresh[18612], Fresh[18611], Fresh[18610], Fresh[18609], Fresh[18608], Fresh[18607], Fresh[18606], Fresh[18605], Fresh[18604], Fresh[18603], Fresh[18602], Fresh[18601], Fresh[18600], Fresh[18599], Fresh[18598], Fresh[18597], Fresh[18596], Fresh[18595], Fresh[18594], Fresh[18593], Fresh[18592], Fresh[18591], Fresh[18590], Fresh[18589], Fresh[18588], Fresh[18587], Fresh[18586], Fresh[18585], Fresh[18584], Fresh[18583], Fresh[18582], Fresh[18581], Fresh[18580], Fresh[18579], Fresh[18578], Fresh[18577], Fresh[18576], Fresh[18575], Fresh[18574], Fresh[18573], Fresh[18572], Fresh[18571], Fresh[18570], Fresh[18569], Fresh[18568], Fresh[18567], Fresh[18566], Fresh[18565], Fresh[18564], Fresh[18563], Fresh[18562], Fresh[18561], Fresh[18560], Fresh[18559], Fresh[18558], Fresh[18557], Fresh[18556], Fresh[18555], Fresh[18554], Fresh[18553], Fresh[18552], Fresh[18551], Fresh[18550], Fresh[18549], Fresh[18548], Fresh[18547], Fresh[18546], Fresh[18545], Fresh[18544], Fresh[18543], Fresh[18542], Fresh[18541], Fresh[18540], Fresh[18539], Fresh[18538], Fresh[18537], Fresh[18536], Fresh[18535], Fresh[18534], Fresh[18533], Fresh[18532], Fresh[18531], Fresh[18530], Fresh[18529], Fresh[18528], Fresh[18527], Fresh[18526], Fresh[18525], Fresh[18524], Fresh[18523], Fresh[18522], Fresh[18521], Fresh[18520], Fresh[18519], Fresh[18518], Fresh[18517], Fresh[18516], Fresh[18515], Fresh[18514], Fresh[18513], Fresh[18512], Fresh[18511], Fresh[18510], Fresh[18509], Fresh[18508], Fresh[18507], Fresh[18506], Fresh[18505], Fresh[18504], Fresh[18503], Fresh[18502], Fresh[18501], Fresh[18500], Fresh[18499], Fresh[18498], Fresh[18497], Fresh[18496], Fresh[18495], Fresh[18494], Fresh[18493], Fresh[18492], Fresh[18491], Fresh[18490], Fresh[18489], Fresh[18488], Fresh[18487], Fresh[18486], Fresh[18485], Fresh[18484], Fresh[18483], Fresh[18482], Fresh[18481], Fresh[18480], Fresh[18479], Fresh[18478], Fresh[18477], Fresh[18476], Fresh[18475], Fresh[18474], Fresh[18473], Fresh[18472], Fresh[18471], Fresh[18470], Fresh[18469], Fresh[18468], Fresh[18467], Fresh[18466], Fresh[18465], Fresh[18464], Fresh[18463], Fresh[18462], Fresh[18461], Fresh[18460], Fresh[18459], Fresh[18458], Fresh[18457], Fresh[18456], Fresh[18455], Fresh[18454], Fresh[18453], Fresh[18452], Fresh[18451], Fresh[18450], Fresh[18449], Fresh[18448], Fresh[18447], Fresh[18446], Fresh[18445], Fresh[18444], Fresh[18443], Fresh[18442], Fresh[18441], Fresh[18440], Fresh[18439], Fresh[18438], Fresh[18437], Fresh[18436], Fresh[18435], Fresh[18434], Fresh[18433], Fresh[18432], Fresh[18431], Fresh[18430], Fresh[18429], Fresh[18428], Fresh[18427], Fresh[18426], Fresh[18425], Fresh[18424], Fresh[18423], Fresh[18422], Fresh[18421], Fresh[18420], Fresh[18419], Fresh[18418], Fresh[18417], Fresh[18416], Fresh[18415], Fresh[18414], Fresh[18413], Fresh[18412], Fresh[18411], Fresh[18410], Fresh[18409], Fresh[18408], Fresh[18407], Fresh[18406], Fresh[18405], Fresh[18404], Fresh[18403], Fresh[18402], Fresh[18401], Fresh[18400], Fresh[18399], Fresh[18398], Fresh[18397], Fresh[18396], Fresh[18395], Fresh[18394], Fresh[18393], Fresh[18392], Fresh[18391], Fresh[18390], Fresh[18389], Fresh[18388], Fresh[18387], Fresh[18386], Fresh[18385], Fresh[18384], Fresh[18383], Fresh[18382], Fresh[18381], Fresh[18380], Fresh[18379], Fresh[18378], Fresh[18377], Fresh[18376], Fresh[18375], Fresh[18374], Fresh[18373], Fresh[18372], Fresh[18371], Fresh[18370], Fresh[18369], Fresh[18368], Fresh[18367], Fresh[18366], Fresh[18365], Fresh[18364], Fresh[18363], Fresh[18362], Fresh[18361], Fresh[18360], Fresh[18359], Fresh[18358], Fresh[18357], Fresh[18356], Fresh[18355], Fresh[18354], Fresh[18353], Fresh[18352], Fresh[18351], Fresh[18350], Fresh[18349], Fresh[18348], Fresh[18347], Fresh[18346], Fresh[18345], Fresh[18344], Fresh[18343], Fresh[18342], Fresh[18341], Fresh[18340], Fresh[18339], Fresh[18338], Fresh[18337], Fresh[18336], Fresh[18335], Fresh[18334], Fresh[18333], Fresh[18332], Fresh[18331], Fresh[18330], Fresh[18329], Fresh[18328], Fresh[18327], Fresh[18326], Fresh[18325], Fresh[18324], Fresh[18323], Fresh[18322], Fresh[18321], Fresh[18320], Fresh[18319], Fresh[18318], Fresh[18317], Fresh[18316], Fresh[18315], Fresh[18314], Fresh[18313], Fresh[18312], Fresh[18311], Fresh[18310], Fresh[18309], Fresh[18308], Fresh[18307], Fresh[18306], Fresh[18305], Fresh[18304], Fresh[18303], Fresh[18302], Fresh[18301], Fresh[18300], Fresh[18299], Fresh[18298], Fresh[18297], Fresh[18296], Fresh[18295], Fresh[18294], Fresh[18293], Fresh[18292], Fresh[18291], Fresh[18290], Fresh[18289], Fresh[18288], Fresh[18287], Fresh[18286], Fresh[18285], Fresh[18284], Fresh[18283], Fresh[18282], Fresh[18281], Fresh[18280], Fresh[18279], Fresh[18278], Fresh[18277], Fresh[18276], Fresh[18275], Fresh[18274], Fresh[18273], Fresh[18272], Fresh[18271], Fresh[18270], Fresh[18269], Fresh[18268], Fresh[18267], Fresh[18266], Fresh[18265], Fresh[18264], Fresh[18263], Fresh[18262], Fresh[18261], Fresh[18260], Fresh[18259], Fresh[18258], Fresh[18257], Fresh[18256], Fresh[18255], Fresh[18254], Fresh[18253], Fresh[18252], Fresh[18251], Fresh[18250], Fresh[18249], Fresh[18248], Fresh[18247], Fresh[18246], Fresh[18245], Fresh[18244], Fresh[18243], Fresh[18242], Fresh[18241], Fresh[18240], Fresh[18239], Fresh[18238], Fresh[18237], Fresh[18236], Fresh[18235], Fresh[18234], Fresh[18233], Fresh[18232], Fresh[18231], Fresh[18230], Fresh[18229], Fresh[18228], Fresh[18227], Fresh[18226], Fresh[18225], Fresh[18224], Fresh[18223], Fresh[18222], Fresh[18221], Fresh[18220], Fresh[18219], Fresh[18218], Fresh[18217], Fresh[18216], Fresh[18215], Fresh[18214], Fresh[18213], Fresh[18212], Fresh[18211], Fresh[18210], Fresh[18209], Fresh[18208], Fresh[18207], Fresh[18206], Fresh[18205], Fresh[18204], Fresh[18203], Fresh[18202], Fresh[18201], Fresh[18200], Fresh[18199], Fresh[18198], Fresh[18197], Fresh[18196], Fresh[18195], Fresh[18194], Fresh[18193], Fresh[18192], Fresh[18191], Fresh[18190], Fresh[18189], Fresh[18188], Fresh[18187], Fresh[18186], Fresh[18185], Fresh[18184], Fresh[18183], Fresh[18182], Fresh[18181], Fresh[18180], Fresh[18179], Fresh[18178], Fresh[18177], Fresh[18176], Fresh[18175], Fresh[18174], Fresh[18173], Fresh[18172], Fresh[18171], Fresh[18170], Fresh[18169], Fresh[18168], Fresh[18167], Fresh[18166], Fresh[18165], Fresh[18164], Fresh[18163], Fresh[18162], Fresh[18161], Fresh[18160], Fresh[18159], Fresh[18158], Fresh[18157], Fresh[18156], Fresh[18155], Fresh[18154], Fresh[18153], Fresh[18152], Fresh[18151], Fresh[18150], Fresh[18149], Fresh[18148], Fresh[18147], Fresh[18146], Fresh[18145], Fresh[18144], Fresh[18143], Fresh[18142], Fresh[18141], Fresh[18140], Fresh[18139], Fresh[18138], Fresh[18137], Fresh[18136], Fresh[18135], Fresh[18134], Fresh[18133], Fresh[18132], Fresh[18131], Fresh[18130], Fresh[18129], Fresh[18128], Fresh[18127], Fresh[18126], Fresh[18125], Fresh[18124], Fresh[18123], Fresh[18122], Fresh[18121], Fresh[18120], Fresh[18119], Fresh[18118], Fresh[18117], Fresh[18116], Fresh[18115], Fresh[18114], Fresh[18113], Fresh[18112], Fresh[18111], Fresh[18110], Fresh[18109], Fresh[18108], Fresh[18107], Fresh[18106], Fresh[18105], Fresh[18104], Fresh[18103], Fresh[18102], Fresh[18101], Fresh[18100], Fresh[18099], Fresh[18098], Fresh[18097], Fresh[18096], Fresh[18095], Fresh[18094], Fresh[18093], Fresh[18092], Fresh[18091], Fresh[18090], Fresh[18089], Fresh[18088], Fresh[18087], Fresh[18086], Fresh[18085], Fresh[18084], Fresh[18083], Fresh[18082], Fresh[18081], Fresh[18080], Fresh[18079], Fresh[18078], Fresh[18077], Fresh[18076], Fresh[18075], Fresh[18074], Fresh[18073], Fresh[18072], Fresh[18071], Fresh[18070], Fresh[18069], Fresh[18068], Fresh[18067], Fresh[18066], Fresh[18065], Fresh[18064], Fresh[18063], Fresh[18062], Fresh[18061], Fresh[18060], Fresh[18059], Fresh[18058], Fresh[18057], Fresh[18056], Fresh[18055], Fresh[18054], Fresh[18053], Fresh[18052], Fresh[18051], Fresh[18050], Fresh[18049], Fresh[18048], Fresh[18047], Fresh[18046], Fresh[18045], Fresh[18044], Fresh[18043], Fresh[18042], Fresh[18041], Fresh[18040], Fresh[18039], Fresh[18038], Fresh[18037], Fresh[18036], Fresh[18035], Fresh[18034], Fresh[18033], Fresh[18032], Fresh[18031], Fresh[18030], Fresh[18029], Fresh[18028], Fresh[18027], Fresh[18026], Fresh[18025], Fresh[18024], Fresh[18023], Fresh[18022], Fresh[18021], Fresh[18020], Fresh[18019], Fresh[18018], Fresh[18017], Fresh[18016], Fresh[18015], Fresh[18014], Fresh[18013], Fresh[18012], Fresh[18011], Fresh[18010], Fresh[18009], Fresh[18008], Fresh[18007], Fresh[18006], Fresh[18005], Fresh[18004], Fresh[18003], Fresh[18002], Fresh[18001], Fresh[18000], Fresh[17999], Fresh[17998], Fresh[17997], Fresh[17996], Fresh[17995], Fresh[17994], Fresh[17993], Fresh[17992], Fresh[17991], Fresh[17990], Fresh[17989], Fresh[17988], Fresh[17987], Fresh[17986], Fresh[17985], Fresh[17984], Fresh[17983], Fresh[17982], Fresh[17981], Fresh[17980], Fresh[17979], Fresh[17978], Fresh[17977], Fresh[17976], Fresh[17975], Fresh[17974], Fresh[17973], Fresh[17972], Fresh[17971], Fresh[17970], Fresh[17969], Fresh[17968], Fresh[17967], Fresh[17966], Fresh[17965], Fresh[17964], Fresh[17963], Fresh[17962], Fresh[17961], Fresh[17960], Fresh[17959], Fresh[17958], Fresh[17957], Fresh[17956], Fresh[17955], Fresh[17954], Fresh[17953], Fresh[17952], Fresh[17951], Fresh[17950], Fresh[17949], Fresh[17948], Fresh[17947], Fresh[17946], Fresh[17945], Fresh[17944], Fresh[17943], Fresh[17942], Fresh[17941], Fresh[17940], Fresh[17939], Fresh[17938], Fresh[17937], Fresh[17936], Fresh[17935], Fresh[17934], Fresh[17933], Fresh[17932], Fresh[17931], Fresh[17930], Fresh[17929], Fresh[17928], Fresh[17927], Fresh[17926], Fresh[17925], Fresh[17924], Fresh[17923], Fresh[17922], Fresh[17921], Fresh[17920], Fresh[17919], Fresh[17918], Fresh[17917], Fresh[17916], Fresh[17915], Fresh[17914], Fresh[17913], Fresh[17912], Fresh[17911], Fresh[17910], Fresh[17909], Fresh[17908], Fresh[17907], Fresh[17906], Fresh[17905], Fresh[17904], Fresh[17903], Fresh[17902], Fresh[17901], Fresh[17900], Fresh[17899], Fresh[17898], Fresh[17897], Fresh[17896], Fresh[17895], Fresh[17894], Fresh[17893], Fresh[17892], Fresh[17891], Fresh[17890], Fresh[17889], Fresh[17888], Fresh[17887], Fresh[17886], Fresh[17885], Fresh[17884], Fresh[17883], Fresh[17882], Fresh[17881], Fresh[17880], Fresh[17879], Fresh[17878], Fresh[17877], Fresh[17876], Fresh[17875], Fresh[17874], Fresh[17873], Fresh[17872], Fresh[17871], Fresh[17870], Fresh[17869], Fresh[17868], Fresh[17867], Fresh[17866], Fresh[17865], Fresh[17864], Fresh[17863], Fresh[17862], Fresh[17861], Fresh[17860], Fresh[17859], Fresh[17858], Fresh[17857], Fresh[17856], Fresh[17855], Fresh[17854], Fresh[17853], Fresh[17852], Fresh[17851], Fresh[17850], Fresh[17849], Fresh[17848], Fresh[17847], Fresh[17846], Fresh[17845], Fresh[17844], Fresh[17843], Fresh[17842], Fresh[17841], Fresh[17840], Fresh[17839], Fresh[17838], Fresh[17837], Fresh[17836], Fresh[17835], Fresh[17834], Fresh[17833], Fresh[17832], Fresh[17831], Fresh[17830], Fresh[17829], Fresh[17828], Fresh[17827], Fresh[17826], Fresh[17825], Fresh[17824], Fresh[17823], Fresh[17822], Fresh[17821], Fresh[17820], Fresh[17819], Fresh[17818], Fresh[17817], Fresh[17816], Fresh[17815], Fresh[17814], Fresh[17813], Fresh[17812], Fresh[17811], Fresh[17810], Fresh[17809], Fresh[17808], Fresh[17807], Fresh[17806], Fresh[17805], Fresh[17804], Fresh[17803], Fresh[17802], Fresh[17801], Fresh[17800], Fresh[17799], Fresh[17798], Fresh[17797], Fresh[17796], Fresh[17795], Fresh[17794], Fresh[17793], Fresh[17792], Fresh[17791], Fresh[17790], Fresh[17789], Fresh[17788], Fresh[17787], Fresh[17786], Fresh[17785], Fresh[17784], Fresh[17783], Fresh[17782], Fresh[17781], Fresh[17780], Fresh[17779], Fresh[17778], Fresh[17777], Fresh[17776], Fresh[17775], Fresh[17774], Fresh[17773], Fresh[17772], Fresh[17771], Fresh[17770], Fresh[17769], Fresh[17768], Fresh[17767], Fresh[17766], Fresh[17765], Fresh[17764], Fresh[17763], Fresh[17762], Fresh[17761], Fresh[17760], Fresh[17759], Fresh[17758], Fresh[17757], Fresh[17756], Fresh[17755], Fresh[17754], Fresh[17753], Fresh[17752], Fresh[17751], Fresh[17750], Fresh[17749], Fresh[17748], Fresh[17747], Fresh[17746], Fresh[17745], Fresh[17744], Fresh[17743], Fresh[17742], Fresh[17741], Fresh[17740], Fresh[17739], Fresh[17738], Fresh[17737], Fresh[17736], Fresh[17735], Fresh[17734], Fresh[17733], Fresh[17732], Fresh[17731], Fresh[17730], Fresh[17729], Fresh[17728], Fresh[17727], Fresh[17726], Fresh[17725], Fresh[17724], Fresh[17723], Fresh[17722], Fresh[17721], Fresh[17720], Fresh[17719], Fresh[17718], Fresh[17717], Fresh[17716], Fresh[17715], Fresh[17714], Fresh[17713], Fresh[17712], Fresh[17711], Fresh[17710], Fresh[17709], Fresh[17708], Fresh[17707], Fresh[17706], Fresh[17705], Fresh[17704], Fresh[17703], Fresh[17702], Fresh[17701], Fresh[17700], Fresh[17699], Fresh[17698], Fresh[17697], Fresh[17696], Fresh[17695], Fresh[17694], Fresh[17693], Fresh[17692], Fresh[17691], Fresh[17690], Fresh[17689], Fresh[17688], Fresh[17687], Fresh[17686], Fresh[17685], Fresh[17684], Fresh[17683], Fresh[17682], Fresh[17681], Fresh[17680], Fresh[17679], Fresh[17678], Fresh[17677], Fresh[17676], Fresh[17675], Fresh[17674], Fresh[17673], Fresh[17672], Fresh[17671], Fresh[17670], Fresh[17669], Fresh[17668], Fresh[17667], Fresh[17666], Fresh[17665], Fresh[17664], Fresh[17663], Fresh[17662], Fresh[17661], Fresh[17660], Fresh[17659], Fresh[17658], Fresh[17657], Fresh[17656], Fresh[17655], Fresh[17654], Fresh[17653], Fresh[17652], Fresh[17651], Fresh[17650], Fresh[17649], Fresh[17648], Fresh[17647], Fresh[17646], Fresh[17645], Fresh[17644], Fresh[17643], Fresh[17642], Fresh[17641], Fresh[17640], Fresh[17639], Fresh[17638], Fresh[17637], Fresh[17636], Fresh[17635], Fresh[17634], Fresh[17633], Fresh[17632], Fresh[17631], Fresh[17630], Fresh[17629], Fresh[17628], Fresh[17627], Fresh[17626], Fresh[17625], Fresh[17624], Fresh[17623], Fresh[17622], Fresh[17621], Fresh[17620], Fresh[17619], Fresh[17618], Fresh[17617], Fresh[17616], Fresh[17615], Fresh[17614], Fresh[17613], Fresh[17612], Fresh[17611], Fresh[17610], Fresh[17609], Fresh[17608], Fresh[17607], Fresh[17606], Fresh[17605], Fresh[17604], Fresh[17603], Fresh[17602], Fresh[17601], Fresh[17600], Fresh[17599], Fresh[17598], Fresh[17597], Fresh[17596], Fresh[17595], Fresh[17594], Fresh[17593], Fresh[17592], Fresh[17591], Fresh[17590], Fresh[17589], Fresh[17588], Fresh[17587], Fresh[17586], Fresh[17585], Fresh[17584], Fresh[17583], Fresh[17582], Fresh[17581], Fresh[17580], Fresh[17579], Fresh[17578], Fresh[17577], Fresh[17576], Fresh[17575], Fresh[17574], Fresh[17573], Fresh[17572], Fresh[17571], Fresh[17570], Fresh[17569], Fresh[17568], Fresh[17567], Fresh[17566], Fresh[17565], Fresh[17564], Fresh[17563], Fresh[17562], Fresh[17561], Fresh[17560], Fresh[17559], Fresh[17558], Fresh[17557], Fresh[17556], Fresh[17555], Fresh[17554], Fresh[17553], Fresh[17552], Fresh[17551], Fresh[17550], Fresh[17549], Fresh[17548], Fresh[17547], Fresh[17546], Fresh[17545], Fresh[17544], Fresh[17543], Fresh[17542], Fresh[17541], Fresh[17540], Fresh[17539], Fresh[17538], Fresh[17537], Fresh[17536], Fresh[17535], Fresh[17534], Fresh[17533], Fresh[17532], Fresh[17531], Fresh[17530], Fresh[17529], Fresh[17528], Fresh[17527], Fresh[17526], Fresh[17525], Fresh[17524], Fresh[17523], Fresh[17522], Fresh[17521], Fresh[17520], Fresh[17519], Fresh[17518], Fresh[17517], Fresh[17516], Fresh[17515], Fresh[17514], Fresh[17513], Fresh[17512], Fresh[17511], Fresh[17510], Fresh[17509], Fresh[17508], Fresh[17507], Fresh[17506], Fresh[17505], Fresh[17504], Fresh[17503], Fresh[17502], Fresh[17501], Fresh[17500], Fresh[17499], Fresh[17498], Fresh[17497], Fresh[17496], Fresh[17495], Fresh[17494], Fresh[17493], Fresh[17492], Fresh[17491], Fresh[17490], Fresh[17489], Fresh[17488], Fresh[17487], Fresh[17486], Fresh[17485], Fresh[17484], Fresh[17483], Fresh[17482], Fresh[17481], Fresh[17480], Fresh[17479], Fresh[17478], Fresh[17477], Fresh[17476], Fresh[17475], Fresh[17474], Fresh[17473], Fresh[17472], Fresh[17471], Fresh[17470], Fresh[17469], Fresh[17468], Fresh[17467], Fresh[17466], Fresh[17465], Fresh[17464], Fresh[17463], Fresh[17462], Fresh[17461], Fresh[17460], Fresh[17459], Fresh[17458], Fresh[17457], Fresh[17456], Fresh[17455], Fresh[17454], Fresh[17453], Fresh[17452], Fresh[17451], Fresh[17450], Fresh[17449], Fresh[17448], Fresh[17447], Fresh[17446], Fresh[17445], Fresh[17444], Fresh[17443], Fresh[17442], Fresh[17441], Fresh[17440], Fresh[17439], Fresh[17438], Fresh[17437], Fresh[17436], Fresh[17435], Fresh[17434], Fresh[17433], Fresh[17432], Fresh[17431], Fresh[17430], Fresh[17429], Fresh[17428], Fresh[17427], Fresh[17426], Fresh[17425], Fresh[17424], Fresh[17423], Fresh[17422], Fresh[17421], Fresh[17420], Fresh[17419], Fresh[17418], Fresh[17417], Fresh[17416], Fresh[17415], Fresh[17414], Fresh[17413], Fresh[17412], Fresh[17411], Fresh[17410], Fresh[17409], Fresh[17408], Fresh[17407], Fresh[17406], Fresh[17405], Fresh[17404], Fresh[17403], Fresh[17402], Fresh[17401], Fresh[17400], Fresh[17399], Fresh[17398], Fresh[17397], Fresh[17396], Fresh[17395], Fresh[17394], Fresh[17393], Fresh[17392], Fresh[17391], Fresh[17390], Fresh[17389], Fresh[17388], Fresh[17387], Fresh[17386], Fresh[17385], Fresh[17384], Fresh[17383], Fresh[17382], Fresh[17381], Fresh[17380], Fresh[17379], Fresh[17378], Fresh[17377], Fresh[17376], Fresh[17375], Fresh[17374], Fresh[17373], Fresh[17372], Fresh[17371], Fresh[17370], Fresh[17369], Fresh[17368], Fresh[17367], Fresh[17366], Fresh[17365], Fresh[17364], Fresh[17363], Fresh[17362], Fresh[17361], Fresh[17360], Fresh[17359], Fresh[17358], Fresh[17357], Fresh[17356], Fresh[17355], Fresh[17354], Fresh[17353], Fresh[17352], Fresh[17351], Fresh[17350], Fresh[17349], Fresh[17348], Fresh[17347], Fresh[17346], Fresh[17345], Fresh[17344], Fresh[17343], Fresh[17342], Fresh[17341], Fresh[17340], Fresh[17339], Fresh[17338], Fresh[17337], Fresh[17336], Fresh[17335], Fresh[17334], Fresh[17333], Fresh[17332], Fresh[17331], Fresh[17330], Fresh[17329], Fresh[17328], Fresh[17327], Fresh[17326], Fresh[17325], Fresh[17324], Fresh[17323], Fresh[17322], Fresh[17321], Fresh[17320], Fresh[17319], Fresh[17318], Fresh[17317], Fresh[17316], Fresh[17315], Fresh[17314], Fresh[17313], Fresh[17312], Fresh[17311], Fresh[17310], Fresh[17309], Fresh[17308], Fresh[17307], Fresh[17306], Fresh[17305], Fresh[17304], Fresh[17303], Fresh[17302], Fresh[17301], Fresh[17300], Fresh[17299], Fresh[17298], Fresh[17297], Fresh[17296], Fresh[17295], Fresh[17294], Fresh[17293], Fresh[17292], Fresh[17291], Fresh[17290], Fresh[17289], Fresh[17288], Fresh[17287], Fresh[17286], Fresh[17285], Fresh[17284], Fresh[17283], Fresh[17282], Fresh[17281], Fresh[17280], Fresh[17279], Fresh[17278], Fresh[17277], Fresh[17276], Fresh[17275], Fresh[17274], Fresh[17273], Fresh[17272], Fresh[17271], Fresh[17270], Fresh[17269], Fresh[17268], Fresh[17267], Fresh[17266], Fresh[17265], Fresh[17264], Fresh[17263], Fresh[17262], Fresh[17261], Fresh[17260], Fresh[17259], Fresh[17258], Fresh[17257], Fresh[17256], Fresh[17255], Fresh[17254], Fresh[17253], Fresh[17252], Fresh[17251], Fresh[17250], Fresh[17249], Fresh[17248], Fresh[17247], Fresh[17246], Fresh[17245], Fresh[17244], Fresh[17243], Fresh[17242], Fresh[17241], Fresh[17240], Fresh[17239], Fresh[17238], Fresh[17237], Fresh[17236], Fresh[17235], Fresh[17234], Fresh[17233], Fresh[17232], Fresh[17231], Fresh[17230], Fresh[17229], Fresh[17228], Fresh[17227], Fresh[17226], Fresh[17225], Fresh[17224], Fresh[17223], Fresh[17222], Fresh[17221], Fresh[17220], Fresh[17219], Fresh[17218], Fresh[17217], Fresh[17216], Fresh[17215], Fresh[17214], Fresh[17213], Fresh[17212], Fresh[17211], Fresh[17210], Fresh[17209], Fresh[17208], Fresh[17207], Fresh[17206], Fresh[17205], Fresh[17204], Fresh[17203], Fresh[17202], Fresh[17201], Fresh[17200], Fresh[17199], Fresh[17198], Fresh[17197], Fresh[17196], Fresh[17195], Fresh[17194], Fresh[17193], Fresh[17192], Fresh[17191], Fresh[17190], Fresh[17189], Fresh[17188], Fresh[17187], Fresh[17186], Fresh[17185], Fresh[17184], Fresh[17183], Fresh[17182], Fresh[17181], Fresh[17180], Fresh[17179], Fresh[17178], Fresh[17177], Fresh[17176], Fresh[17175], Fresh[17174], Fresh[17173], Fresh[17172], Fresh[17171], Fresh[17170], Fresh[17169], Fresh[17168], Fresh[17167], Fresh[17166], Fresh[17165], Fresh[17164], Fresh[17163], Fresh[17162], Fresh[17161], Fresh[17160], Fresh[17159], Fresh[17158], Fresh[17157], Fresh[17156], Fresh[17155], Fresh[17154], Fresh[17153], Fresh[17152], Fresh[17151], Fresh[17150], Fresh[17149], Fresh[17148], Fresh[17147], Fresh[17146], Fresh[17145], Fresh[17144], Fresh[17143], Fresh[17142], Fresh[17141], Fresh[17140], Fresh[17139], Fresh[17138], Fresh[17137], Fresh[17136], Fresh[17135], Fresh[17134], Fresh[17133], Fresh[17132], Fresh[17131], Fresh[17130], Fresh[17129], Fresh[17128], Fresh[17127], Fresh[17126], Fresh[17125], Fresh[17124], Fresh[17123], Fresh[17122], Fresh[17121], Fresh[17120], Fresh[17119], Fresh[17118], Fresh[17117], Fresh[17116], Fresh[17115], Fresh[17114], Fresh[17113], Fresh[17112], Fresh[17111], Fresh[17110], Fresh[17109], Fresh[17108], Fresh[17107], Fresh[17106], Fresh[17105], Fresh[17104], Fresh[17103], Fresh[17102], Fresh[17101], Fresh[17100], Fresh[17099], Fresh[17098], Fresh[17097], Fresh[17096], Fresh[17095], Fresh[17094], Fresh[17093], Fresh[17092], Fresh[17091], Fresh[17090], Fresh[17089], Fresh[17088], Fresh[17087], Fresh[17086], Fresh[17085], Fresh[17084], Fresh[17083], Fresh[17082], Fresh[17081], Fresh[17080], Fresh[17079], Fresh[17078], Fresh[17077], Fresh[17076], Fresh[17075], Fresh[17074], Fresh[17073], Fresh[17072], Fresh[17071], Fresh[17070], Fresh[17069], Fresh[17068], Fresh[17067], Fresh[17066], Fresh[17065], Fresh[17064], Fresh[17063], Fresh[17062], Fresh[17061], Fresh[17060], Fresh[17059], Fresh[17058], Fresh[17057], Fresh[17056], Fresh[17055], Fresh[17054], Fresh[17053], Fresh[17052], Fresh[17051], Fresh[17050], Fresh[17049], Fresh[17048], Fresh[17047], Fresh[17046], Fresh[17045], Fresh[17044], Fresh[17043], Fresh[17042], Fresh[17041], Fresh[17040], Fresh[17039], Fresh[17038], Fresh[17037], Fresh[17036], Fresh[17035], Fresh[17034], Fresh[17033], Fresh[17032], Fresh[17031], Fresh[17030], Fresh[17029], Fresh[17028], Fresh[17027], Fresh[17026], Fresh[17025], Fresh[17024], Fresh[17023], Fresh[17022], Fresh[17021], Fresh[17020], Fresh[17019], Fresh[17018], Fresh[17017], Fresh[17016], Fresh[17015], Fresh[17014], Fresh[17013], Fresh[17012], Fresh[17011], Fresh[17010], Fresh[17009], Fresh[17008], Fresh[17007], Fresh[17006], Fresh[17005], Fresh[17004], Fresh[17003], Fresh[17002], Fresh[17001], Fresh[17000], Fresh[16999], Fresh[16998], Fresh[16997], Fresh[16996], Fresh[16995], Fresh[16994], Fresh[16993], Fresh[16992], Fresh[16991], Fresh[16990], Fresh[16989], Fresh[16988], Fresh[16987], Fresh[16986], Fresh[16985], Fresh[16984], Fresh[16983], Fresh[16982], Fresh[16981], Fresh[16980], Fresh[16979], Fresh[16978], Fresh[16977], Fresh[16976], Fresh[16975], Fresh[16974], Fresh[16973], Fresh[16972], Fresh[16971], Fresh[16970], Fresh[16969], Fresh[16968], Fresh[16967], Fresh[16966], Fresh[16965], Fresh[16964], Fresh[16963], Fresh[16962], Fresh[16961], Fresh[16960], Fresh[16959], Fresh[16958], Fresh[16957], Fresh[16956], Fresh[16955], Fresh[16954], Fresh[16953], Fresh[16952], Fresh[16951], Fresh[16950], Fresh[16949], Fresh[16948], Fresh[16947], Fresh[16946], Fresh[16945], Fresh[16944], Fresh[16943], Fresh[16942], Fresh[16941], Fresh[16940], Fresh[16939], Fresh[16938], Fresh[16937], Fresh[16936], Fresh[16935], Fresh[16934], Fresh[16933], Fresh[16932], Fresh[16931], Fresh[16930], Fresh[16929], Fresh[16928], Fresh[16927], Fresh[16926], Fresh[16925], Fresh[16924], Fresh[16923], Fresh[16922], Fresh[16921], Fresh[16920], Fresh[16919], Fresh[16918], Fresh[16917], Fresh[16916], Fresh[16915], Fresh[16914], Fresh[16913], Fresh[16912], Fresh[16911], Fresh[16910], Fresh[16909], Fresh[16908], Fresh[16907], Fresh[16906], Fresh[16905], Fresh[16904], Fresh[16903], Fresh[16902], Fresh[16901], Fresh[16900], Fresh[16899], Fresh[16898], Fresh[16897], Fresh[16896], Fresh[16895], Fresh[16894], Fresh[16893], Fresh[16892], Fresh[16891], Fresh[16890], Fresh[16889], Fresh[16888], Fresh[16887], Fresh[16886], Fresh[16885], Fresh[16884], Fresh[16883], Fresh[16882], Fresh[16881], Fresh[16880], Fresh[16879], Fresh[16878], Fresh[16877], Fresh[16876], Fresh[16875], Fresh[16874], Fresh[16873], Fresh[16872], Fresh[16871], Fresh[16870], Fresh[16869], Fresh[16868], Fresh[16867], Fresh[16866], Fresh[16865], Fresh[16864], Fresh[16863], Fresh[16862], Fresh[16861], Fresh[16860], Fresh[16859], Fresh[16858], Fresh[16857], Fresh[16856], Fresh[16855], Fresh[16854], Fresh[16853], Fresh[16852], Fresh[16851], Fresh[16850], Fresh[16849], Fresh[16848], Fresh[16847], Fresh[16846], Fresh[16845], Fresh[16844], Fresh[16843], Fresh[16842], Fresh[16841], Fresh[16840], Fresh[16839], Fresh[16838], Fresh[16837], Fresh[16836], Fresh[16835], Fresh[16834], Fresh[16833], Fresh[16832], Fresh[16831], Fresh[16830], Fresh[16829], Fresh[16828], Fresh[16827], Fresh[16826], Fresh[16825], Fresh[16824], Fresh[16823], Fresh[16822], Fresh[16821], Fresh[16820], Fresh[16819], Fresh[16818], Fresh[16817], Fresh[16816], Fresh[16815], Fresh[16814], Fresh[16813], Fresh[16812], Fresh[16811], Fresh[16810], Fresh[16809], Fresh[16808], Fresh[16807], Fresh[16806], Fresh[16805], Fresh[16804], Fresh[16803], Fresh[16802], Fresh[16801], Fresh[16800], Fresh[16799], Fresh[16798], Fresh[16797], Fresh[16796], Fresh[16795], Fresh[16794], Fresh[16793], Fresh[16792], Fresh[16791], Fresh[16790], Fresh[16789], Fresh[16788], Fresh[16787], Fresh[16786], Fresh[16785], Fresh[16784], Fresh[16783], Fresh[16782], Fresh[16781], Fresh[16780], Fresh[16779], Fresh[16778], Fresh[16777], Fresh[16776], Fresh[16775], Fresh[16774], Fresh[16773], Fresh[16772], Fresh[16771], Fresh[16770], Fresh[16769], Fresh[16768], Fresh[16767], Fresh[16766], Fresh[16765], Fresh[16764], Fresh[16763], Fresh[16762], Fresh[16761], Fresh[16760], Fresh[16759], Fresh[16758], Fresh[16757], Fresh[16756], Fresh[16755], Fresh[16754], Fresh[16753], Fresh[16752], Fresh[16751], Fresh[16750], Fresh[16749], Fresh[16748], Fresh[16747], Fresh[16746], Fresh[16745], Fresh[16744], Fresh[16743], Fresh[16742], Fresh[16741], Fresh[16740], Fresh[16739], Fresh[16738], Fresh[16737], Fresh[16736], Fresh[16735], Fresh[16734], Fresh[16733], Fresh[16732], Fresh[16731], Fresh[16730], Fresh[16729], Fresh[16728], Fresh[16727], Fresh[16726], Fresh[16725], Fresh[16724], Fresh[16723], Fresh[16722], Fresh[16721], Fresh[16720], Fresh[16719], Fresh[16718], Fresh[16717], Fresh[16716], Fresh[16715], Fresh[16714], Fresh[16713], Fresh[16712], Fresh[16711], Fresh[16710], Fresh[16709], Fresh[16708], Fresh[16707], Fresh[16706], Fresh[16705], Fresh[16704], Fresh[16703], Fresh[16702], Fresh[16701], Fresh[16700], Fresh[16699], Fresh[16698], Fresh[16697], Fresh[16696], Fresh[16695], Fresh[16694], Fresh[16693], Fresh[16692], Fresh[16691], Fresh[16690], Fresh[16689], Fresh[16688], Fresh[16687], Fresh[16686], Fresh[16685], Fresh[16684], Fresh[16683], Fresh[16682], Fresh[16681], Fresh[16680], Fresh[16679], Fresh[16678], Fresh[16677], Fresh[16676], Fresh[16675], Fresh[16674], Fresh[16673], Fresh[16672], Fresh[16671], Fresh[16670], Fresh[16669], Fresh[16668], Fresh[16667], Fresh[16666], Fresh[16665], Fresh[16664], Fresh[16663], Fresh[16662], Fresh[16661], Fresh[16660], Fresh[16659], Fresh[16658], Fresh[16657], Fresh[16656], Fresh[16655], Fresh[16654], Fresh[16653], Fresh[16652], Fresh[16651], Fresh[16650], Fresh[16649], Fresh[16648], Fresh[16647], Fresh[16646], Fresh[16645], Fresh[16644], Fresh[16643], Fresh[16642], Fresh[16641], Fresh[16640], Fresh[16639], Fresh[16638], Fresh[16637], Fresh[16636], Fresh[16635], Fresh[16634], Fresh[16633], Fresh[16632], Fresh[16631], Fresh[16630], Fresh[16629], Fresh[16628], Fresh[16627], Fresh[16626], Fresh[16625], Fresh[16624], Fresh[16623], Fresh[16622], Fresh[16621], Fresh[16620], Fresh[16619], Fresh[16618], Fresh[16617], Fresh[16616], Fresh[16615], Fresh[16614], Fresh[16613], Fresh[16612], Fresh[16611], Fresh[16610], Fresh[16609], Fresh[16608], Fresh[16607], Fresh[16606], Fresh[16605], Fresh[16604], Fresh[16603], Fresh[16602], Fresh[16601], Fresh[16600], Fresh[16599], Fresh[16598], Fresh[16597], Fresh[16596], Fresh[16595], Fresh[16594], Fresh[16593], Fresh[16592], Fresh[16591], Fresh[16590], Fresh[16589], Fresh[16588], Fresh[16587], Fresh[16586], Fresh[16585], Fresh[16584], Fresh[16583], Fresh[16582], Fresh[16581], Fresh[16580], Fresh[16579], Fresh[16578], Fresh[16577], Fresh[16576], Fresh[16575], Fresh[16574], Fresh[16573], Fresh[16572], Fresh[16571], Fresh[16570], Fresh[16569], Fresh[16568], Fresh[16567], Fresh[16566], Fresh[16565], Fresh[16564], Fresh[16563], Fresh[16562], Fresh[16561], Fresh[16560], Fresh[16559], Fresh[16558], Fresh[16557], Fresh[16556], Fresh[16555], Fresh[16554], Fresh[16553], Fresh[16552], Fresh[16551], Fresh[16550], Fresh[16549], Fresh[16548], Fresh[16547], Fresh[16546], Fresh[16545], Fresh[16544], Fresh[16543], Fresh[16542], Fresh[16541], Fresh[16540], Fresh[16539], Fresh[16538], Fresh[16537], Fresh[16536], Fresh[16535], Fresh[16534], Fresh[16533], Fresh[16532], Fresh[16531], Fresh[16530], Fresh[16529], Fresh[16528], Fresh[16527], Fresh[16526], Fresh[16525], Fresh[16524], Fresh[16523], Fresh[16522], Fresh[16521], Fresh[16520], Fresh[16519], Fresh[16518], Fresh[16517], Fresh[16516], Fresh[16515], Fresh[16514], Fresh[16513], Fresh[16512], Fresh[16511], Fresh[16510], Fresh[16509], Fresh[16508], Fresh[16507], Fresh[16506], Fresh[16505], Fresh[16504], Fresh[16503], Fresh[16502], Fresh[16501], Fresh[16500], Fresh[16499], Fresh[16498], Fresh[16497], Fresh[16496], Fresh[16495], Fresh[16494], Fresh[16493], Fresh[16492], Fresh[16491], Fresh[16490], Fresh[16489], Fresh[16488], Fresh[16487], Fresh[16486], Fresh[16485], Fresh[16484], Fresh[16483], Fresh[16482], Fresh[16481], Fresh[16480], Fresh[16479], Fresh[16478], Fresh[16477], Fresh[16476], Fresh[16475], Fresh[16474], Fresh[16473], Fresh[16472], Fresh[16471], Fresh[16470], Fresh[16469], Fresh[16468], Fresh[16467], Fresh[16466], Fresh[16465], Fresh[16464], Fresh[16463], Fresh[16462], Fresh[16461], Fresh[16460], Fresh[16459], Fresh[16458], Fresh[16457], Fresh[16456], Fresh[16455], Fresh[16454], Fresh[16453], Fresh[16452], Fresh[16451], Fresh[16450], Fresh[16449], Fresh[16448], Fresh[16447], Fresh[16446], Fresh[16445], Fresh[16444], Fresh[16443], Fresh[16442], Fresh[16441], Fresh[16440], Fresh[16439], Fresh[16438], Fresh[16437], Fresh[16436], Fresh[16435], Fresh[16434], Fresh[16433], Fresh[16432], Fresh[16431], Fresh[16430], Fresh[16429], Fresh[16428], Fresh[16427], Fresh[16426], Fresh[16425], Fresh[16424], Fresh[16423], Fresh[16422], Fresh[16421], Fresh[16420], Fresh[16419], Fresh[16418], Fresh[16417], Fresh[16416], Fresh[16415], Fresh[16414], Fresh[16413], Fresh[16412], Fresh[16411], Fresh[16410], Fresh[16409], Fresh[16408], Fresh[16407], Fresh[16406], Fresh[16405], Fresh[16404], Fresh[16403], Fresh[16402], Fresh[16401], Fresh[16400], Fresh[16399], Fresh[16398], Fresh[16397], Fresh[16396], Fresh[16395], Fresh[16394], Fresh[16393], Fresh[16392], Fresh[16391], Fresh[16390], Fresh[16389], Fresh[16388], Fresh[16387], Fresh[16386], Fresh[16385], Fresh[16384], Fresh[16383], Fresh[16382], Fresh[16381], Fresh[16380], Fresh[16379], Fresh[16378], Fresh[16377], Fresh[16376], Fresh[16375], Fresh[16374], Fresh[16373], Fresh[16372], Fresh[16371], Fresh[16370], Fresh[16369], Fresh[16368], Fresh[16367], Fresh[16366], Fresh[16365], Fresh[16364], Fresh[16363], Fresh[16362], Fresh[16361], Fresh[16360], Fresh[16359], Fresh[16358], Fresh[16357], Fresh[16356], Fresh[16355], Fresh[16354], Fresh[16353], Fresh[16352], Fresh[16351], Fresh[16350], Fresh[16349], Fresh[16348], Fresh[16347], Fresh[16346], Fresh[16345], Fresh[16344], Fresh[16343], Fresh[16342], Fresh[16341], Fresh[16340], Fresh[16339], Fresh[16338], Fresh[16337], Fresh[16336], Fresh[16335], Fresh[16334], Fresh[16333], Fresh[16332], Fresh[16331], Fresh[16330], Fresh[16329], Fresh[16328], Fresh[16327], Fresh[16326], Fresh[16325], Fresh[16324], Fresh[16323], Fresh[16322], Fresh[16321], Fresh[16320], Fresh[16319], Fresh[16318], Fresh[16317], Fresh[16316], Fresh[16315], Fresh[16314], Fresh[16313], Fresh[16312], Fresh[16311], Fresh[16310], Fresh[16309], Fresh[16308], Fresh[16307], Fresh[16306], Fresh[16305], Fresh[16304], Fresh[16303], Fresh[16302], Fresh[16301], Fresh[16300], Fresh[16299], Fresh[16298], Fresh[16297], Fresh[16296], Fresh[16295], Fresh[16294], Fresh[16293], Fresh[16292], Fresh[16291], Fresh[16290], Fresh[16289], Fresh[16288], Fresh[16287], Fresh[16286], Fresh[16285], Fresh[16284], Fresh[16283], Fresh[16282], Fresh[16281], Fresh[16280], Fresh[16279], Fresh[16278], Fresh[16277], Fresh[16276], Fresh[16275], Fresh[16274], Fresh[16273], Fresh[16272], Fresh[16271], Fresh[16270], Fresh[16269], Fresh[16268], Fresh[16267], Fresh[16266], Fresh[16265], Fresh[16264], Fresh[16263], Fresh[16262], Fresh[16261], Fresh[16260], Fresh[16259], Fresh[16258], Fresh[16257], Fresh[16256], Fresh[16255], Fresh[16254], Fresh[16253], Fresh[16252], Fresh[16251], Fresh[16250], Fresh[16249], Fresh[16248], Fresh[16247], Fresh[16246], Fresh[16245], Fresh[16244], Fresh[16243], Fresh[16242], Fresh[16241], Fresh[16240], Fresh[16239], Fresh[16238], Fresh[16237], Fresh[16236], Fresh[16235], Fresh[16234], Fresh[16233], Fresh[16232], Fresh[16231], Fresh[16230], Fresh[16229], Fresh[16228], Fresh[16227], Fresh[16226], Fresh[16225], Fresh[16224], Fresh[16223], Fresh[16222], Fresh[16221], Fresh[16220], Fresh[16219], Fresh[16218], Fresh[16217], Fresh[16216], Fresh[16215], Fresh[16214], Fresh[16213], Fresh[16212], Fresh[16211], Fresh[16210], Fresh[16209], Fresh[16208], Fresh[16207], Fresh[16206], Fresh[16205], Fresh[16204], Fresh[16203], Fresh[16202], Fresh[16201], Fresh[16200], Fresh[16199], Fresh[16198], Fresh[16197], Fresh[16196], Fresh[16195], Fresh[16194], Fresh[16193], Fresh[16192], Fresh[16191], Fresh[16190], Fresh[16189], Fresh[16188], Fresh[16187], Fresh[16186], Fresh[16185], Fresh[16184], Fresh[16183], Fresh[16182], Fresh[16181], Fresh[16180], Fresh[16179], Fresh[16178], Fresh[16177], Fresh[16176], Fresh[16175], Fresh[16174], Fresh[16173], Fresh[16172], Fresh[16171], Fresh[16170], Fresh[16169], Fresh[16168], Fresh[16167], Fresh[16166], Fresh[16165], Fresh[16164], Fresh[16163], Fresh[16162], Fresh[16161], Fresh[16160], Fresh[16159], Fresh[16158], Fresh[16157], Fresh[16156], Fresh[16155], Fresh[16154], Fresh[16153], Fresh[16152], Fresh[16151], Fresh[16150], Fresh[16149], Fresh[16148], Fresh[16147], Fresh[16146], Fresh[16145], Fresh[16144], Fresh[16143], Fresh[16142], Fresh[16141], Fresh[16140], Fresh[16139], Fresh[16138], Fresh[16137], Fresh[16136], Fresh[16135], Fresh[16134], Fresh[16133], Fresh[16132], Fresh[16131], Fresh[16130], Fresh[16129], Fresh[16128], Fresh[16127], Fresh[16126], Fresh[16125], Fresh[16124], Fresh[16123], Fresh[16122], Fresh[16121], Fresh[16120], Fresh[16119], Fresh[16118], Fresh[16117], Fresh[16116], Fresh[16115], Fresh[16114], Fresh[16113], Fresh[16112], Fresh[16111], Fresh[16110], Fresh[16109], Fresh[16108], Fresh[16107], Fresh[16106], Fresh[16105], Fresh[16104], Fresh[16103], Fresh[16102], Fresh[16101], Fresh[16100], Fresh[16099], Fresh[16098], Fresh[16097], Fresh[16096], Fresh[16095], Fresh[16094], Fresh[16093], Fresh[16092], Fresh[16091], Fresh[16090], Fresh[16089], Fresh[16088], Fresh[16087], Fresh[16086], Fresh[16085], Fresh[16084], Fresh[16083], Fresh[16082], Fresh[16081], Fresh[16080], Fresh[16079], Fresh[16078], Fresh[16077], Fresh[16076], Fresh[16075], Fresh[16074], Fresh[16073], Fresh[16072], Fresh[16071], Fresh[16070], Fresh[16069], Fresh[16068], Fresh[16067], Fresh[16066], Fresh[16065], Fresh[16064], Fresh[16063], Fresh[16062], Fresh[16061], Fresh[16060], Fresh[16059], Fresh[16058], Fresh[16057], Fresh[16056], Fresh[16055], Fresh[16054], Fresh[16053], Fresh[16052], Fresh[16051], Fresh[16050], Fresh[16049], Fresh[16048], Fresh[16047], Fresh[16046], Fresh[16045], Fresh[16044], Fresh[16043], Fresh[16042], Fresh[16041], Fresh[16040], Fresh[16039], Fresh[16038], Fresh[16037], Fresh[16036], Fresh[16035], Fresh[16034], Fresh[16033], Fresh[16032], Fresh[16031], Fresh[16030], Fresh[16029], Fresh[16028], Fresh[16027], Fresh[16026], Fresh[16025], Fresh[16024], Fresh[16023], Fresh[16022], Fresh[16021], Fresh[16020], Fresh[16019], Fresh[16018], Fresh[16017], Fresh[16016], Fresh[16015], Fresh[16014], Fresh[16013], Fresh[16012], Fresh[16011], Fresh[16010], Fresh[16009], Fresh[16008], Fresh[16007], Fresh[16006], Fresh[16005], Fresh[16004], Fresh[16003], Fresh[16002], Fresh[16001], Fresh[16000], Fresh[15999], Fresh[15998], Fresh[15997], Fresh[15996], Fresh[15995], Fresh[15994], Fresh[15993], Fresh[15992], Fresh[15991], Fresh[15990], Fresh[15989], Fresh[15988], Fresh[15987], Fresh[15986], Fresh[15985], Fresh[15984], Fresh[15983], Fresh[15982], Fresh[15981], Fresh[15980], Fresh[15979], Fresh[15978], Fresh[15977], Fresh[15976], Fresh[15975], Fresh[15974], Fresh[15973], Fresh[15972], Fresh[15971], Fresh[15970], Fresh[15969], Fresh[15968], Fresh[15967], Fresh[15966], Fresh[15965], Fresh[15964], Fresh[15963], Fresh[15962], Fresh[15961], Fresh[15960], Fresh[15959], Fresh[15958], Fresh[15957], Fresh[15956], Fresh[15955], Fresh[15954], Fresh[15953], Fresh[15952], Fresh[15951], Fresh[15950], Fresh[15949], Fresh[15948], Fresh[15947], Fresh[15946], Fresh[15945], Fresh[15944], Fresh[15943], Fresh[15942], Fresh[15941], Fresh[15940], Fresh[15939], Fresh[15938], Fresh[15937], Fresh[15936], Fresh[15935], Fresh[15934], Fresh[15933], Fresh[15932], Fresh[15931], Fresh[15930], Fresh[15929], Fresh[15928], Fresh[15927], Fresh[15926], Fresh[15925], Fresh[15924], Fresh[15923], Fresh[15922], Fresh[15921], Fresh[15920], Fresh[15919], Fresh[15918], Fresh[15917], Fresh[15916], Fresh[15915], Fresh[15914], Fresh[15913], Fresh[15912], Fresh[15911], Fresh[15910], Fresh[15909], Fresh[15908], Fresh[15907], Fresh[15906], Fresh[15905], Fresh[15904], Fresh[15903], Fresh[15902], Fresh[15901], Fresh[15900], Fresh[15899], Fresh[15898], Fresh[15897], Fresh[15896], Fresh[15895], Fresh[15894], Fresh[15893], Fresh[15892], Fresh[15891], Fresh[15890], Fresh[15889], Fresh[15888], Fresh[15887], Fresh[15886], Fresh[15885], Fresh[15884], Fresh[15883], Fresh[15882], Fresh[15881], Fresh[15880], Fresh[15879], Fresh[15878], Fresh[15877], Fresh[15876], Fresh[15875], Fresh[15874], Fresh[15873], Fresh[15872], Fresh[15871], Fresh[15870], Fresh[15869], Fresh[15868], Fresh[15867], Fresh[15866], Fresh[15865], Fresh[15864], Fresh[15863], Fresh[15862], Fresh[15861], Fresh[15860], Fresh[15859], Fresh[15858], Fresh[15857], Fresh[15856], Fresh[15855], Fresh[15854], Fresh[15853], Fresh[15852], Fresh[15851], Fresh[15850], Fresh[15849], Fresh[15848], Fresh[15847], Fresh[15846], Fresh[15845], Fresh[15844], Fresh[15843], Fresh[15842], Fresh[15841], Fresh[15840], Fresh[15839], Fresh[15838], Fresh[15837], Fresh[15836], Fresh[15835], Fresh[15834], Fresh[15833], Fresh[15832], Fresh[15831], Fresh[15830], Fresh[15829], Fresh[15828], Fresh[15827], Fresh[15826], Fresh[15825], Fresh[15824], Fresh[15823], Fresh[15822], Fresh[15821], Fresh[15820], Fresh[15819], Fresh[15818], Fresh[15817], Fresh[15816], Fresh[15815], Fresh[15814], Fresh[15813], Fresh[15812], Fresh[15811], Fresh[15810], Fresh[15809], Fresh[15808], Fresh[15807], Fresh[15806], Fresh[15805], Fresh[15804], Fresh[15803], Fresh[15802], Fresh[15801], Fresh[15800], Fresh[15799], Fresh[15798], Fresh[15797], Fresh[15796], Fresh[15795], Fresh[15794], Fresh[15793], Fresh[15792], Fresh[15791], Fresh[15790], Fresh[15789], Fresh[15788], Fresh[15787], Fresh[15786], Fresh[15785], Fresh[15784], Fresh[15783], Fresh[15782], Fresh[15781], Fresh[15780], Fresh[15779], Fresh[15778], Fresh[15777], Fresh[15776], Fresh[15775], Fresh[15774], Fresh[15773], Fresh[15772], Fresh[15771], Fresh[15770], Fresh[15769], Fresh[15768], Fresh[15767], Fresh[15766], Fresh[15765], Fresh[15764], Fresh[15763], Fresh[15762], Fresh[15761], Fresh[15760], Fresh[15759], Fresh[15758], Fresh[15757], Fresh[15756], Fresh[15755], Fresh[15754], Fresh[15753], Fresh[15752], Fresh[15751], Fresh[15750], Fresh[15749], Fresh[15748], Fresh[15747], Fresh[15746], Fresh[15745], Fresh[15744], Fresh[15743], Fresh[15742], Fresh[15741], Fresh[15740], Fresh[15739], Fresh[15738], Fresh[15737], Fresh[15736], Fresh[15735], Fresh[15734], Fresh[15733], Fresh[15732], Fresh[15731], Fresh[15730], Fresh[15729], Fresh[15728], Fresh[15727], Fresh[15726], Fresh[15725], Fresh[15724], Fresh[15723], Fresh[15722], Fresh[15721], Fresh[15720], Fresh[15719], Fresh[15718], Fresh[15717], Fresh[15716], Fresh[15715], Fresh[15714], Fresh[15713], Fresh[15712], Fresh[15711], Fresh[15710], Fresh[15709], Fresh[15708], Fresh[15707], Fresh[15706], Fresh[15705], Fresh[15704], Fresh[15703], Fresh[15702], Fresh[15701], Fresh[15700], Fresh[15699], Fresh[15698], Fresh[15697], Fresh[15696], Fresh[15695], Fresh[15694], Fresh[15693], Fresh[15692], Fresh[15691], Fresh[15690], Fresh[15689], Fresh[15688], Fresh[15687], Fresh[15686], Fresh[15685], Fresh[15684], Fresh[15683], Fresh[15682], Fresh[15681], Fresh[15680], Fresh[15679], Fresh[15678], Fresh[15677], Fresh[15676], Fresh[15675], Fresh[15674], Fresh[15673], Fresh[15672], Fresh[15671], Fresh[15670], Fresh[15669], Fresh[15668], Fresh[15667], Fresh[15666], Fresh[15665], Fresh[15664], Fresh[15663], Fresh[15662], Fresh[15661], Fresh[15660], Fresh[15659], Fresh[15658], Fresh[15657], Fresh[15656], Fresh[15655], Fresh[15654], Fresh[15653], Fresh[15652], Fresh[15651], Fresh[15650], Fresh[15649], Fresh[15648], Fresh[15647], Fresh[15646], Fresh[15645], Fresh[15644], Fresh[15643], Fresh[15642], Fresh[15641], Fresh[15640], Fresh[15639], Fresh[15638], Fresh[15637], Fresh[15636], Fresh[15635], Fresh[15634], Fresh[15633], Fresh[15632], Fresh[15631], Fresh[15630], Fresh[15629], Fresh[15628], Fresh[15627], Fresh[15626], Fresh[15625], Fresh[15624], Fresh[15623], Fresh[15622], Fresh[15621], Fresh[15620], Fresh[15619], Fresh[15618], Fresh[15617], Fresh[15616], Fresh[15615], Fresh[15614], Fresh[15613], Fresh[15612], Fresh[15611], Fresh[15610], Fresh[15609], Fresh[15608], Fresh[15607], Fresh[15606], Fresh[15605], Fresh[15604], Fresh[15603], Fresh[15602], Fresh[15601], Fresh[15600], Fresh[15599], Fresh[15598], Fresh[15597], Fresh[15596], Fresh[15595], Fresh[15594], Fresh[15593], Fresh[15592], Fresh[15591], Fresh[15590], Fresh[15589], Fresh[15588], Fresh[15587], Fresh[15586], Fresh[15585], Fresh[15584], Fresh[15583], Fresh[15582], Fresh[15581], Fresh[15580], Fresh[15579], Fresh[15578], Fresh[15577], Fresh[15576], Fresh[15575], Fresh[15574], Fresh[15573], Fresh[15572], Fresh[15571], Fresh[15570], Fresh[15569], Fresh[15568], Fresh[15567], Fresh[15566], Fresh[15565], Fresh[15564], Fresh[15563], Fresh[15562], Fresh[15561], Fresh[15560], Fresh[15559], Fresh[15558], Fresh[15557], Fresh[15556], Fresh[15555], Fresh[15554], Fresh[15553], Fresh[15552], Fresh[15551], Fresh[15550], Fresh[15549], Fresh[15548], Fresh[15547], Fresh[15546], Fresh[15545], Fresh[15544], Fresh[15543], Fresh[15542], Fresh[15541], Fresh[15540], Fresh[15539], Fresh[15538], Fresh[15537], Fresh[15536], Fresh[15535], Fresh[15534], Fresh[15533], Fresh[15532], Fresh[15531], Fresh[15530], Fresh[15529], Fresh[15528], Fresh[15527], Fresh[15526], Fresh[15525], Fresh[15524], Fresh[15523], Fresh[15522], Fresh[15521], Fresh[15520], Fresh[15519], Fresh[15518], Fresh[15517], Fresh[15516], Fresh[15515], Fresh[15514], Fresh[15513], Fresh[15512], Fresh[15511], Fresh[15510], Fresh[15509], Fresh[15508], Fresh[15507], Fresh[15506], Fresh[15505], Fresh[15504], Fresh[15503], Fresh[15502], Fresh[15501], Fresh[15500], Fresh[15499], Fresh[15498], Fresh[15497], Fresh[15496], Fresh[15495], Fresh[15494], Fresh[15493], Fresh[15492], Fresh[15491], Fresh[15490], Fresh[15489], Fresh[15488], Fresh[15487], Fresh[15486], Fresh[15485], Fresh[15484], Fresh[15483], Fresh[15482], Fresh[15481], Fresh[15480], Fresh[15479], Fresh[15478], Fresh[15477], Fresh[15476], Fresh[15475], Fresh[15474], Fresh[15473], Fresh[15472], Fresh[15471], Fresh[15470], Fresh[15469], Fresh[15468], Fresh[15467], Fresh[15466], Fresh[15465], Fresh[15464], Fresh[15463], Fresh[15462], Fresh[15461], Fresh[15460], Fresh[15459], Fresh[15458], Fresh[15457], Fresh[15456], Fresh[15455], Fresh[15454], Fresh[15453], Fresh[15452], Fresh[15451], Fresh[15450], Fresh[15449], Fresh[15448], Fresh[15447], Fresh[15446], Fresh[15445], Fresh[15444], Fresh[15443], Fresh[15442], Fresh[15441], Fresh[15440], Fresh[15439], Fresh[15438], Fresh[15437], Fresh[15436], Fresh[15435], Fresh[15434], Fresh[15433], Fresh[15432], Fresh[15431], Fresh[15430], Fresh[15429], Fresh[15428], Fresh[15427], Fresh[15426], Fresh[15425], Fresh[15424], Fresh[15423], Fresh[15422], Fresh[15421], Fresh[15420], Fresh[15419], Fresh[15418], Fresh[15417], Fresh[15416], Fresh[15415], Fresh[15414], Fresh[15413], Fresh[15412], Fresh[15411], Fresh[15410], Fresh[15409], Fresh[15408], Fresh[15407], Fresh[15406], Fresh[15405], Fresh[15404], Fresh[15403], Fresh[15402], Fresh[15401], Fresh[15400], Fresh[15399], Fresh[15398], Fresh[15397], Fresh[15396], Fresh[15395], Fresh[15394], Fresh[15393], Fresh[15392], Fresh[15391], Fresh[15390], Fresh[15389], Fresh[15388], Fresh[15387], Fresh[15386], Fresh[15385], Fresh[15384], Fresh[15383], Fresh[15382], Fresh[15381], Fresh[15380], Fresh[15379], Fresh[15378], Fresh[15377], Fresh[15376], Fresh[15375], Fresh[15374], Fresh[15373], Fresh[15372], Fresh[15371], Fresh[15370], Fresh[15369], Fresh[15368], Fresh[15367], Fresh[15366], Fresh[15365], Fresh[15364], Fresh[15363], Fresh[15362], Fresh[15361], Fresh[15360], Fresh[15359], Fresh[15358], Fresh[15357], Fresh[15356], Fresh[15355], Fresh[15354], Fresh[15353], Fresh[15352], Fresh[15351], Fresh[15350], Fresh[15349], Fresh[15348], Fresh[15347], Fresh[15346], Fresh[15345], Fresh[15344], Fresh[15343], Fresh[15342], Fresh[15341], Fresh[15340], Fresh[15339], Fresh[15338], Fresh[15337], Fresh[15336], Fresh[15335], Fresh[15334], Fresh[15333], Fresh[15332], Fresh[15331], Fresh[15330], Fresh[15329], Fresh[15328], Fresh[15327], Fresh[15326], Fresh[15325], Fresh[15324], Fresh[15323], Fresh[15322], Fresh[15321], Fresh[15320], Fresh[15319], Fresh[15318], Fresh[15317], Fresh[15316], Fresh[15315], Fresh[15314], Fresh[15313], Fresh[15312], Fresh[15311], Fresh[15310], Fresh[15309], Fresh[15308], Fresh[15307], Fresh[15306], Fresh[15305], Fresh[15304], Fresh[15303], Fresh[15302], Fresh[15301], Fresh[15300], Fresh[15299], Fresh[15298], Fresh[15297], Fresh[15296], Fresh[15295], Fresh[15294], Fresh[15293], Fresh[15292], Fresh[15291], Fresh[15290], Fresh[15289], Fresh[15288], Fresh[15287], Fresh[15286], Fresh[15285], Fresh[15284], Fresh[15283], Fresh[15282], Fresh[15281], Fresh[15280], Fresh[15279], Fresh[15278], Fresh[15277], Fresh[15276], Fresh[15275], Fresh[15274], Fresh[15273], Fresh[15272], Fresh[15271], Fresh[15270], Fresh[15269], Fresh[15268], Fresh[15267], Fresh[15266], Fresh[15265], Fresh[15264], Fresh[15263], Fresh[15262], Fresh[15261], Fresh[15260], Fresh[15259], Fresh[15258], Fresh[15257], Fresh[15256], Fresh[15255], Fresh[15254], Fresh[15253], Fresh[15252], Fresh[15251], Fresh[15250], Fresh[15249], Fresh[15248], Fresh[15247], Fresh[15246], Fresh[15245], Fresh[15244], Fresh[15243], Fresh[15242], Fresh[15241], Fresh[15240], Fresh[15239], Fresh[15238], Fresh[15237], Fresh[15236], Fresh[15235], Fresh[15234], Fresh[15233], Fresh[15232], Fresh[15231], Fresh[15230], Fresh[15229], Fresh[15228], Fresh[15227], Fresh[15226], Fresh[15225], Fresh[15224], Fresh[15223], Fresh[15222], Fresh[15221], Fresh[15220], Fresh[15219], Fresh[15218], Fresh[15217], Fresh[15216], Fresh[15215], Fresh[15214], Fresh[15213], Fresh[15212], Fresh[15211], Fresh[15210], Fresh[15209], Fresh[15208], Fresh[15207], Fresh[15206], Fresh[15205], Fresh[15204], Fresh[15203], Fresh[15202], Fresh[15201], Fresh[15200], Fresh[15199], Fresh[15198], Fresh[15197], Fresh[15196], Fresh[15195], Fresh[15194], Fresh[15193], Fresh[15192], Fresh[15191], Fresh[15190], Fresh[15189], Fresh[15188], Fresh[15187], Fresh[15186], Fresh[15185], Fresh[15184], Fresh[15183], Fresh[15182], Fresh[15181], Fresh[15180], Fresh[15179], Fresh[15178], Fresh[15177], Fresh[15176], Fresh[15175], Fresh[15174], Fresh[15173], Fresh[15172], Fresh[15171], Fresh[15170], Fresh[15169], Fresh[15168], Fresh[15167], Fresh[15166], Fresh[15165], Fresh[15164], Fresh[15163], Fresh[15162], Fresh[15161], Fresh[15160], Fresh[15159], Fresh[15158], Fresh[15157], Fresh[15156], Fresh[15155], Fresh[15154], Fresh[15153], Fresh[15152], Fresh[15151], Fresh[15150], Fresh[15149], Fresh[15148], Fresh[15147], Fresh[15146], Fresh[15145], Fresh[15144], Fresh[15143], Fresh[15142], Fresh[15141], Fresh[15140], Fresh[15139], Fresh[15138], Fresh[15137], Fresh[15136], Fresh[15135], Fresh[15134], Fresh[15133], Fresh[15132], Fresh[15131], Fresh[15130], Fresh[15129], Fresh[15128], Fresh[15127], Fresh[15126], Fresh[15125], Fresh[15124], Fresh[15123], Fresh[15122], Fresh[15121], Fresh[15120], Fresh[15119], Fresh[15118], Fresh[15117], Fresh[15116], Fresh[15115], Fresh[15114], Fresh[15113], Fresh[15112], Fresh[15111], Fresh[15110], Fresh[15109], Fresh[15108], Fresh[15107], Fresh[15106], Fresh[15105], Fresh[15104], Fresh[15103], Fresh[15102], Fresh[15101], Fresh[15100], Fresh[15099], Fresh[15098], Fresh[15097], Fresh[15096], Fresh[15095], Fresh[15094], Fresh[15093], Fresh[15092], Fresh[15091], Fresh[15090], Fresh[15089], Fresh[15088], Fresh[15087], Fresh[15086], Fresh[15085], Fresh[15084], Fresh[15083], Fresh[15082], Fresh[15081], Fresh[15080], Fresh[15079], Fresh[15078], Fresh[15077], Fresh[15076], Fresh[15075], Fresh[15074], Fresh[15073], Fresh[15072], Fresh[15071], Fresh[15070], Fresh[15069], Fresh[15068], Fresh[15067], Fresh[15066], Fresh[15065], Fresh[15064], Fresh[15063], Fresh[15062], Fresh[15061], Fresh[15060], Fresh[15059], Fresh[15058], Fresh[15057], Fresh[15056], Fresh[15055], Fresh[15054], Fresh[15053], Fresh[15052], Fresh[15051], Fresh[15050], Fresh[15049], Fresh[15048], Fresh[15047], Fresh[15046], Fresh[15045], Fresh[15044], Fresh[15043], Fresh[15042], Fresh[15041], Fresh[15040], Fresh[15039], Fresh[15038], Fresh[15037], Fresh[15036], Fresh[15035], Fresh[15034], Fresh[15033], Fresh[15032], Fresh[15031], Fresh[15030], Fresh[15029], Fresh[15028], Fresh[15027], Fresh[15026], Fresh[15025], Fresh[15024], Fresh[15023], Fresh[15022], Fresh[15021], Fresh[15020], Fresh[15019], Fresh[15018], Fresh[15017], Fresh[15016], Fresh[15015], Fresh[15014], Fresh[15013], Fresh[15012], Fresh[15011], Fresh[15010], Fresh[15009], Fresh[15008], Fresh[15007], Fresh[15006], Fresh[15005], Fresh[15004], Fresh[15003], Fresh[15002], Fresh[15001], Fresh[15000], Fresh[14999], Fresh[14998], Fresh[14997], Fresh[14996], Fresh[14995], Fresh[14994], Fresh[14993], Fresh[14992], Fresh[14991], Fresh[14990], Fresh[14989], Fresh[14988], Fresh[14987], Fresh[14986], Fresh[14985], Fresh[14984], Fresh[14983], Fresh[14982], Fresh[14981], Fresh[14980], Fresh[14979], Fresh[14978], Fresh[14977], Fresh[14976], Fresh[14975], Fresh[14974], Fresh[14973], Fresh[14972], Fresh[14971], Fresh[14970], Fresh[14969], Fresh[14968], Fresh[14967], Fresh[14966], Fresh[14965], Fresh[14964], Fresh[14963], Fresh[14962], Fresh[14961], Fresh[14960], Fresh[14959], Fresh[14958], Fresh[14957], Fresh[14956], Fresh[14955], Fresh[14954], Fresh[14953], Fresh[14952], Fresh[14951], Fresh[14950], Fresh[14949], Fresh[14948], Fresh[14947], Fresh[14946], Fresh[14945], Fresh[14944], Fresh[14943], Fresh[14942], Fresh[14941], Fresh[14940], Fresh[14939], Fresh[14938], Fresh[14937], Fresh[14936], Fresh[14935], Fresh[14934], Fresh[14933], Fresh[14932], Fresh[14931], Fresh[14930], Fresh[14929], Fresh[14928], Fresh[14927], Fresh[14926], Fresh[14925], Fresh[14924], Fresh[14923], Fresh[14922], Fresh[14921], Fresh[14920], Fresh[14919], Fresh[14918], Fresh[14917], Fresh[14916], Fresh[14915], Fresh[14914], Fresh[14913], Fresh[14912], Fresh[14911], Fresh[14910], Fresh[14909], Fresh[14908], Fresh[14907], Fresh[14906], Fresh[14905], Fresh[14904], Fresh[14903], Fresh[14902], Fresh[14901], Fresh[14900], Fresh[14899], Fresh[14898], Fresh[14897], Fresh[14896], Fresh[14895], Fresh[14894], Fresh[14893], Fresh[14892], Fresh[14891], Fresh[14890], Fresh[14889], Fresh[14888], Fresh[14887], Fresh[14886], Fresh[14885], Fresh[14884], Fresh[14883], Fresh[14882], Fresh[14881], Fresh[14880], Fresh[14879], Fresh[14878], Fresh[14877], Fresh[14876], Fresh[14875], Fresh[14874], Fresh[14873], Fresh[14872], Fresh[14871], Fresh[14870], Fresh[14869], Fresh[14868], Fresh[14867], Fresh[14866], Fresh[14865], Fresh[14864], Fresh[14863], Fresh[14862], Fresh[14861], Fresh[14860], Fresh[14859], Fresh[14858], Fresh[14857], Fresh[14856], Fresh[14855], Fresh[14854], Fresh[14853], Fresh[14852], Fresh[14851], Fresh[14850], Fresh[14849], Fresh[14848], Fresh[14847], Fresh[14846], Fresh[14845], Fresh[14844], Fresh[14843], Fresh[14842], Fresh[14841], Fresh[14840], Fresh[14839], Fresh[14838], Fresh[14837], Fresh[14836], Fresh[14835], Fresh[14834], Fresh[14833], Fresh[14832], Fresh[14831], Fresh[14830], Fresh[14829], Fresh[14828], Fresh[14827], Fresh[14826], Fresh[14825], Fresh[14824], Fresh[14823], Fresh[14822], Fresh[14821], Fresh[14820], Fresh[14819], Fresh[14818], Fresh[14817], Fresh[14816], Fresh[14815], Fresh[14814], Fresh[14813], Fresh[14812], Fresh[14811], Fresh[14810], Fresh[14809], Fresh[14808], Fresh[14807], Fresh[14806], Fresh[14805], Fresh[14804], Fresh[14803], Fresh[14802], Fresh[14801], Fresh[14800], Fresh[14799], Fresh[14798], Fresh[14797], Fresh[14796], Fresh[14795], Fresh[14794], Fresh[14793], Fresh[14792], Fresh[14791], Fresh[14790], Fresh[14789], Fresh[14788], Fresh[14787], Fresh[14786], Fresh[14785], Fresh[14784], Fresh[14783], Fresh[14782], Fresh[14781], Fresh[14780], Fresh[14779], Fresh[14778], Fresh[14777], Fresh[14776], Fresh[14775], Fresh[14774], Fresh[14773], Fresh[14772], Fresh[14771], Fresh[14770], Fresh[14769], Fresh[14768], Fresh[14767], Fresh[14766], Fresh[14765], Fresh[14764], Fresh[14763], Fresh[14762], Fresh[14761], Fresh[14760], Fresh[14759], Fresh[14758], Fresh[14757], Fresh[14756], Fresh[14755], Fresh[14754], Fresh[14753], Fresh[14752], Fresh[14751], Fresh[14750], Fresh[14749], Fresh[14748], Fresh[14747], Fresh[14746], Fresh[14745], Fresh[14744], Fresh[14743], Fresh[14742], Fresh[14741], Fresh[14740], Fresh[14739], Fresh[14738], Fresh[14737], Fresh[14736], Fresh[14735], Fresh[14734], Fresh[14733], Fresh[14732], Fresh[14731], Fresh[14730], Fresh[14729], Fresh[14728], Fresh[14727], Fresh[14726], Fresh[14725], Fresh[14724], Fresh[14723], Fresh[14722], Fresh[14721], Fresh[14720], Fresh[14719], Fresh[14718], Fresh[14717], Fresh[14716], Fresh[14715], Fresh[14714], Fresh[14713], Fresh[14712], Fresh[14711], Fresh[14710], Fresh[14709], Fresh[14708], Fresh[14707], Fresh[14706], Fresh[14705], Fresh[14704], Fresh[14703], Fresh[14702], Fresh[14701], Fresh[14700], Fresh[14699], Fresh[14698], Fresh[14697], Fresh[14696], Fresh[14695], Fresh[14694], Fresh[14693], Fresh[14692], Fresh[14691], Fresh[14690], Fresh[14689], Fresh[14688], Fresh[14687], Fresh[14686], Fresh[14685], Fresh[14684], Fresh[14683], Fresh[14682], Fresh[14681], Fresh[14680], Fresh[14679], Fresh[14678], Fresh[14677], Fresh[14676], Fresh[14675], Fresh[14674], Fresh[14673], Fresh[14672], Fresh[14671], Fresh[14670], Fresh[14669], Fresh[14668], Fresh[14667], Fresh[14666], Fresh[14665], Fresh[14664], Fresh[14663], Fresh[14662], Fresh[14661], Fresh[14660], Fresh[14659], Fresh[14658], Fresh[14657], Fresh[14656], Fresh[14655], Fresh[14654], Fresh[14653], Fresh[14652], Fresh[14651], Fresh[14650], Fresh[14649], Fresh[14648], Fresh[14647], Fresh[14646], Fresh[14645], Fresh[14644], Fresh[14643], Fresh[14642], Fresh[14641], Fresh[14640], Fresh[14639], Fresh[14638], Fresh[14637], Fresh[14636], Fresh[14635], Fresh[14634], Fresh[14633], Fresh[14632], Fresh[14631], Fresh[14630], Fresh[14629], Fresh[14628], Fresh[14627], Fresh[14626], Fresh[14625], Fresh[14624], Fresh[14623], Fresh[14622], Fresh[14621], Fresh[14620], Fresh[14619], Fresh[14618], Fresh[14617], Fresh[14616], Fresh[14615], Fresh[14614], Fresh[14613], Fresh[14612], Fresh[14611], Fresh[14610], Fresh[14609], Fresh[14608], Fresh[14607], Fresh[14606], Fresh[14605], Fresh[14604], Fresh[14603], Fresh[14602], Fresh[14601], Fresh[14600], Fresh[14599], Fresh[14598], Fresh[14597], Fresh[14596], Fresh[14595], Fresh[14594], Fresh[14593], Fresh[14592], Fresh[14591], Fresh[14590], Fresh[14589], Fresh[14588], Fresh[14587], Fresh[14586], Fresh[14585], Fresh[14584], Fresh[14583], Fresh[14582], Fresh[14581], Fresh[14580], Fresh[14579], Fresh[14578], Fresh[14577], Fresh[14576], Fresh[14575], Fresh[14574], Fresh[14573], Fresh[14572], Fresh[14571], Fresh[14570], Fresh[14569], Fresh[14568], Fresh[14567], Fresh[14566], Fresh[14565], Fresh[14564], Fresh[14563], Fresh[14562], Fresh[14561], Fresh[14560], Fresh[14559], Fresh[14558], Fresh[14557], Fresh[14556], Fresh[14555], Fresh[14554], Fresh[14553], Fresh[14552], Fresh[14551], Fresh[14550], Fresh[14549], Fresh[14548], Fresh[14547], Fresh[14546], Fresh[14545], Fresh[14544], Fresh[14543], Fresh[14542], Fresh[14541], Fresh[14540], Fresh[14539], Fresh[14538], Fresh[14537], Fresh[14536], Fresh[14535], Fresh[14534], Fresh[14533], Fresh[14532], Fresh[14531], Fresh[14530], Fresh[14529], Fresh[14528], Fresh[14527], Fresh[14526], Fresh[14525], Fresh[14524], Fresh[14523], Fresh[14522], Fresh[14521], Fresh[14520], Fresh[14519], Fresh[14518], Fresh[14517], Fresh[14516], Fresh[14515], Fresh[14514], Fresh[14513], Fresh[14512], Fresh[14511], Fresh[14510], Fresh[14509], Fresh[14508], Fresh[14507], Fresh[14506], Fresh[14505], Fresh[14504], Fresh[14503], Fresh[14502], Fresh[14501], Fresh[14500], Fresh[14499], Fresh[14498], Fresh[14497], Fresh[14496], Fresh[14495], Fresh[14494], Fresh[14493], Fresh[14492], Fresh[14491], Fresh[14490], Fresh[14489], Fresh[14488], Fresh[14487], Fresh[14486], Fresh[14485], Fresh[14484], Fresh[14483], Fresh[14482], Fresh[14481], Fresh[14480], Fresh[14479], Fresh[14478], Fresh[14477], Fresh[14476], Fresh[14475], Fresh[14474], Fresh[14473], Fresh[14472], Fresh[14471], Fresh[14470], Fresh[14469], Fresh[14468], Fresh[14467], Fresh[14466], Fresh[14465], Fresh[14464], Fresh[14463], Fresh[14462], Fresh[14461], Fresh[14460], Fresh[14459], Fresh[14458], Fresh[14457], Fresh[14456], Fresh[14455], Fresh[14454], Fresh[14453], Fresh[14452], Fresh[14451], Fresh[14450], Fresh[14449], Fresh[14448], Fresh[14447], Fresh[14446], Fresh[14445], Fresh[14444], Fresh[14443], Fresh[14442], Fresh[14441], Fresh[14440], Fresh[14439], Fresh[14438], Fresh[14437], Fresh[14436], Fresh[14435], Fresh[14434], Fresh[14433], Fresh[14432], Fresh[14431], Fresh[14430], Fresh[14429], Fresh[14428], Fresh[14427], Fresh[14426], Fresh[14425], Fresh[14424], Fresh[14423], Fresh[14422], Fresh[14421], Fresh[14420], Fresh[14419], Fresh[14418], Fresh[14417], Fresh[14416], Fresh[14415], Fresh[14414], Fresh[14413], Fresh[14412], Fresh[14411], Fresh[14410], Fresh[14409], Fresh[14408], Fresh[14407], Fresh[14406], Fresh[14405], Fresh[14404], Fresh[14403], Fresh[14402], Fresh[14401], Fresh[14400], Fresh[14399], Fresh[14398], Fresh[14397], Fresh[14396], Fresh[14395], Fresh[14394], Fresh[14393], Fresh[14392], Fresh[14391], Fresh[14390], Fresh[14389], Fresh[14388], Fresh[14387], Fresh[14386], Fresh[14385], Fresh[14384], Fresh[14383], Fresh[14382], Fresh[14381], Fresh[14380], Fresh[14379], Fresh[14378], Fresh[14377], Fresh[14376], Fresh[14375], Fresh[14374], Fresh[14373], Fresh[14372], Fresh[14371], Fresh[14370], Fresh[14369], Fresh[14368], Fresh[14367], Fresh[14366], Fresh[14365], Fresh[14364], Fresh[14363], Fresh[14362], Fresh[14361], Fresh[14360], Fresh[14359], Fresh[14358], Fresh[14357], Fresh[14356], Fresh[14355], Fresh[14354], Fresh[14353], Fresh[14352], Fresh[14351], Fresh[14350], Fresh[14349], Fresh[14348], Fresh[14347], Fresh[14346], Fresh[14345], Fresh[14344], Fresh[14343], Fresh[14342], Fresh[14341], Fresh[14340], Fresh[14339], Fresh[14338], Fresh[14337], Fresh[14336], Fresh[14335], Fresh[14334], Fresh[14333], Fresh[14332], Fresh[14331], Fresh[14330], Fresh[14329], Fresh[14328], Fresh[14327], Fresh[14326], Fresh[14325], Fresh[14324], Fresh[14323], Fresh[14322], Fresh[14321], Fresh[14320], Fresh[14319], Fresh[14318], Fresh[14317], Fresh[14316], Fresh[14315], Fresh[14314], Fresh[14313], Fresh[14312], Fresh[14311], Fresh[14310], Fresh[14309], Fresh[14308], Fresh[14307], Fresh[14306], Fresh[14305], Fresh[14304], Fresh[14303], Fresh[14302], Fresh[14301], Fresh[14300], Fresh[14299], Fresh[14298], Fresh[14297], Fresh[14296], Fresh[14295], Fresh[14294], Fresh[14293], Fresh[14292], Fresh[14291], Fresh[14290], Fresh[14289], Fresh[14288], Fresh[14287], Fresh[14286], Fresh[14285], Fresh[14284], Fresh[14283], Fresh[14282], Fresh[14281], Fresh[14280], Fresh[14279], Fresh[14278], Fresh[14277], Fresh[14276], Fresh[14275], Fresh[14274], Fresh[14273], Fresh[14272], Fresh[14271], Fresh[14270], Fresh[14269], Fresh[14268], Fresh[14267], Fresh[14266], Fresh[14265], Fresh[14264], Fresh[14263], Fresh[14262], Fresh[14261], Fresh[14260], Fresh[14259], Fresh[14258], Fresh[14257], Fresh[14256], Fresh[14255], Fresh[14254], Fresh[14253], Fresh[14252], Fresh[14251], Fresh[14250], Fresh[14249], Fresh[14248], Fresh[14247], Fresh[14246], Fresh[14245], Fresh[14244], Fresh[14243], Fresh[14242], Fresh[14241], Fresh[14240], Fresh[14239], Fresh[14238], Fresh[14237], Fresh[14236], Fresh[14235], Fresh[14234], Fresh[14233], Fresh[14232], Fresh[14231], Fresh[14230], Fresh[14229], Fresh[14228], Fresh[14227], Fresh[14226], Fresh[14225], Fresh[14224], Fresh[14223], Fresh[14222], Fresh[14221], Fresh[14220], Fresh[14219], Fresh[14218], Fresh[14217], Fresh[14216], Fresh[14215], Fresh[14214], Fresh[14213], Fresh[14212], Fresh[14211], Fresh[14210], Fresh[14209], Fresh[14208], Fresh[14207], Fresh[14206], Fresh[14205], Fresh[14204], Fresh[14203], Fresh[14202], Fresh[14201], Fresh[14200], Fresh[14199], Fresh[14198], Fresh[14197], Fresh[14196], Fresh[14195], Fresh[14194], Fresh[14193], Fresh[14192], Fresh[14191], Fresh[14190], Fresh[14189], Fresh[14188], Fresh[14187], Fresh[14186], Fresh[14185], Fresh[14184], Fresh[14183], Fresh[14182], Fresh[14181], Fresh[14180], Fresh[14179], Fresh[14178], Fresh[14177], Fresh[14176], Fresh[14175], Fresh[14174], Fresh[14173], Fresh[14172], Fresh[14171], Fresh[14170], Fresh[14169], Fresh[14168], Fresh[14167], Fresh[14166], Fresh[14165], Fresh[14164], Fresh[14163], Fresh[14162], Fresh[14161], Fresh[14160], Fresh[14159], Fresh[14158], Fresh[14157], Fresh[14156], Fresh[14155], Fresh[14154], Fresh[14153], Fresh[14152], Fresh[14151], Fresh[14150], Fresh[14149], Fresh[14148], Fresh[14147], Fresh[14146], Fresh[14145], Fresh[14144], Fresh[14143], Fresh[14142], Fresh[14141], Fresh[14140], Fresh[14139], Fresh[14138], Fresh[14137], Fresh[14136], Fresh[14135], Fresh[14134], Fresh[14133], Fresh[14132], Fresh[14131], Fresh[14130], Fresh[14129], Fresh[14128], Fresh[14127], Fresh[14126], Fresh[14125], Fresh[14124], Fresh[14123], Fresh[14122], Fresh[14121], Fresh[14120], Fresh[14119], Fresh[14118], Fresh[14117], Fresh[14116], Fresh[14115], Fresh[14114], Fresh[14113], Fresh[14112], Fresh[14111], Fresh[14110], Fresh[14109], Fresh[14108], Fresh[14107], Fresh[14106], Fresh[14105], Fresh[14104], Fresh[14103], Fresh[14102], Fresh[14101], Fresh[14100], Fresh[14099], Fresh[14098], Fresh[14097], Fresh[14096], Fresh[14095], Fresh[14094], Fresh[14093], Fresh[14092], Fresh[14091], Fresh[14090], Fresh[14089], Fresh[14088], Fresh[14087], Fresh[14086], Fresh[14085], Fresh[14084], Fresh[14083], Fresh[14082], Fresh[14081], Fresh[14080], Fresh[14079], Fresh[14078], Fresh[14077], Fresh[14076], Fresh[14075], Fresh[14074], Fresh[14073], Fresh[14072], Fresh[14071], Fresh[14070], Fresh[14069], Fresh[14068], Fresh[14067], Fresh[14066], Fresh[14065], Fresh[14064], Fresh[14063], Fresh[14062], Fresh[14061], Fresh[14060], Fresh[14059], Fresh[14058], Fresh[14057], Fresh[14056], Fresh[14055], Fresh[14054], Fresh[14053], Fresh[14052], Fresh[14051], Fresh[14050], Fresh[14049], Fresh[14048], Fresh[14047], Fresh[14046], Fresh[14045], Fresh[14044], Fresh[14043], Fresh[14042], Fresh[14041], Fresh[14040], Fresh[14039], Fresh[14038], Fresh[14037], Fresh[14036], Fresh[14035], Fresh[14034], Fresh[14033], Fresh[14032], Fresh[14031], Fresh[14030], Fresh[14029], Fresh[14028], Fresh[14027], Fresh[14026], Fresh[14025], Fresh[14024], Fresh[14023], Fresh[14022], Fresh[14021], Fresh[14020], Fresh[14019], Fresh[14018], Fresh[14017], Fresh[14016], Fresh[14015], Fresh[14014], Fresh[14013], Fresh[14012], Fresh[14011], Fresh[14010], Fresh[14009], Fresh[14008], Fresh[14007], Fresh[14006], Fresh[14005], Fresh[14004], Fresh[14003], Fresh[14002], Fresh[14001], Fresh[14000], Fresh[13999], Fresh[13998], Fresh[13997], Fresh[13996], Fresh[13995], Fresh[13994], Fresh[13993], Fresh[13992], Fresh[13991], Fresh[13990], Fresh[13989], Fresh[13988], Fresh[13987], Fresh[13986], Fresh[13985], Fresh[13984], Fresh[13983], Fresh[13982], Fresh[13981], Fresh[13980], Fresh[13979], Fresh[13978], Fresh[13977], Fresh[13976], Fresh[13975], Fresh[13974], Fresh[13973], Fresh[13972], Fresh[13971], Fresh[13970], Fresh[13969], Fresh[13968], Fresh[13967], Fresh[13966], Fresh[13965], Fresh[13964], Fresh[13963], Fresh[13962], Fresh[13961], Fresh[13960], Fresh[13959], Fresh[13958], Fresh[13957], Fresh[13956], Fresh[13955], Fresh[13954], Fresh[13953], Fresh[13952], Fresh[13951], Fresh[13950], Fresh[13949], Fresh[13948], Fresh[13947], Fresh[13946], Fresh[13945], Fresh[13944], Fresh[13943], Fresh[13942], Fresh[13941], Fresh[13940], Fresh[13939], Fresh[13938], Fresh[13937], Fresh[13936], Fresh[13935], Fresh[13934], Fresh[13933], Fresh[13932], Fresh[13931], Fresh[13930], Fresh[13929], Fresh[13928], Fresh[13927], Fresh[13926], Fresh[13925], Fresh[13924], Fresh[13923], Fresh[13922], Fresh[13921], Fresh[13920], Fresh[13919], Fresh[13918], Fresh[13917], Fresh[13916], Fresh[13915], Fresh[13914], Fresh[13913], Fresh[13912], Fresh[13911], Fresh[13910], Fresh[13909], Fresh[13908], Fresh[13907], Fresh[13906], Fresh[13905], Fresh[13904], Fresh[13903], Fresh[13902], Fresh[13901], Fresh[13900], Fresh[13899], Fresh[13898], Fresh[13897], Fresh[13896], Fresh[13895], Fresh[13894], Fresh[13893], Fresh[13892], Fresh[13891], Fresh[13890], Fresh[13889], Fresh[13888], Fresh[13887], Fresh[13886], Fresh[13885], Fresh[13884], Fresh[13883], Fresh[13882], Fresh[13881], Fresh[13880], Fresh[13879], Fresh[13878], Fresh[13877], Fresh[13876], Fresh[13875], Fresh[13874], Fresh[13873], Fresh[13872], Fresh[13871], Fresh[13870], Fresh[13869], Fresh[13868], Fresh[13867], Fresh[13866], Fresh[13865], Fresh[13864], Fresh[13863], Fresh[13862], Fresh[13861], Fresh[13860], Fresh[13859], Fresh[13858], Fresh[13857], Fresh[13856], Fresh[13855], Fresh[13854], Fresh[13853], Fresh[13852], Fresh[13851], Fresh[13850], Fresh[13849], Fresh[13848], Fresh[13847], Fresh[13846], Fresh[13845], Fresh[13844], Fresh[13843], Fresh[13842], Fresh[13841], Fresh[13840], Fresh[13839], Fresh[13838], Fresh[13837], Fresh[13836], Fresh[13835], Fresh[13834], Fresh[13833], Fresh[13832], Fresh[13831], Fresh[13830], Fresh[13829], Fresh[13828], Fresh[13827], Fresh[13826], Fresh[13825], Fresh[13824], Fresh[13823], Fresh[13822], Fresh[13821], Fresh[13820], Fresh[13819], Fresh[13818], Fresh[13817], Fresh[13816], Fresh[13815], Fresh[13814], Fresh[13813], Fresh[13812], Fresh[13811], Fresh[13810], Fresh[13809], Fresh[13808], Fresh[13807], Fresh[13806], Fresh[13805], Fresh[13804], Fresh[13803], Fresh[13802], Fresh[13801], Fresh[13800], Fresh[13799], Fresh[13798], Fresh[13797], Fresh[13796], Fresh[13795], Fresh[13794], Fresh[13793], Fresh[13792], Fresh[13791], Fresh[13790], Fresh[13789], Fresh[13788], Fresh[13787], Fresh[13786], Fresh[13785], Fresh[13784], Fresh[13783], Fresh[13782], Fresh[13781], Fresh[13780], Fresh[13779], Fresh[13778], Fresh[13777], Fresh[13776], Fresh[13775], Fresh[13774], Fresh[13773], Fresh[13772], Fresh[13771], Fresh[13770], Fresh[13769], Fresh[13768], Fresh[13767], Fresh[13766], Fresh[13765], Fresh[13764], Fresh[13763], Fresh[13762], Fresh[13761], Fresh[13760], Fresh[13759], Fresh[13758], Fresh[13757], Fresh[13756], Fresh[13755], Fresh[13754], Fresh[13753], Fresh[13752], Fresh[13751], Fresh[13750], Fresh[13749], Fresh[13748], Fresh[13747], Fresh[13746], Fresh[13745], Fresh[13744], Fresh[13743], Fresh[13742], Fresh[13741], Fresh[13740], Fresh[13739], Fresh[13738], Fresh[13737], Fresh[13736], Fresh[13735], Fresh[13734], Fresh[13733], Fresh[13732], Fresh[13731], Fresh[13730], Fresh[13729], Fresh[13728], Fresh[13727], Fresh[13726], Fresh[13725], Fresh[13724], Fresh[13723], Fresh[13722], Fresh[13721], Fresh[13720], Fresh[13719], Fresh[13718], Fresh[13717], Fresh[13716], Fresh[13715], Fresh[13714], Fresh[13713], Fresh[13712], Fresh[13711], Fresh[13710], Fresh[13709], Fresh[13708], Fresh[13707], Fresh[13706], Fresh[13705], Fresh[13704], Fresh[13703], Fresh[13702], Fresh[13701], Fresh[13700], Fresh[13699], Fresh[13698], Fresh[13697], Fresh[13696], Fresh[13695], Fresh[13694], Fresh[13693], Fresh[13692], Fresh[13691], Fresh[13690], Fresh[13689], Fresh[13688], Fresh[13687], Fresh[13686], Fresh[13685], Fresh[13684], Fresh[13683], Fresh[13682], Fresh[13681], Fresh[13680], Fresh[13679], Fresh[13678], Fresh[13677], Fresh[13676], Fresh[13675], Fresh[13674], Fresh[13673], Fresh[13672], Fresh[13671], Fresh[13670], Fresh[13669], Fresh[13668], Fresh[13667], Fresh[13666], Fresh[13665], Fresh[13664], Fresh[13663], Fresh[13662], Fresh[13661], Fresh[13660], Fresh[13659], Fresh[13658], Fresh[13657], Fresh[13656], Fresh[13655], Fresh[13654], Fresh[13653], Fresh[13652], Fresh[13651], Fresh[13650], Fresh[13649], Fresh[13648], Fresh[13647], Fresh[13646], Fresh[13645], Fresh[13644], Fresh[13643], Fresh[13642], Fresh[13641], Fresh[13640], Fresh[13639], Fresh[13638], Fresh[13637], Fresh[13636], Fresh[13635], Fresh[13634], Fresh[13633], Fresh[13632], Fresh[13631], Fresh[13630], Fresh[13629], Fresh[13628], Fresh[13627], Fresh[13626], Fresh[13625], Fresh[13624], Fresh[13623], Fresh[13622], Fresh[13621], Fresh[13620], Fresh[13619], Fresh[13618], Fresh[13617], Fresh[13616], Fresh[13615], Fresh[13614], Fresh[13613], Fresh[13612], Fresh[13611], Fresh[13610], Fresh[13609], Fresh[13608], Fresh[13607], Fresh[13606], Fresh[13605], Fresh[13604], Fresh[13603], Fresh[13602], Fresh[13601], Fresh[13600], Fresh[13599], Fresh[13598], Fresh[13597], Fresh[13596], Fresh[13595], Fresh[13594], Fresh[13593], Fresh[13592], Fresh[13591], Fresh[13590], Fresh[13589], Fresh[13588], Fresh[13587], Fresh[13586], Fresh[13585], Fresh[13584], Fresh[13583], Fresh[13582], Fresh[13581], Fresh[13580], Fresh[13579], Fresh[13578], Fresh[13577], Fresh[13576], Fresh[13575], Fresh[13574], Fresh[13573], Fresh[13572], Fresh[13571], Fresh[13570], Fresh[13569], Fresh[13568], Fresh[13567], Fresh[13566], Fresh[13565], Fresh[13564], Fresh[13563], Fresh[13562], Fresh[13561], Fresh[13560], Fresh[13559], Fresh[13558], Fresh[13557], Fresh[13556], Fresh[13555], Fresh[13554], Fresh[13553], Fresh[13552], Fresh[13551], Fresh[13550], Fresh[13549], Fresh[13548], Fresh[13547], Fresh[13546], Fresh[13545], Fresh[13544], Fresh[13543], Fresh[13542], Fresh[13541], Fresh[13540], Fresh[13539], Fresh[13538], Fresh[13537], Fresh[13536], Fresh[13535], Fresh[13534], Fresh[13533], Fresh[13532], Fresh[13531], Fresh[13530], Fresh[13529], Fresh[13528], Fresh[13527], Fresh[13526], Fresh[13525], Fresh[13524], Fresh[13523], Fresh[13522], Fresh[13521], Fresh[13520], Fresh[13519], Fresh[13518], Fresh[13517], Fresh[13516], Fresh[13515], Fresh[13514], Fresh[13513], Fresh[13512], Fresh[13511], Fresh[13510], Fresh[13509], Fresh[13508], Fresh[13507], Fresh[13506], Fresh[13505], Fresh[13504], Fresh[13503], Fresh[13502], Fresh[13501], Fresh[13500], Fresh[13499], Fresh[13498], Fresh[13497], Fresh[13496], Fresh[13495], Fresh[13494], Fresh[13493], Fresh[13492], Fresh[13491], Fresh[13490], Fresh[13489], Fresh[13488], Fresh[13487], Fresh[13486], Fresh[13485], Fresh[13484], Fresh[13483], Fresh[13482], Fresh[13481], Fresh[13480], Fresh[13479], Fresh[13478], Fresh[13477], Fresh[13476], Fresh[13475], Fresh[13474], Fresh[13473], Fresh[13472], Fresh[13471], Fresh[13470], Fresh[13469], Fresh[13468], Fresh[13467], Fresh[13466], Fresh[13465], Fresh[13464], Fresh[13463], Fresh[13462], Fresh[13461], Fresh[13460], Fresh[13459], Fresh[13458], Fresh[13457], Fresh[13456], Fresh[13455], Fresh[13454], Fresh[13453], Fresh[13452], Fresh[13451], Fresh[13450], Fresh[13449], Fresh[13448], Fresh[13447], Fresh[13446], Fresh[13445], Fresh[13444], Fresh[13443], Fresh[13442], Fresh[13441], Fresh[13440], Fresh[13439], Fresh[13438], Fresh[13437], Fresh[13436], Fresh[13435], Fresh[13434], Fresh[13433], Fresh[13432], Fresh[13431], Fresh[13430], Fresh[13429], Fresh[13428], Fresh[13427], Fresh[13426], Fresh[13425], Fresh[13424], Fresh[13423], Fresh[13422], Fresh[13421], Fresh[13420], Fresh[13419], Fresh[13418], Fresh[13417], Fresh[13416], Fresh[13415], Fresh[13414], Fresh[13413], Fresh[13412], Fresh[13411], Fresh[13410], Fresh[13409], Fresh[13408], Fresh[13407], Fresh[13406], Fresh[13405], Fresh[13404], Fresh[13403], Fresh[13402], Fresh[13401], Fresh[13400], Fresh[13399], Fresh[13398], Fresh[13397], Fresh[13396], Fresh[13395], Fresh[13394], Fresh[13393], Fresh[13392], Fresh[13391], Fresh[13390], Fresh[13389], Fresh[13388], Fresh[13387], Fresh[13386], Fresh[13385], Fresh[13384], Fresh[13383], Fresh[13382], Fresh[13381], Fresh[13380], Fresh[13379], Fresh[13378], Fresh[13377], Fresh[13376], Fresh[13375], Fresh[13374], Fresh[13373], Fresh[13372], Fresh[13371], Fresh[13370], Fresh[13369], Fresh[13368], Fresh[13367], Fresh[13366], Fresh[13365], Fresh[13364], Fresh[13363], Fresh[13362], Fresh[13361], Fresh[13360], Fresh[13359], Fresh[13358], Fresh[13357], Fresh[13356], Fresh[13355], Fresh[13354], Fresh[13353], Fresh[13352], Fresh[13351], Fresh[13350], Fresh[13349], Fresh[13348], Fresh[13347], Fresh[13346], Fresh[13345], Fresh[13344], Fresh[13343], Fresh[13342], Fresh[13341], Fresh[13340], Fresh[13339], Fresh[13338], Fresh[13337], Fresh[13336], Fresh[13335], Fresh[13334], Fresh[13333], Fresh[13332], Fresh[13331], Fresh[13330], Fresh[13329], Fresh[13328], Fresh[13327], Fresh[13326], Fresh[13325], Fresh[13324], Fresh[13323], Fresh[13322], Fresh[13321], Fresh[13320], Fresh[13319], Fresh[13318], Fresh[13317], Fresh[13316], Fresh[13315], Fresh[13314], Fresh[13313], Fresh[13312], Fresh[13311], Fresh[13310], Fresh[13309], Fresh[13308], Fresh[13307], Fresh[13306], Fresh[13305], Fresh[13304], Fresh[13303], Fresh[13302], Fresh[13301], Fresh[13300], Fresh[13299], Fresh[13298], Fresh[13297], Fresh[13296], Fresh[13295], Fresh[13294], Fresh[13293], Fresh[13292], Fresh[13291], Fresh[13290], Fresh[13289], Fresh[13288], Fresh[13287], Fresh[13286], Fresh[13285], Fresh[13284], Fresh[13283], Fresh[13282], Fresh[13281], Fresh[13280], Fresh[13279], Fresh[13278], Fresh[13277], Fresh[13276], Fresh[13275], Fresh[13274], Fresh[13273], Fresh[13272], Fresh[13271], Fresh[13270], Fresh[13269], Fresh[13268], Fresh[13267], Fresh[13266], Fresh[13265], Fresh[13264], Fresh[13263], Fresh[13262], Fresh[13261], Fresh[13260], Fresh[13259], Fresh[13258], Fresh[13257], Fresh[13256], Fresh[13255], Fresh[13254], Fresh[13253], Fresh[13252], Fresh[13251], Fresh[13250], Fresh[13249], Fresh[13248], Fresh[13247], Fresh[13246], Fresh[13245], Fresh[13244], Fresh[13243], Fresh[13242], Fresh[13241], Fresh[13240], Fresh[13239], Fresh[13238], Fresh[13237], Fresh[13236], Fresh[13235], Fresh[13234], Fresh[13233], Fresh[13232], Fresh[13231], Fresh[13230], Fresh[13229], Fresh[13228], Fresh[13227], Fresh[13226], Fresh[13225], Fresh[13224], Fresh[13223], Fresh[13222], Fresh[13221], Fresh[13220], Fresh[13219], Fresh[13218], Fresh[13217], Fresh[13216], Fresh[13215], Fresh[13214], Fresh[13213], Fresh[13212], Fresh[13211], Fresh[13210], Fresh[13209], Fresh[13208], Fresh[13207], Fresh[13206], Fresh[13205], Fresh[13204], Fresh[13203], Fresh[13202], Fresh[13201], Fresh[13200], Fresh[13199], Fresh[13198], Fresh[13197], Fresh[13196], Fresh[13195], Fresh[13194], Fresh[13193], Fresh[13192], Fresh[13191], Fresh[13190], Fresh[13189], Fresh[13188], Fresh[13187], Fresh[13186], Fresh[13185], Fresh[13184], Fresh[13183], Fresh[13182], Fresh[13181], Fresh[13180], Fresh[13179], Fresh[13178], Fresh[13177], Fresh[13176], Fresh[13175], Fresh[13174], Fresh[13173], Fresh[13172], Fresh[13171], Fresh[13170], Fresh[13169], Fresh[13168], Fresh[13167], Fresh[13166], Fresh[13165], Fresh[13164], Fresh[13163], Fresh[13162], Fresh[13161], Fresh[13160], Fresh[13159], Fresh[13158], Fresh[13157], Fresh[13156], Fresh[13155], Fresh[13154], Fresh[13153], Fresh[13152], Fresh[13151], Fresh[13150], Fresh[13149], Fresh[13148], Fresh[13147], Fresh[13146], Fresh[13145], Fresh[13144], Fresh[13143], Fresh[13142], Fresh[13141], Fresh[13140], Fresh[13139], Fresh[13138], Fresh[13137], Fresh[13136], Fresh[13135], Fresh[13134], Fresh[13133], Fresh[13132], Fresh[13131], Fresh[13130], Fresh[13129], Fresh[13128], Fresh[13127], Fresh[13126], Fresh[13125], Fresh[13124], Fresh[13123], Fresh[13122], Fresh[13121], Fresh[13120], Fresh[13119], Fresh[13118], Fresh[13117], Fresh[13116], Fresh[13115], Fresh[13114], Fresh[13113], Fresh[13112], Fresh[13111], Fresh[13110], Fresh[13109], Fresh[13108], Fresh[13107], Fresh[13106], Fresh[13105], Fresh[13104], Fresh[13103], Fresh[13102], Fresh[13101], Fresh[13100], Fresh[13099], Fresh[13098], Fresh[13097], Fresh[13096], Fresh[13095], Fresh[13094], Fresh[13093], Fresh[13092], Fresh[13091], Fresh[13090], Fresh[13089], Fresh[13088], Fresh[13087], Fresh[13086], Fresh[13085], Fresh[13084], Fresh[13083], Fresh[13082], Fresh[13081], Fresh[13080], Fresh[13079], Fresh[13078], Fresh[13077], Fresh[13076], Fresh[13075], Fresh[13074], Fresh[13073], Fresh[13072], Fresh[13071], Fresh[13070], Fresh[13069], Fresh[13068], Fresh[13067], Fresh[13066], Fresh[13065], Fresh[13064], Fresh[13063], Fresh[13062], Fresh[13061], Fresh[13060], Fresh[13059], Fresh[13058], Fresh[13057], Fresh[13056], Fresh[13055], Fresh[13054], Fresh[13053], Fresh[13052], Fresh[13051], Fresh[13050], Fresh[13049], Fresh[13048], Fresh[13047], Fresh[13046], Fresh[13045], Fresh[13044], Fresh[13043], Fresh[13042], Fresh[13041], Fresh[13040], Fresh[13039], Fresh[13038], Fresh[13037], Fresh[13036], Fresh[13035], Fresh[13034], Fresh[13033], Fresh[13032], Fresh[13031], Fresh[13030], Fresh[13029], Fresh[13028], Fresh[13027], Fresh[13026], Fresh[13025], Fresh[13024], Fresh[13023], Fresh[13022], Fresh[13021], Fresh[13020], Fresh[13019], Fresh[13018], Fresh[13017], Fresh[13016], Fresh[13015], Fresh[13014], Fresh[13013], Fresh[13012], Fresh[13011], Fresh[13010], Fresh[13009], Fresh[13008], Fresh[13007], Fresh[13006], Fresh[13005], Fresh[13004], Fresh[13003], Fresh[13002], Fresh[13001], Fresh[13000], Fresh[12999], Fresh[12998], Fresh[12997], Fresh[12996], Fresh[12995], Fresh[12994], Fresh[12993], Fresh[12992], Fresh[12991], Fresh[12990], Fresh[12989], Fresh[12988], Fresh[12987], Fresh[12986], Fresh[12985], Fresh[12984], Fresh[12983], Fresh[12982], Fresh[12981], Fresh[12980], Fresh[12979], Fresh[12978], Fresh[12977], Fresh[12976], Fresh[12975], Fresh[12974], Fresh[12973], Fresh[12972], Fresh[12971], Fresh[12970], Fresh[12969], Fresh[12968], Fresh[12967], Fresh[12966], Fresh[12965], Fresh[12964], Fresh[12963], Fresh[12962], Fresh[12961], Fresh[12960], Fresh[12959], Fresh[12958], Fresh[12957], Fresh[12956], Fresh[12955], Fresh[12954], Fresh[12953], Fresh[12952], Fresh[12951], Fresh[12950], Fresh[12949], Fresh[12948], Fresh[12947], Fresh[12946], Fresh[12945], Fresh[12944], Fresh[12943], Fresh[12942], Fresh[12941], Fresh[12940], Fresh[12939], Fresh[12938], Fresh[12937], Fresh[12936], Fresh[12935], Fresh[12934], Fresh[12933], Fresh[12932], Fresh[12931], Fresh[12930], Fresh[12929], Fresh[12928], Fresh[12927], Fresh[12926], Fresh[12925], Fresh[12924], Fresh[12923], Fresh[12922], Fresh[12921], Fresh[12920], Fresh[12919], Fresh[12918], Fresh[12917], Fresh[12916], Fresh[12915], Fresh[12914], Fresh[12913], Fresh[12912], Fresh[12911], Fresh[12910], Fresh[12909], Fresh[12908], Fresh[12907], Fresh[12906], Fresh[12905], Fresh[12904], Fresh[12903], Fresh[12902], Fresh[12901], Fresh[12900], Fresh[12899], Fresh[12898], Fresh[12897], Fresh[12896], Fresh[12895], Fresh[12894], Fresh[12893], Fresh[12892], Fresh[12891], Fresh[12890], Fresh[12889], Fresh[12888], Fresh[12887], Fresh[12886], Fresh[12885], Fresh[12884], Fresh[12883], Fresh[12882], Fresh[12881], Fresh[12880], Fresh[12879], Fresh[12878], Fresh[12877], Fresh[12876], Fresh[12875], Fresh[12874], Fresh[12873], Fresh[12872], Fresh[12871], Fresh[12870], Fresh[12869], Fresh[12868], Fresh[12867], Fresh[12866], Fresh[12865], Fresh[12864], Fresh[12863], Fresh[12862], Fresh[12861], Fresh[12860], Fresh[12859], Fresh[12858], Fresh[12857], Fresh[12856], Fresh[12855], Fresh[12854], Fresh[12853], Fresh[12852], Fresh[12851], Fresh[12850], Fresh[12849], Fresh[12848], Fresh[12847], Fresh[12846], Fresh[12845], Fresh[12844], Fresh[12843], Fresh[12842], Fresh[12841], Fresh[12840], Fresh[12839], Fresh[12838], Fresh[12837], Fresh[12836], Fresh[12835], Fresh[12834], Fresh[12833], Fresh[12832], Fresh[12831], Fresh[12830], Fresh[12829], Fresh[12828], Fresh[12827], Fresh[12826], Fresh[12825], Fresh[12824], Fresh[12823], Fresh[12822], Fresh[12821], Fresh[12820], Fresh[12819], Fresh[12818], Fresh[12817], Fresh[12816], Fresh[12815], Fresh[12814], Fresh[12813], Fresh[12812], Fresh[12811], Fresh[12810], Fresh[12809], Fresh[12808], Fresh[12807], Fresh[12806], Fresh[12805], Fresh[12804], Fresh[12803], Fresh[12802], Fresh[12801], Fresh[12800], Fresh[12799], Fresh[12798], Fresh[12797], Fresh[12796], Fresh[12795], Fresh[12794], Fresh[12793], Fresh[12792], Fresh[12791], Fresh[12790], Fresh[12789], Fresh[12788], Fresh[12787], Fresh[12786], Fresh[12785], Fresh[12784], Fresh[12783], Fresh[12782], Fresh[12781], Fresh[12780], Fresh[12779], Fresh[12778], Fresh[12777], Fresh[12776], Fresh[12775], Fresh[12774], Fresh[12773], Fresh[12772], Fresh[12771], Fresh[12770], Fresh[12769], Fresh[12768], Fresh[12767], Fresh[12766], Fresh[12765], Fresh[12764], Fresh[12763], Fresh[12762], Fresh[12761], Fresh[12760], Fresh[12759], Fresh[12758], Fresh[12757], Fresh[12756], Fresh[12755], Fresh[12754], Fresh[12753], Fresh[12752], Fresh[12751], Fresh[12750], Fresh[12749], Fresh[12748], Fresh[12747], Fresh[12746], Fresh[12745], Fresh[12744], Fresh[12743], Fresh[12742], Fresh[12741], Fresh[12740], Fresh[12739], Fresh[12738], Fresh[12737], Fresh[12736], Fresh[12735], Fresh[12734], Fresh[12733], Fresh[12732], Fresh[12731], Fresh[12730], Fresh[12729], Fresh[12728], Fresh[12727], Fresh[12726], Fresh[12725], Fresh[12724], Fresh[12723], Fresh[12722], Fresh[12721], Fresh[12720], Fresh[12719], Fresh[12718], Fresh[12717], Fresh[12716], Fresh[12715], Fresh[12714], Fresh[12713], Fresh[12712], Fresh[12711], Fresh[12710], Fresh[12709], Fresh[12708], Fresh[12707], Fresh[12706], Fresh[12705], Fresh[12704], Fresh[12703], Fresh[12702], Fresh[12701], Fresh[12700], Fresh[12699], Fresh[12698], Fresh[12697], Fresh[12696], Fresh[12695], Fresh[12694], Fresh[12693], Fresh[12692], Fresh[12691], Fresh[12690], Fresh[12689], Fresh[12688], Fresh[12687], Fresh[12686], Fresh[12685], Fresh[12684], Fresh[12683], Fresh[12682], Fresh[12681], Fresh[12680], Fresh[12679], Fresh[12678], Fresh[12677], Fresh[12676], Fresh[12675], Fresh[12674], Fresh[12673], Fresh[12672], Fresh[12671], Fresh[12670], Fresh[12669], Fresh[12668], Fresh[12667], Fresh[12666], Fresh[12665], Fresh[12664], Fresh[12663], Fresh[12662], Fresh[12661], Fresh[12660], Fresh[12659], Fresh[12658], Fresh[12657], Fresh[12656], Fresh[12655], Fresh[12654], Fresh[12653], Fresh[12652], Fresh[12651], Fresh[12650], Fresh[12649], Fresh[12648], Fresh[12647], Fresh[12646], Fresh[12645], Fresh[12644], Fresh[12643], Fresh[12642], Fresh[12641], Fresh[12640], Fresh[12639], Fresh[12638], Fresh[12637], Fresh[12636], Fresh[12635], Fresh[12634], Fresh[12633], Fresh[12632], Fresh[12631], Fresh[12630], Fresh[12629], Fresh[12628], Fresh[12627], Fresh[12626], Fresh[12625], Fresh[12624], Fresh[12623], Fresh[12622], Fresh[12621], Fresh[12620], Fresh[12619], Fresh[12618], Fresh[12617], Fresh[12616], Fresh[12615], Fresh[12614], Fresh[12613], Fresh[12612], Fresh[12611], Fresh[12610], Fresh[12609], Fresh[12608], Fresh[12607], Fresh[12606], Fresh[12605], Fresh[12604], Fresh[12603], Fresh[12602], Fresh[12601], Fresh[12600], Fresh[12599], Fresh[12598], Fresh[12597], Fresh[12596], Fresh[12595], Fresh[12594], Fresh[12593], Fresh[12592], Fresh[12591], Fresh[12590], Fresh[12589], Fresh[12588], Fresh[12587], Fresh[12586], Fresh[12585], Fresh[12584], Fresh[12583], Fresh[12582], Fresh[12581], Fresh[12580], Fresh[12579], Fresh[12578], Fresh[12577], Fresh[12576], Fresh[12575], Fresh[12574], Fresh[12573], Fresh[12572], Fresh[12571], Fresh[12570], Fresh[12569], Fresh[12568], Fresh[12567], Fresh[12566], Fresh[12565], Fresh[12564], Fresh[12563], Fresh[12562], Fresh[12561], Fresh[12560], Fresh[12559], Fresh[12558], Fresh[12557], Fresh[12556], Fresh[12555], Fresh[12554], Fresh[12553], Fresh[12552], Fresh[12551], Fresh[12550], Fresh[12549], Fresh[12548], Fresh[12547], Fresh[12546], Fresh[12545], Fresh[12544], Fresh[12543], Fresh[12542], Fresh[12541], Fresh[12540], Fresh[12539], Fresh[12538], Fresh[12537], Fresh[12536], Fresh[12535], Fresh[12534], Fresh[12533], Fresh[12532], Fresh[12531], Fresh[12530], Fresh[12529], Fresh[12528], Fresh[12527], Fresh[12526], Fresh[12525], Fresh[12524], Fresh[12523], Fresh[12522], Fresh[12521], Fresh[12520], Fresh[12519], Fresh[12518], Fresh[12517], Fresh[12516], Fresh[12515], Fresh[12514], Fresh[12513], Fresh[12512], Fresh[12511], Fresh[12510], Fresh[12509], Fresh[12508], Fresh[12507], Fresh[12506], Fresh[12505], Fresh[12504], Fresh[12503], Fresh[12502], Fresh[12501], Fresh[12500], Fresh[12499], Fresh[12498], Fresh[12497], Fresh[12496], Fresh[12495], Fresh[12494], Fresh[12493], Fresh[12492], Fresh[12491], Fresh[12490], Fresh[12489], Fresh[12488], Fresh[12487], Fresh[12486], Fresh[12485], Fresh[12484], Fresh[12483], Fresh[12482], Fresh[12481], Fresh[12480], Fresh[12479], Fresh[12478], Fresh[12477], Fresh[12476], Fresh[12475], Fresh[12474], Fresh[12473], Fresh[12472], Fresh[12471], Fresh[12470], Fresh[12469], Fresh[12468], Fresh[12467], Fresh[12466], Fresh[12465], Fresh[12464], Fresh[12463], Fresh[12462], Fresh[12461], Fresh[12460], Fresh[12459], Fresh[12458], Fresh[12457], Fresh[12456], Fresh[12455], Fresh[12454], Fresh[12453], Fresh[12452], Fresh[12451], Fresh[12450], Fresh[12449], Fresh[12448], Fresh[12447], Fresh[12446], Fresh[12445], Fresh[12444], Fresh[12443], Fresh[12442], Fresh[12441], Fresh[12440], Fresh[12439], Fresh[12438], Fresh[12437], Fresh[12436], Fresh[12435], Fresh[12434], Fresh[12433], Fresh[12432], Fresh[12431], Fresh[12430], Fresh[12429], Fresh[12428], Fresh[12427], Fresh[12426], Fresh[12425], Fresh[12424], Fresh[12423], Fresh[12422], Fresh[12421], Fresh[12420], Fresh[12419], Fresh[12418], Fresh[12417], Fresh[12416], Fresh[12415], Fresh[12414], Fresh[12413], Fresh[12412], Fresh[12411], Fresh[12410], Fresh[12409], Fresh[12408], Fresh[12407], Fresh[12406], Fresh[12405], Fresh[12404], Fresh[12403], Fresh[12402], Fresh[12401], Fresh[12400], Fresh[12399], Fresh[12398], Fresh[12397], Fresh[12396], Fresh[12395], Fresh[12394], Fresh[12393], Fresh[12392], Fresh[12391], Fresh[12390], Fresh[12389], Fresh[12388], Fresh[12387], Fresh[12386], Fresh[12385], Fresh[12384], Fresh[12383], Fresh[12382], Fresh[12381], Fresh[12380], Fresh[12379], Fresh[12378], Fresh[12377], Fresh[12376], Fresh[12375], Fresh[12374], Fresh[12373], Fresh[12372], Fresh[12371], Fresh[12370], Fresh[12369], Fresh[12368], Fresh[12367], Fresh[12366], Fresh[12365], Fresh[12364], Fresh[12363], Fresh[12362], Fresh[12361], Fresh[12360], Fresh[12359], Fresh[12358], Fresh[12357], Fresh[12356], Fresh[12355], Fresh[12354], Fresh[12353], Fresh[12352], Fresh[12351], Fresh[12350], Fresh[12349], Fresh[12348], Fresh[12347], Fresh[12346], Fresh[12345], Fresh[12344], Fresh[12343], Fresh[12342], Fresh[12341], Fresh[12340], Fresh[12339], Fresh[12338], Fresh[12337], Fresh[12336], Fresh[12335], Fresh[12334], Fresh[12333], Fresh[12332], Fresh[12331], Fresh[12330], Fresh[12329], Fresh[12328], Fresh[12327], Fresh[12326], Fresh[12325], Fresh[12324], Fresh[12323], Fresh[12322], Fresh[12321], Fresh[12320], Fresh[12319], Fresh[12318], Fresh[12317], Fresh[12316], Fresh[12315], Fresh[12314], Fresh[12313], Fresh[12312], Fresh[12311], Fresh[12310], Fresh[12309], Fresh[12308], Fresh[12307], Fresh[12306], Fresh[12305], Fresh[12304], Fresh[12303], Fresh[12302], Fresh[12301], Fresh[12300], Fresh[12299], Fresh[12298], Fresh[12297], Fresh[12296], Fresh[12295], Fresh[12294], Fresh[12293], Fresh[12292], Fresh[12291], Fresh[12290], Fresh[12289], Fresh[12288], Fresh[12287], Fresh[12286], Fresh[12285], Fresh[12284], Fresh[12283], Fresh[12282], Fresh[12281], Fresh[12280], Fresh[12279], Fresh[12278], Fresh[12277], Fresh[12276], Fresh[12275], Fresh[12274], Fresh[12273], Fresh[12272], Fresh[12271], Fresh[12270], Fresh[12269], Fresh[12268], Fresh[12267], Fresh[12266], Fresh[12265], Fresh[12264], Fresh[12263], Fresh[12262], Fresh[12261], Fresh[12260], Fresh[12259], Fresh[12258], Fresh[12257], Fresh[12256], Fresh[12255], Fresh[12254], Fresh[12253], Fresh[12252], Fresh[12251], Fresh[12250], Fresh[12249], Fresh[12248], Fresh[12247], Fresh[12246], Fresh[12245], Fresh[12244], Fresh[12243], Fresh[12242], Fresh[12241], Fresh[12240], Fresh[12239], Fresh[12238], Fresh[12237], Fresh[12236], Fresh[12235], Fresh[12234], Fresh[12233], Fresh[12232], Fresh[12231], Fresh[12230], Fresh[12229], Fresh[12228], Fresh[12227], Fresh[12226], Fresh[12225], Fresh[12224], Fresh[12223], Fresh[12222], Fresh[12221], Fresh[12220], Fresh[12219], Fresh[12218], Fresh[12217], Fresh[12216], Fresh[12215], Fresh[12214], Fresh[12213], Fresh[12212], Fresh[12211], Fresh[12210], Fresh[12209], Fresh[12208], Fresh[12207], Fresh[12206], Fresh[12205], Fresh[12204], Fresh[12203], Fresh[12202], Fresh[12201], Fresh[12200], Fresh[12199], Fresh[12198], Fresh[12197], Fresh[12196], Fresh[12195], Fresh[12194], Fresh[12193], Fresh[12192], Fresh[12191], Fresh[12190], Fresh[12189], Fresh[12188], Fresh[12187], Fresh[12186], Fresh[12185], Fresh[12184], Fresh[12183], Fresh[12182], Fresh[12181], Fresh[12180], Fresh[12179], Fresh[12178], Fresh[12177], Fresh[12176], Fresh[12175], Fresh[12174], Fresh[12173], Fresh[12172], Fresh[12171], Fresh[12170], Fresh[12169], Fresh[12168], Fresh[12167], Fresh[12166], Fresh[12165], Fresh[12164], Fresh[12163], Fresh[12162], Fresh[12161], Fresh[12160], Fresh[12159], Fresh[12158], Fresh[12157], Fresh[12156], Fresh[12155], Fresh[12154], Fresh[12153], Fresh[12152], Fresh[12151], Fresh[12150], Fresh[12149], Fresh[12148], Fresh[12147], Fresh[12146], Fresh[12145], Fresh[12144], Fresh[12143], Fresh[12142], Fresh[12141], Fresh[12140], Fresh[12139], Fresh[12138], Fresh[12137], Fresh[12136], Fresh[12135], Fresh[12134], Fresh[12133], Fresh[12132], Fresh[12131], Fresh[12130], Fresh[12129], Fresh[12128], Fresh[12127], Fresh[12126], Fresh[12125], Fresh[12124], Fresh[12123], Fresh[12122], Fresh[12121], Fresh[12120], Fresh[12119], Fresh[12118], Fresh[12117], Fresh[12116], Fresh[12115], Fresh[12114], Fresh[12113], Fresh[12112], Fresh[12111], Fresh[12110], Fresh[12109], Fresh[12108], Fresh[12107], Fresh[12106], Fresh[12105], Fresh[12104], Fresh[12103], Fresh[12102], Fresh[12101], Fresh[12100], Fresh[12099], Fresh[12098], Fresh[12097], Fresh[12096], Fresh[12095], Fresh[12094], Fresh[12093], Fresh[12092], Fresh[12091], Fresh[12090], Fresh[12089], Fresh[12088], Fresh[12087], Fresh[12086], Fresh[12085], Fresh[12084], Fresh[12083], Fresh[12082], Fresh[12081], Fresh[12080], Fresh[12079], Fresh[12078], Fresh[12077], Fresh[12076], Fresh[12075], Fresh[12074], Fresh[12073], Fresh[12072], Fresh[12071], Fresh[12070], Fresh[12069], Fresh[12068], Fresh[12067], Fresh[12066], Fresh[12065], Fresh[12064], Fresh[12063], Fresh[12062], Fresh[12061], Fresh[12060], Fresh[12059], Fresh[12058], Fresh[12057], Fresh[12056], Fresh[12055], Fresh[12054], Fresh[12053], Fresh[12052], Fresh[12051], Fresh[12050], Fresh[12049], Fresh[12048], Fresh[12047], Fresh[12046], Fresh[12045], Fresh[12044], Fresh[12043], Fresh[12042], Fresh[12041], Fresh[12040], Fresh[12039], Fresh[12038], Fresh[12037], Fresh[12036], Fresh[12035], Fresh[12034], Fresh[12033], Fresh[12032], Fresh[12031], Fresh[12030], Fresh[12029], Fresh[12028], Fresh[12027], Fresh[12026], Fresh[12025], Fresh[12024], Fresh[12023], Fresh[12022], Fresh[12021], Fresh[12020], Fresh[12019], Fresh[12018], Fresh[12017], Fresh[12016], Fresh[12015], Fresh[12014], Fresh[12013], Fresh[12012], Fresh[12011], Fresh[12010], Fresh[12009], Fresh[12008], Fresh[12007], Fresh[12006], Fresh[12005], Fresh[12004], Fresh[12003], Fresh[12002], Fresh[12001], Fresh[12000], Fresh[11999], Fresh[11998], Fresh[11997], Fresh[11996], Fresh[11995], Fresh[11994], Fresh[11993], Fresh[11992], Fresh[11991], Fresh[11990], Fresh[11989], Fresh[11988], Fresh[11987], Fresh[11986], Fresh[11985], Fresh[11984], Fresh[11983], Fresh[11982], Fresh[11981], Fresh[11980], Fresh[11979], Fresh[11978], Fresh[11977], Fresh[11976], Fresh[11975], Fresh[11974], Fresh[11973], Fresh[11972], Fresh[11971], Fresh[11970], Fresh[11969], Fresh[11968], Fresh[11967], Fresh[11966], Fresh[11965], Fresh[11964], Fresh[11963], Fresh[11962], Fresh[11961], Fresh[11960], Fresh[11959], Fresh[11958], Fresh[11957], Fresh[11956], Fresh[11955], Fresh[11954], Fresh[11953], Fresh[11952], Fresh[11951], Fresh[11950], Fresh[11949], Fresh[11948], Fresh[11947], Fresh[11946], Fresh[11945], Fresh[11944], Fresh[11943], Fresh[11942], Fresh[11941], Fresh[11940], Fresh[11939], Fresh[11938], Fresh[11937], Fresh[11936], Fresh[11935], Fresh[11934], Fresh[11933], Fresh[11932], Fresh[11931], Fresh[11930], Fresh[11929], Fresh[11928], Fresh[11927], Fresh[11926], Fresh[11925], Fresh[11924], Fresh[11923], Fresh[11922], Fresh[11921], Fresh[11920], Fresh[11919], Fresh[11918], Fresh[11917], Fresh[11916], Fresh[11915], Fresh[11914], Fresh[11913], Fresh[11912], Fresh[11911], Fresh[11910], Fresh[11909], Fresh[11908], Fresh[11907], Fresh[11906], Fresh[11905], Fresh[11904], Fresh[11903], Fresh[11902], Fresh[11901], Fresh[11900], Fresh[11899], Fresh[11898], Fresh[11897], Fresh[11896], Fresh[11895], Fresh[11894], Fresh[11893], Fresh[11892], Fresh[11891], Fresh[11890], Fresh[11889], Fresh[11888], Fresh[11887], Fresh[11886], Fresh[11885], Fresh[11884], Fresh[11883], Fresh[11882], Fresh[11881], Fresh[11880], Fresh[11879], Fresh[11878], Fresh[11877], Fresh[11876], Fresh[11875], Fresh[11874], Fresh[11873], Fresh[11872], Fresh[11871], Fresh[11870], Fresh[11869], Fresh[11868], Fresh[11867], Fresh[11866], Fresh[11865], Fresh[11864], Fresh[11863], Fresh[11862], Fresh[11861], Fresh[11860], Fresh[11859], Fresh[11858], Fresh[11857], Fresh[11856], Fresh[11855], Fresh[11854], Fresh[11853], Fresh[11852], Fresh[11851], Fresh[11850], Fresh[11849], Fresh[11848], Fresh[11847], Fresh[11846], Fresh[11845], Fresh[11844], Fresh[11843], Fresh[11842], Fresh[11841], Fresh[11840], Fresh[11839], Fresh[11838], Fresh[11837], Fresh[11836], Fresh[11835], Fresh[11834], Fresh[11833], Fresh[11832], Fresh[11831], Fresh[11830], Fresh[11829], Fresh[11828], Fresh[11827], Fresh[11826], Fresh[11825], Fresh[11824], Fresh[11823], Fresh[11822], Fresh[11821], Fresh[11820], Fresh[11819], Fresh[11818], Fresh[11817], Fresh[11816], Fresh[11815], Fresh[11814], Fresh[11813], Fresh[11812], Fresh[11811], Fresh[11810], Fresh[11809], Fresh[11808], Fresh[11807], Fresh[11806], Fresh[11805], Fresh[11804], Fresh[11803], Fresh[11802], Fresh[11801], Fresh[11800], Fresh[11799], Fresh[11798], Fresh[11797], Fresh[11796], Fresh[11795], Fresh[11794], Fresh[11793], Fresh[11792], Fresh[11791], Fresh[11790], Fresh[11789], Fresh[11788], Fresh[11787], Fresh[11786], Fresh[11785], Fresh[11784], Fresh[11783], Fresh[11782], Fresh[11781], Fresh[11780], Fresh[11779], Fresh[11778], Fresh[11777], Fresh[11776], Fresh[11775], Fresh[11774], Fresh[11773], Fresh[11772], Fresh[11771], Fresh[11770], Fresh[11769], Fresh[11768], Fresh[11767], Fresh[11766], Fresh[11765], Fresh[11764], Fresh[11763], Fresh[11762], Fresh[11761], Fresh[11760], Fresh[11759], Fresh[11758], Fresh[11757], Fresh[11756], Fresh[11755], Fresh[11754], Fresh[11753], Fresh[11752], Fresh[11751], Fresh[11750], Fresh[11749], Fresh[11748], Fresh[11747], Fresh[11746], Fresh[11745], Fresh[11744], Fresh[11743], Fresh[11742], Fresh[11741], Fresh[11740], Fresh[11739], Fresh[11738], Fresh[11737], Fresh[11736], Fresh[11735], Fresh[11734], Fresh[11733], Fresh[11732], Fresh[11731], Fresh[11730], Fresh[11729], Fresh[11728], Fresh[11727], Fresh[11726], Fresh[11725], Fresh[11724], Fresh[11723], Fresh[11722], Fresh[11721], Fresh[11720], Fresh[11719], Fresh[11718], Fresh[11717], Fresh[11716], Fresh[11715], Fresh[11714], Fresh[11713], Fresh[11712], Fresh[11711], Fresh[11710], Fresh[11709], Fresh[11708], Fresh[11707], Fresh[11706], Fresh[11705], Fresh[11704], Fresh[11703], Fresh[11702], Fresh[11701], Fresh[11700], Fresh[11699], Fresh[11698], Fresh[11697], Fresh[11696], Fresh[11695], Fresh[11694], Fresh[11693], Fresh[11692], Fresh[11691], Fresh[11690], Fresh[11689], Fresh[11688], Fresh[11687], Fresh[11686], Fresh[11685], Fresh[11684], Fresh[11683], Fresh[11682], Fresh[11681], Fresh[11680], Fresh[11679], Fresh[11678], Fresh[11677], Fresh[11676], Fresh[11675], Fresh[11674], Fresh[11673], Fresh[11672], Fresh[11671], Fresh[11670], Fresh[11669], Fresh[11668], Fresh[11667], Fresh[11666], Fresh[11665], Fresh[11664], Fresh[11663], Fresh[11662], Fresh[11661], Fresh[11660], Fresh[11659], Fresh[11658], Fresh[11657], Fresh[11656], Fresh[11655], Fresh[11654], Fresh[11653], Fresh[11652], Fresh[11651], Fresh[11650], Fresh[11649], Fresh[11648], Fresh[11647], Fresh[11646], Fresh[11645], Fresh[11644], Fresh[11643], Fresh[11642], Fresh[11641], Fresh[11640], Fresh[11639], Fresh[11638], Fresh[11637], Fresh[11636], Fresh[11635], Fresh[11634], Fresh[11633], Fresh[11632], Fresh[11631], Fresh[11630], Fresh[11629], Fresh[11628], Fresh[11627], Fresh[11626], Fresh[11625], Fresh[11624], Fresh[11623], Fresh[11622], Fresh[11621], Fresh[11620], Fresh[11619], Fresh[11618], Fresh[11617], Fresh[11616], Fresh[11615], Fresh[11614], Fresh[11613], Fresh[11612], Fresh[11611], Fresh[11610], Fresh[11609], Fresh[11608], Fresh[11607], Fresh[11606], Fresh[11605], Fresh[11604], Fresh[11603], Fresh[11602], Fresh[11601], Fresh[11600], Fresh[11599], Fresh[11598], Fresh[11597], Fresh[11596], Fresh[11595], Fresh[11594], Fresh[11593], Fresh[11592], Fresh[11591], Fresh[11590], Fresh[11589], Fresh[11588], Fresh[11587], Fresh[11586], Fresh[11585], Fresh[11584], Fresh[11583], Fresh[11582], Fresh[11581], Fresh[11580], Fresh[11579], Fresh[11578], Fresh[11577], Fresh[11576], Fresh[11575], Fresh[11574], Fresh[11573], Fresh[11572], Fresh[11571], Fresh[11570], Fresh[11569], Fresh[11568], Fresh[11567], Fresh[11566], Fresh[11565], Fresh[11564], Fresh[11563], Fresh[11562], Fresh[11561], Fresh[11560], Fresh[11559], Fresh[11558], Fresh[11557], Fresh[11556], Fresh[11555], Fresh[11554], Fresh[11553], Fresh[11552], Fresh[11551], Fresh[11550], Fresh[11549], Fresh[11548], Fresh[11547], Fresh[11546], Fresh[11545], Fresh[11544], Fresh[11543], Fresh[11542], Fresh[11541], Fresh[11540], Fresh[11539], Fresh[11538], Fresh[11537], Fresh[11536], Fresh[11535], Fresh[11534], Fresh[11533], Fresh[11532], Fresh[11531], Fresh[11530], Fresh[11529], Fresh[11528], Fresh[11527], Fresh[11526], Fresh[11525], Fresh[11524], Fresh[11523], Fresh[11522], Fresh[11521], Fresh[11520], Fresh[11519], Fresh[11518], Fresh[11517], Fresh[11516], Fresh[11515], Fresh[11514], Fresh[11513], Fresh[11512], Fresh[11511], Fresh[11510], Fresh[11509], Fresh[11508], Fresh[11507], Fresh[11506], Fresh[11505], Fresh[11504], Fresh[11503], Fresh[11502], Fresh[11501], Fresh[11500], Fresh[11499], Fresh[11498], Fresh[11497], Fresh[11496], Fresh[11495], Fresh[11494], Fresh[11493], Fresh[11492], Fresh[11491], Fresh[11490], Fresh[11489], Fresh[11488], Fresh[11487], Fresh[11486], Fresh[11485], Fresh[11484], Fresh[11483], Fresh[11482], Fresh[11481], Fresh[11480], Fresh[11479], Fresh[11478], Fresh[11477], Fresh[11476], Fresh[11475], Fresh[11474], Fresh[11473], Fresh[11472], Fresh[11471], Fresh[11470], Fresh[11469], Fresh[11468], Fresh[11467], Fresh[11466], Fresh[11465], Fresh[11464], Fresh[11463], Fresh[11462], Fresh[11461], Fresh[11460], Fresh[11459], Fresh[11458], Fresh[11457], Fresh[11456], Fresh[11455], Fresh[11454], Fresh[11453], Fresh[11452], Fresh[11451], Fresh[11450], Fresh[11449], Fresh[11448], Fresh[11447], Fresh[11446], Fresh[11445], Fresh[11444], Fresh[11443], Fresh[11442], Fresh[11441], Fresh[11440], Fresh[11439], Fresh[11438], Fresh[11437], Fresh[11436], Fresh[11435], Fresh[11434], Fresh[11433], Fresh[11432], Fresh[11431], Fresh[11430], Fresh[11429], Fresh[11428], Fresh[11427], Fresh[11426], Fresh[11425], Fresh[11424], Fresh[11423], Fresh[11422], Fresh[11421], Fresh[11420], Fresh[11419], Fresh[11418], Fresh[11417], Fresh[11416], Fresh[11415], Fresh[11414], Fresh[11413], Fresh[11412], Fresh[11411], Fresh[11410], Fresh[11409], Fresh[11408], Fresh[11407], Fresh[11406], Fresh[11405], Fresh[11404], Fresh[11403], Fresh[11402], Fresh[11401], Fresh[11400], Fresh[11399], Fresh[11398], Fresh[11397], Fresh[11396], Fresh[11395], Fresh[11394], Fresh[11393], Fresh[11392], Fresh[11391], Fresh[11390], Fresh[11389], Fresh[11388], Fresh[11387], Fresh[11386], Fresh[11385], Fresh[11384], Fresh[11383], Fresh[11382], Fresh[11381], Fresh[11380], Fresh[11379], Fresh[11378], Fresh[11377], Fresh[11376], Fresh[11375], Fresh[11374], Fresh[11373], Fresh[11372], Fresh[11371], Fresh[11370], Fresh[11369], Fresh[11368], Fresh[11367], Fresh[11366], Fresh[11365], Fresh[11364], Fresh[11363], Fresh[11362], Fresh[11361], Fresh[11360], Fresh[11359], Fresh[11358], Fresh[11357], Fresh[11356], Fresh[11355], Fresh[11354], Fresh[11353], Fresh[11352], Fresh[11351], Fresh[11350], Fresh[11349], Fresh[11348], Fresh[11347], Fresh[11346], Fresh[11345], Fresh[11344], Fresh[11343], Fresh[11342], Fresh[11341], Fresh[11340], Fresh[11339], Fresh[11338], Fresh[11337], Fresh[11336], Fresh[11335], Fresh[11334], Fresh[11333], Fresh[11332], Fresh[11331], Fresh[11330], Fresh[11329], Fresh[11328], Fresh[11327], Fresh[11326], Fresh[11325], Fresh[11324], Fresh[11323], Fresh[11322], Fresh[11321], Fresh[11320], Fresh[11319], Fresh[11318], Fresh[11317], Fresh[11316], Fresh[11315], Fresh[11314], Fresh[11313], Fresh[11312], Fresh[11311], Fresh[11310], Fresh[11309], Fresh[11308], Fresh[11307], Fresh[11306], Fresh[11305], Fresh[11304], Fresh[11303], Fresh[11302], Fresh[11301], Fresh[11300], Fresh[11299], Fresh[11298], Fresh[11297], Fresh[11296], Fresh[11295], Fresh[11294], Fresh[11293], Fresh[11292], Fresh[11291], Fresh[11290], Fresh[11289], Fresh[11288], Fresh[11287], Fresh[11286], Fresh[11285], Fresh[11284], Fresh[11283], Fresh[11282], Fresh[11281], Fresh[11280], Fresh[11279], Fresh[11278], Fresh[11277], Fresh[11276], Fresh[11275], Fresh[11274], Fresh[11273], Fresh[11272], Fresh[11271], Fresh[11270], Fresh[11269], Fresh[11268], Fresh[11267], Fresh[11266], Fresh[11265], Fresh[11264], Fresh[11263], Fresh[11262], Fresh[11261], Fresh[11260], Fresh[11259], Fresh[11258], Fresh[11257], Fresh[11256], Fresh[11255], Fresh[11254], Fresh[11253], Fresh[11252], Fresh[11251], Fresh[11250], Fresh[11249], Fresh[11248], Fresh[11247], Fresh[11246], Fresh[11245], Fresh[11244], Fresh[11243], Fresh[11242], Fresh[11241], Fresh[11240], Fresh[11239], Fresh[11238], Fresh[11237], Fresh[11236], Fresh[11235], Fresh[11234], Fresh[11233], Fresh[11232], Fresh[11231], Fresh[11230], Fresh[11229], Fresh[11228], Fresh[11227], Fresh[11226], Fresh[11225], Fresh[11224], Fresh[11223], Fresh[11222], Fresh[11221], Fresh[11220], Fresh[11219], Fresh[11218], Fresh[11217], Fresh[11216], Fresh[11215], Fresh[11214], Fresh[11213], Fresh[11212], Fresh[11211], Fresh[11210], Fresh[11209], Fresh[11208], Fresh[11207], Fresh[11206], Fresh[11205], Fresh[11204], Fresh[11203], Fresh[11202], Fresh[11201], Fresh[11200], Fresh[11199], Fresh[11198], Fresh[11197], Fresh[11196], Fresh[11195], Fresh[11194], Fresh[11193], Fresh[11192], Fresh[11191], Fresh[11190], Fresh[11189], Fresh[11188], Fresh[11187], Fresh[11186], Fresh[11185], Fresh[11184], Fresh[11183], Fresh[11182], Fresh[11181], Fresh[11180], Fresh[11179], Fresh[11178], Fresh[11177], Fresh[11176], Fresh[11175], Fresh[11174], Fresh[11173], Fresh[11172], Fresh[11171], Fresh[11170], Fresh[11169], Fresh[11168], Fresh[11167], Fresh[11166], Fresh[11165], Fresh[11164], Fresh[11163], Fresh[11162], Fresh[11161], Fresh[11160], Fresh[11159], Fresh[11158], Fresh[11157], Fresh[11156], Fresh[11155], Fresh[11154], Fresh[11153], Fresh[11152], Fresh[11151], Fresh[11150], Fresh[11149], Fresh[11148], Fresh[11147], Fresh[11146], Fresh[11145], Fresh[11144], Fresh[11143], Fresh[11142], Fresh[11141], Fresh[11140], Fresh[11139], Fresh[11138], Fresh[11137], Fresh[11136], Fresh[11135], Fresh[11134], Fresh[11133], Fresh[11132], Fresh[11131], Fresh[11130], Fresh[11129], Fresh[11128], Fresh[11127], Fresh[11126], Fresh[11125], Fresh[11124], Fresh[11123], Fresh[11122], Fresh[11121], Fresh[11120], Fresh[11119], Fresh[11118], Fresh[11117], Fresh[11116], Fresh[11115], Fresh[11114], Fresh[11113], Fresh[11112], Fresh[11111], Fresh[11110], Fresh[11109], Fresh[11108], Fresh[11107], Fresh[11106], Fresh[11105], Fresh[11104], Fresh[11103], Fresh[11102], Fresh[11101], Fresh[11100], Fresh[11099], Fresh[11098], Fresh[11097], Fresh[11096], Fresh[11095], Fresh[11094], Fresh[11093], Fresh[11092], Fresh[11091], Fresh[11090], Fresh[11089], Fresh[11088], Fresh[11087], Fresh[11086], Fresh[11085], Fresh[11084], Fresh[11083], Fresh[11082], Fresh[11081], Fresh[11080], Fresh[11079], Fresh[11078], Fresh[11077], Fresh[11076], Fresh[11075], Fresh[11074], Fresh[11073], Fresh[11072], Fresh[11071], Fresh[11070], Fresh[11069], Fresh[11068], Fresh[11067], Fresh[11066], Fresh[11065], Fresh[11064], Fresh[11063], Fresh[11062], Fresh[11061], Fresh[11060], Fresh[11059], Fresh[11058], Fresh[11057], Fresh[11056], Fresh[11055], Fresh[11054], Fresh[11053], Fresh[11052], Fresh[11051], Fresh[11050], Fresh[11049], Fresh[11048], Fresh[11047], Fresh[11046], Fresh[11045], Fresh[11044], Fresh[11043], Fresh[11042], Fresh[11041], Fresh[11040], Fresh[11039], Fresh[11038], Fresh[11037], Fresh[11036], Fresh[11035], Fresh[11034], Fresh[11033], Fresh[11032], Fresh[11031], Fresh[11030], Fresh[11029], Fresh[11028], Fresh[11027], Fresh[11026], Fresh[11025], Fresh[11024], Fresh[11023], Fresh[11022], Fresh[11021], Fresh[11020], Fresh[11019], Fresh[11018], Fresh[11017], Fresh[11016], Fresh[11015], Fresh[11014], Fresh[11013], Fresh[11012], Fresh[11011], Fresh[11010], Fresh[11009], Fresh[11008], Fresh[11007], Fresh[11006], Fresh[11005], Fresh[11004], Fresh[11003], Fresh[11002], Fresh[11001], Fresh[11000], Fresh[10999], Fresh[10998], Fresh[10997], Fresh[10996], Fresh[10995], Fresh[10994], Fresh[10993], Fresh[10992], Fresh[10991], Fresh[10990], Fresh[10989], Fresh[10988], Fresh[10987], Fresh[10986], Fresh[10985], Fresh[10984], Fresh[10983], Fresh[10982], Fresh[10981], Fresh[10980], Fresh[10979], Fresh[10978], Fresh[10977], Fresh[10976], Fresh[10975], Fresh[10974], Fresh[10973], Fresh[10972], Fresh[10971], Fresh[10970], Fresh[10969], Fresh[10968], Fresh[10967], Fresh[10966], Fresh[10965], Fresh[10964], Fresh[10963], Fresh[10962], Fresh[10961], Fresh[10960], Fresh[10959], Fresh[10958], Fresh[10957], Fresh[10956], Fresh[10955], Fresh[10954], Fresh[10953], Fresh[10952], Fresh[10951], Fresh[10950], Fresh[10949], Fresh[10948], Fresh[10947], Fresh[10946], Fresh[10945], Fresh[10944], Fresh[10943], Fresh[10942], Fresh[10941], Fresh[10940], Fresh[10939], Fresh[10938], Fresh[10937], Fresh[10936], Fresh[10935], Fresh[10934], Fresh[10933], Fresh[10932], Fresh[10931], Fresh[10930], Fresh[10929], Fresh[10928], Fresh[10927], Fresh[10926], Fresh[10925], Fresh[10924], Fresh[10923], Fresh[10922], Fresh[10921], Fresh[10920], Fresh[10919], Fresh[10918], Fresh[10917], Fresh[10916], Fresh[10915], Fresh[10914], Fresh[10913], Fresh[10912], Fresh[10911], Fresh[10910], Fresh[10909], Fresh[10908], Fresh[10907], Fresh[10906], Fresh[10905], Fresh[10904], Fresh[10903], Fresh[10902], Fresh[10901], Fresh[10900], Fresh[10899], Fresh[10898], Fresh[10897], Fresh[10896], Fresh[10895], Fresh[10894], Fresh[10893], Fresh[10892], Fresh[10891], Fresh[10890], Fresh[10889], Fresh[10888], Fresh[10887], Fresh[10886], Fresh[10885], Fresh[10884], Fresh[10883], Fresh[10882], Fresh[10881], Fresh[10880], Fresh[10879], Fresh[10878], Fresh[10877], Fresh[10876], Fresh[10875], Fresh[10874], Fresh[10873], Fresh[10872], Fresh[10871], Fresh[10870], Fresh[10869], Fresh[10868], Fresh[10867], Fresh[10866], Fresh[10865], Fresh[10864], Fresh[10863], Fresh[10862], Fresh[10861], Fresh[10860], Fresh[10859], Fresh[10858], Fresh[10857], Fresh[10856], Fresh[10855], Fresh[10854], Fresh[10853], Fresh[10852], Fresh[10851], Fresh[10850], Fresh[10849], Fresh[10848], Fresh[10847], Fresh[10846], Fresh[10845], Fresh[10844], Fresh[10843], Fresh[10842], Fresh[10841], Fresh[10840], Fresh[10839], Fresh[10838], Fresh[10837], Fresh[10836], Fresh[10835], Fresh[10834], Fresh[10833], Fresh[10832], Fresh[10831], Fresh[10830], Fresh[10829], Fresh[10828], Fresh[10827], Fresh[10826], Fresh[10825], Fresh[10824], Fresh[10823], Fresh[10822], Fresh[10821], Fresh[10820], Fresh[10819], Fresh[10818], Fresh[10817], Fresh[10816], Fresh[10815], Fresh[10814], Fresh[10813], Fresh[10812], Fresh[10811], Fresh[10810], Fresh[10809], Fresh[10808], Fresh[10807], Fresh[10806], Fresh[10805], Fresh[10804], Fresh[10803], Fresh[10802], Fresh[10801], Fresh[10800], Fresh[10799], Fresh[10798], Fresh[10797], Fresh[10796], Fresh[10795], Fresh[10794], Fresh[10793], Fresh[10792], Fresh[10791], Fresh[10790], Fresh[10789], Fresh[10788], Fresh[10787], Fresh[10786], Fresh[10785], Fresh[10784], Fresh[10783], Fresh[10782], Fresh[10781], Fresh[10780], Fresh[10779], Fresh[10778], Fresh[10777], Fresh[10776], Fresh[10775], Fresh[10774], Fresh[10773], Fresh[10772], Fresh[10771], Fresh[10770], Fresh[10769], Fresh[10768], Fresh[10767], Fresh[10766], Fresh[10765], Fresh[10764], Fresh[10763], Fresh[10762], Fresh[10761], Fresh[10760], Fresh[10759], Fresh[10758], Fresh[10757], Fresh[10756], Fresh[10755], Fresh[10754], Fresh[10753], Fresh[10752], Fresh[10751], Fresh[10750], Fresh[10749], Fresh[10748], Fresh[10747], Fresh[10746], Fresh[10745], Fresh[10744], Fresh[10743], Fresh[10742], Fresh[10741], Fresh[10740], Fresh[10739], Fresh[10738], Fresh[10737], Fresh[10736], Fresh[10735], Fresh[10734], Fresh[10733], Fresh[10732], Fresh[10731], Fresh[10730], Fresh[10729], Fresh[10728], Fresh[10727], Fresh[10726], Fresh[10725], Fresh[10724], Fresh[10723], Fresh[10722], Fresh[10721], Fresh[10720], Fresh[10719], Fresh[10718], Fresh[10717], Fresh[10716], Fresh[10715], Fresh[10714], Fresh[10713], Fresh[10712], Fresh[10711], Fresh[10710], Fresh[10709], Fresh[10708], Fresh[10707], Fresh[10706], Fresh[10705], Fresh[10704], Fresh[10703], Fresh[10702], Fresh[10701], Fresh[10700], Fresh[10699], Fresh[10698], Fresh[10697], Fresh[10696], Fresh[10695], Fresh[10694], Fresh[10693], Fresh[10692], Fresh[10691], Fresh[10690], Fresh[10689], Fresh[10688], Fresh[10687], Fresh[10686], Fresh[10685], Fresh[10684], Fresh[10683], Fresh[10682], Fresh[10681], Fresh[10680], Fresh[10679], Fresh[10678], Fresh[10677], Fresh[10676], Fresh[10675], Fresh[10674], Fresh[10673], Fresh[10672], Fresh[10671], Fresh[10670], Fresh[10669], Fresh[10668], Fresh[10667], Fresh[10666], Fresh[10665], Fresh[10664], Fresh[10663], Fresh[10662], Fresh[10661], Fresh[10660], Fresh[10659], Fresh[10658], Fresh[10657], Fresh[10656], Fresh[10655], Fresh[10654], Fresh[10653], Fresh[10652], Fresh[10651], Fresh[10650], Fresh[10649], Fresh[10648], Fresh[10647], Fresh[10646], Fresh[10645], Fresh[10644], Fresh[10643], Fresh[10642], Fresh[10641], Fresh[10640], Fresh[10639], Fresh[10638], Fresh[10637], Fresh[10636], Fresh[10635], Fresh[10634], Fresh[10633], Fresh[10632], Fresh[10631], Fresh[10630], Fresh[10629], Fresh[10628], Fresh[10627], Fresh[10626], Fresh[10625], Fresh[10624], Fresh[10623], Fresh[10622], Fresh[10621], Fresh[10620], Fresh[10619], Fresh[10618], Fresh[10617], Fresh[10616], Fresh[10615], Fresh[10614], Fresh[10613], Fresh[10612], Fresh[10611], Fresh[10610], Fresh[10609], Fresh[10608], Fresh[10607], Fresh[10606], Fresh[10605], Fresh[10604], Fresh[10603], Fresh[10602], Fresh[10601], Fresh[10600], Fresh[10599], Fresh[10598], Fresh[10597], Fresh[10596], Fresh[10595], Fresh[10594], Fresh[10593], Fresh[10592], Fresh[10591], Fresh[10590], Fresh[10589], Fresh[10588], Fresh[10587], Fresh[10586], Fresh[10585], Fresh[10584], Fresh[10583], Fresh[10582], Fresh[10581], Fresh[10580], Fresh[10579], Fresh[10578], Fresh[10577], Fresh[10576], Fresh[10575], Fresh[10574], Fresh[10573], Fresh[10572], Fresh[10571], Fresh[10570], Fresh[10569], Fresh[10568], Fresh[10567], Fresh[10566], Fresh[10565], Fresh[10564], Fresh[10563], Fresh[10562], Fresh[10561], Fresh[10560], Fresh[10559], Fresh[10558], Fresh[10557], Fresh[10556], Fresh[10555], Fresh[10554], Fresh[10553], Fresh[10552], Fresh[10551], Fresh[10550], Fresh[10549], Fresh[10548], Fresh[10547], Fresh[10546], Fresh[10545], Fresh[10544], Fresh[10543], Fresh[10542], Fresh[10541], Fresh[10540], Fresh[10539], Fresh[10538], Fresh[10537], Fresh[10536], Fresh[10535], Fresh[10534], Fresh[10533], Fresh[10532], Fresh[10531], Fresh[10530], Fresh[10529], Fresh[10528], Fresh[10527], Fresh[10526], Fresh[10525], Fresh[10524], Fresh[10523], Fresh[10522], Fresh[10521], Fresh[10520], Fresh[10519], Fresh[10518], Fresh[10517], Fresh[10516], Fresh[10515], Fresh[10514], Fresh[10513], Fresh[10512], Fresh[10511], Fresh[10510], Fresh[10509], Fresh[10508], Fresh[10507], Fresh[10506], Fresh[10505], Fresh[10504], Fresh[10503], Fresh[10502], Fresh[10501], Fresh[10500], Fresh[10499], Fresh[10498], Fresh[10497], Fresh[10496], Fresh[10495], Fresh[10494], Fresh[10493], Fresh[10492], Fresh[10491], Fresh[10490], Fresh[10489], Fresh[10488], Fresh[10487], Fresh[10486], Fresh[10485], Fresh[10484], Fresh[10483], Fresh[10482], Fresh[10481], Fresh[10480], Fresh[10479], Fresh[10478], Fresh[10477], Fresh[10476], Fresh[10475], Fresh[10474], Fresh[10473], Fresh[10472], Fresh[10471], Fresh[10470], Fresh[10469], Fresh[10468], Fresh[10467], Fresh[10466], Fresh[10465], Fresh[10464], Fresh[10463], Fresh[10462], Fresh[10461], Fresh[10460], Fresh[10459], Fresh[10458], Fresh[10457], Fresh[10456], Fresh[10455], Fresh[10454], Fresh[10453], Fresh[10452], Fresh[10451], Fresh[10450], Fresh[10449], Fresh[10448], Fresh[10447], Fresh[10446], Fresh[10445], Fresh[10444], Fresh[10443], Fresh[10442], Fresh[10441], Fresh[10440], Fresh[10439], Fresh[10438], Fresh[10437], Fresh[10436], Fresh[10435], Fresh[10434], Fresh[10433], Fresh[10432], Fresh[10431], Fresh[10430], Fresh[10429], Fresh[10428], Fresh[10427], Fresh[10426], Fresh[10425], Fresh[10424], Fresh[10423], Fresh[10422], Fresh[10421], Fresh[10420], Fresh[10419], Fresh[10418], Fresh[10417], Fresh[10416], Fresh[10415], Fresh[10414], Fresh[10413], Fresh[10412], Fresh[10411], Fresh[10410], Fresh[10409], Fresh[10408], Fresh[10407], Fresh[10406], Fresh[10405], Fresh[10404], Fresh[10403], Fresh[10402], Fresh[10401], Fresh[10400], Fresh[10399], Fresh[10398], Fresh[10397], Fresh[10396], Fresh[10395], Fresh[10394], Fresh[10393], Fresh[10392], Fresh[10391], Fresh[10390], Fresh[10389], Fresh[10388], Fresh[10387], Fresh[10386], Fresh[10385], Fresh[10384], Fresh[10383], Fresh[10382], Fresh[10381], Fresh[10380], Fresh[10379], Fresh[10378], Fresh[10377], Fresh[10376], Fresh[10375], Fresh[10374], Fresh[10373], Fresh[10372], Fresh[10371], Fresh[10370], Fresh[10369], Fresh[10368], Fresh[10367], Fresh[10366], Fresh[10365], Fresh[10364], Fresh[10363], Fresh[10362], Fresh[10361], Fresh[10360], Fresh[10359], Fresh[10358], Fresh[10357], Fresh[10356], Fresh[10355], Fresh[10354], Fresh[10353], Fresh[10352], Fresh[10351], Fresh[10350], Fresh[10349], Fresh[10348], Fresh[10347], Fresh[10346], Fresh[10345], Fresh[10344], Fresh[10343], Fresh[10342], Fresh[10341], Fresh[10340], Fresh[10339], Fresh[10338], Fresh[10337], Fresh[10336], Fresh[10335], Fresh[10334], Fresh[10333], Fresh[10332], Fresh[10331], Fresh[10330], Fresh[10329], Fresh[10328], Fresh[10327], Fresh[10326], Fresh[10325], Fresh[10324], Fresh[10323], Fresh[10322], Fresh[10321], Fresh[10320], Fresh[10319], Fresh[10318], Fresh[10317], Fresh[10316], Fresh[10315], Fresh[10314], Fresh[10313], Fresh[10312], Fresh[10311], Fresh[10310], Fresh[10309], Fresh[10308], Fresh[10307], Fresh[10306], Fresh[10305], Fresh[10304], Fresh[10303], Fresh[10302], Fresh[10301], Fresh[10300], Fresh[10299], Fresh[10298], Fresh[10297], Fresh[10296], Fresh[10295], Fresh[10294], Fresh[10293], Fresh[10292], Fresh[10291], Fresh[10290], Fresh[10289], Fresh[10288], Fresh[10287], Fresh[10286], Fresh[10285], Fresh[10284], Fresh[10283], Fresh[10282], Fresh[10281], Fresh[10280], Fresh[10279], Fresh[10278], Fresh[10277], Fresh[10276], Fresh[10275], Fresh[10274], Fresh[10273], Fresh[10272], Fresh[10271], Fresh[10270], Fresh[10269], Fresh[10268], Fresh[10267], Fresh[10266], Fresh[10265], Fresh[10264], Fresh[10263], Fresh[10262], Fresh[10261], Fresh[10260], Fresh[10259], Fresh[10258], Fresh[10257], Fresh[10256], Fresh[10255], Fresh[10254], Fresh[10253], Fresh[10252], Fresh[10251], Fresh[10250], Fresh[10249], Fresh[10248], Fresh[10247], Fresh[10246], Fresh[10245], Fresh[10244], Fresh[10243], Fresh[10242], Fresh[10241], Fresh[10240], Fresh[10239], Fresh[10238], Fresh[10237], Fresh[10236], Fresh[10235], Fresh[10234], Fresh[10233], Fresh[10232], Fresh[10231], Fresh[10230], Fresh[10229], Fresh[10228], Fresh[10227], Fresh[10226], Fresh[10225], Fresh[10224], Fresh[10223], Fresh[10222], Fresh[10221], Fresh[10220], Fresh[10219], Fresh[10218], Fresh[10217], Fresh[10216], Fresh[10215], Fresh[10214], Fresh[10213], Fresh[10212], Fresh[10211], Fresh[10210], Fresh[10209], Fresh[10208], Fresh[10207], Fresh[10206], Fresh[10205], Fresh[10204], Fresh[10203], Fresh[10202], Fresh[10201], Fresh[10200], Fresh[10199], Fresh[10198], Fresh[10197], Fresh[10196], Fresh[10195], Fresh[10194], Fresh[10193], Fresh[10192], Fresh[10191], Fresh[10190], Fresh[10189], Fresh[10188], Fresh[10187], Fresh[10186], Fresh[10185], Fresh[10184], Fresh[10183], Fresh[10182], Fresh[10181], Fresh[10180], Fresh[10179], Fresh[10178], Fresh[10177], Fresh[10176], Fresh[10175], Fresh[10174], Fresh[10173], Fresh[10172], Fresh[10171], Fresh[10170], Fresh[10169], Fresh[10168], Fresh[10167], Fresh[10166], Fresh[10165], Fresh[10164], Fresh[10163], Fresh[10162], Fresh[10161], Fresh[10160], Fresh[10159], Fresh[10158], Fresh[10157], Fresh[10156], Fresh[10155], Fresh[10154], Fresh[10153], Fresh[10152], Fresh[10151], Fresh[10150], Fresh[10149], Fresh[10148], Fresh[10147], Fresh[10146], Fresh[10145], Fresh[10144], Fresh[10143], Fresh[10142], Fresh[10141], Fresh[10140], Fresh[10139], Fresh[10138], Fresh[10137], Fresh[10136], Fresh[10135], Fresh[10134], Fresh[10133], Fresh[10132], Fresh[10131], Fresh[10130], Fresh[10129], Fresh[10128], Fresh[10127], Fresh[10126], Fresh[10125], Fresh[10124], Fresh[10123], Fresh[10122], Fresh[10121], Fresh[10120], Fresh[10119], Fresh[10118], Fresh[10117], Fresh[10116], Fresh[10115], Fresh[10114], Fresh[10113], Fresh[10112], Fresh[10111], Fresh[10110], Fresh[10109], Fresh[10108], Fresh[10107], Fresh[10106], Fresh[10105], Fresh[10104], Fresh[10103], Fresh[10102], Fresh[10101], Fresh[10100], Fresh[10099], Fresh[10098], Fresh[10097], Fresh[10096], Fresh[10095], Fresh[10094], Fresh[10093], Fresh[10092], Fresh[10091], Fresh[10090], Fresh[10089], Fresh[10088], Fresh[10087], Fresh[10086], Fresh[10085], Fresh[10084], Fresh[10083], Fresh[10082], Fresh[10081], Fresh[10080], Fresh[10079], Fresh[10078], Fresh[10077], Fresh[10076], Fresh[10075], Fresh[10074], Fresh[10073], Fresh[10072], Fresh[10071], Fresh[10070], Fresh[10069], Fresh[10068], Fresh[10067], Fresh[10066], Fresh[10065], Fresh[10064], Fresh[10063], Fresh[10062], Fresh[10061], Fresh[10060], Fresh[10059], Fresh[10058], Fresh[10057], Fresh[10056], Fresh[10055], Fresh[10054], Fresh[10053], Fresh[10052], Fresh[10051], Fresh[10050], Fresh[10049], Fresh[10048], Fresh[10047], Fresh[10046], Fresh[10045], Fresh[10044], Fresh[10043], Fresh[10042], Fresh[10041], Fresh[10040], Fresh[10039], Fresh[10038], Fresh[10037], Fresh[10036], Fresh[10035], Fresh[10034], Fresh[10033], Fresh[10032], Fresh[10031], Fresh[10030], Fresh[10029], Fresh[10028], Fresh[10027], Fresh[10026], Fresh[10025], Fresh[10024], Fresh[10023], Fresh[10022], Fresh[10021], Fresh[10020], Fresh[10019], Fresh[10018], Fresh[10017], Fresh[10016], Fresh[10015], Fresh[10014], Fresh[10013], Fresh[10012], Fresh[10011], Fresh[10010], Fresh[10009], Fresh[10008], Fresh[10007], Fresh[10006], Fresh[10005], Fresh[10004], Fresh[10003], Fresh[10002], Fresh[10001], Fresh[10000], Fresh[9999], Fresh[9998], Fresh[9997], Fresh[9996], Fresh[9995], Fresh[9994], Fresh[9993], Fresh[9992], Fresh[9991], Fresh[9990], Fresh[9989], Fresh[9988], Fresh[9987], Fresh[9986], Fresh[9985], Fresh[9984], Fresh[9983], Fresh[9982], Fresh[9981], Fresh[9980], Fresh[9979], Fresh[9978], Fresh[9977], Fresh[9976], Fresh[9975], Fresh[9974], Fresh[9973], Fresh[9972], Fresh[9971], Fresh[9970], Fresh[9969], Fresh[9968], Fresh[9967], Fresh[9966], Fresh[9965], Fresh[9964], Fresh[9963], Fresh[9962], Fresh[9961], Fresh[9960], Fresh[9959], Fresh[9958], Fresh[9957], Fresh[9956], Fresh[9955], Fresh[9954], Fresh[9953], Fresh[9952], Fresh[9951], Fresh[9950], Fresh[9949], Fresh[9948], Fresh[9947], Fresh[9946], Fresh[9945], Fresh[9944], Fresh[9943], Fresh[9942], Fresh[9941], Fresh[9940], Fresh[9939], Fresh[9938], Fresh[9937], Fresh[9936], Fresh[9935], Fresh[9934], Fresh[9933], Fresh[9932], Fresh[9931], Fresh[9930], Fresh[9929], Fresh[9928], Fresh[9927], Fresh[9926], Fresh[9925], Fresh[9924], Fresh[9923], Fresh[9922], Fresh[9921], Fresh[9920], Fresh[9919], Fresh[9918], Fresh[9917], Fresh[9916], Fresh[9915], Fresh[9914], Fresh[9913], Fresh[9912], Fresh[9911], Fresh[9910], Fresh[9909], Fresh[9908], Fresh[9907], Fresh[9906], Fresh[9905], Fresh[9904], Fresh[9903], Fresh[9902], Fresh[9901], Fresh[9900], Fresh[9899], Fresh[9898], Fresh[9897], Fresh[9896], Fresh[9895], Fresh[9894], Fresh[9893], Fresh[9892], Fresh[9891], Fresh[9890], Fresh[9889], Fresh[9888], Fresh[9887], Fresh[9886], Fresh[9885], Fresh[9884], Fresh[9883], Fresh[9882], Fresh[9881], Fresh[9880], Fresh[9879], Fresh[9878], Fresh[9877], Fresh[9876], Fresh[9875], Fresh[9874], Fresh[9873], Fresh[9872], Fresh[9871], Fresh[9870], Fresh[9869], Fresh[9868], Fresh[9867], Fresh[9866], Fresh[9865], Fresh[9864], Fresh[9863], Fresh[9862], Fresh[9861], Fresh[9860], Fresh[9859], Fresh[9858], Fresh[9857], Fresh[9856], Fresh[9855], Fresh[9854], Fresh[9853], Fresh[9852], Fresh[9851], Fresh[9850], Fresh[9849], Fresh[9848], Fresh[9847], Fresh[9846], Fresh[9845], Fresh[9844], Fresh[9843], Fresh[9842], Fresh[9841], Fresh[9840], Fresh[9839], Fresh[9838], Fresh[9837], Fresh[9836], Fresh[9835], Fresh[9834], Fresh[9833], Fresh[9832], Fresh[9831], Fresh[9830], Fresh[9829], Fresh[9828], Fresh[9827], Fresh[9826], Fresh[9825], Fresh[9824], Fresh[9823], Fresh[9822], Fresh[9821], Fresh[9820], Fresh[9819], Fresh[9818], Fresh[9817], Fresh[9816], Fresh[9815], Fresh[9814], Fresh[9813], Fresh[9812], Fresh[9811], Fresh[9810], Fresh[9809], Fresh[9808], Fresh[9807], Fresh[9806], Fresh[9805], Fresh[9804], Fresh[9803], Fresh[9802], Fresh[9801], Fresh[9800], Fresh[9799], Fresh[9798], Fresh[9797], Fresh[9796], Fresh[9795], Fresh[9794], Fresh[9793], Fresh[9792], Fresh[9791], Fresh[9790], Fresh[9789], Fresh[9788], Fresh[9787], Fresh[9786], Fresh[9785], Fresh[9784], Fresh[9783], Fresh[9782], Fresh[9781], Fresh[9780], Fresh[9779], Fresh[9778], Fresh[9777], Fresh[9776], Fresh[9775], Fresh[9774], Fresh[9773], Fresh[9772], Fresh[9771], Fresh[9770], Fresh[9769], Fresh[9768], Fresh[9767], Fresh[9766], Fresh[9765], Fresh[9764], Fresh[9763], Fresh[9762], Fresh[9761], Fresh[9760], Fresh[9759], Fresh[9758], Fresh[9757], Fresh[9756], Fresh[9755], Fresh[9754], Fresh[9753], Fresh[9752], Fresh[9751], Fresh[9750], Fresh[9749], Fresh[9748], Fresh[9747], Fresh[9746], Fresh[9745], Fresh[9744], Fresh[9743], Fresh[9742], Fresh[9741], Fresh[9740], Fresh[9739], Fresh[9738], Fresh[9737], Fresh[9736], Fresh[9735], Fresh[9734], Fresh[9733], Fresh[9732], Fresh[9731], Fresh[9730], Fresh[9729], Fresh[9728], Fresh[9727], Fresh[9726], Fresh[9725], Fresh[9724], Fresh[9723], Fresh[9722], Fresh[9721], Fresh[9720], Fresh[9719], Fresh[9718], Fresh[9717], Fresh[9716], Fresh[9715], Fresh[9714], Fresh[9713], Fresh[9712], Fresh[9711], Fresh[9710], Fresh[9709], Fresh[9708], Fresh[9707], Fresh[9706], Fresh[9705], Fresh[9704], Fresh[9703], Fresh[9702], Fresh[9701], Fresh[9700], Fresh[9699], Fresh[9698], Fresh[9697], Fresh[9696], Fresh[9695], Fresh[9694], Fresh[9693], Fresh[9692], Fresh[9691], Fresh[9690], Fresh[9689], Fresh[9688], Fresh[9687], Fresh[9686], Fresh[9685], Fresh[9684], Fresh[9683], Fresh[9682], Fresh[9681], Fresh[9680], Fresh[9679], Fresh[9678], Fresh[9677], Fresh[9676], Fresh[9675], Fresh[9674], Fresh[9673], Fresh[9672], Fresh[9671], Fresh[9670], Fresh[9669], Fresh[9668], Fresh[9667], Fresh[9666], Fresh[9665], Fresh[9664], Fresh[9663], Fresh[9662], Fresh[9661], Fresh[9660], Fresh[9659], Fresh[9658], Fresh[9657], Fresh[9656], Fresh[9655], Fresh[9654], Fresh[9653], Fresh[9652], Fresh[9651], Fresh[9650], Fresh[9649], Fresh[9648], Fresh[9647], Fresh[9646], Fresh[9645], Fresh[9644], Fresh[9643], Fresh[9642], Fresh[9641], Fresh[9640], Fresh[9639], Fresh[9638], Fresh[9637], Fresh[9636], Fresh[9635], Fresh[9634], Fresh[9633], Fresh[9632], Fresh[9631], Fresh[9630], Fresh[9629], Fresh[9628], Fresh[9627], Fresh[9626], Fresh[9625], Fresh[9624], Fresh[9623], Fresh[9622], Fresh[9621], Fresh[9620], Fresh[9619], Fresh[9618], Fresh[9617], Fresh[9616], Fresh[9615], Fresh[9614], Fresh[9613], Fresh[9612], Fresh[9611], Fresh[9610], Fresh[9609], Fresh[9608], Fresh[9607], Fresh[9606], Fresh[9605], Fresh[9604], Fresh[9603], Fresh[9602], Fresh[9601], Fresh[9600], Fresh[9599], Fresh[9598], Fresh[9597], Fresh[9596], Fresh[9595], Fresh[9594], Fresh[9593], Fresh[9592], Fresh[9591], Fresh[9590], Fresh[9589], Fresh[9588], Fresh[9587], Fresh[9586], Fresh[9585], Fresh[9584], Fresh[9583], Fresh[9582], Fresh[9581], Fresh[9580], Fresh[9579], Fresh[9578], Fresh[9577], Fresh[9576], Fresh[9575], Fresh[9574], Fresh[9573], Fresh[9572], Fresh[9571], Fresh[9570], Fresh[9569], Fresh[9568], Fresh[9567], Fresh[9566], Fresh[9565], Fresh[9564], Fresh[9563], Fresh[9562], Fresh[9561], Fresh[9560], Fresh[9559], Fresh[9558], Fresh[9557], Fresh[9556], Fresh[9555], Fresh[9554], Fresh[9553], Fresh[9552], Fresh[9551], Fresh[9550], Fresh[9549], Fresh[9548], Fresh[9547], Fresh[9546], Fresh[9545], Fresh[9544], Fresh[9543], Fresh[9542], Fresh[9541], Fresh[9540], Fresh[9539], Fresh[9538], Fresh[9537], Fresh[9536], Fresh[9535], Fresh[9534], Fresh[9533], Fresh[9532], Fresh[9531], Fresh[9530], Fresh[9529], Fresh[9528], Fresh[9527], Fresh[9526], Fresh[9525], Fresh[9524], Fresh[9523], Fresh[9522], Fresh[9521], Fresh[9520], Fresh[9519], Fresh[9518], Fresh[9517], Fresh[9516], Fresh[9515], Fresh[9514], Fresh[9513], Fresh[9512], Fresh[9511], Fresh[9510], Fresh[9509], Fresh[9508], Fresh[9507], Fresh[9506], Fresh[9505], Fresh[9504], Fresh[9503], Fresh[9502], Fresh[9501], Fresh[9500], Fresh[9499], Fresh[9498], Fresh[9497], Fresh[9496], Fresh[9495], Fresh[9494], Fresh[9493], Fresh[9492], Fresh[9491], Fresh[9490], Fresh[9489], Fresh[9488], Fresh[9487], Fresh[9486], Fresh[9485], Fresh[9484], Fresh[9483], Fresh[9482], Fresh[9481], Fresh[9480], Fresh[9479], Fresh[9478], Fresh[9477], Fresh[9476], Fresh[9475], Fresh[9474], Fresh[9473], Fresh[9472], Fresh[9471], Fresh[9470], Fresh[9469], Fresh[9468], Fresh[9467], Fresh[9466], Fresh[9465], Fresh[9464], Fresh[9463], Fresh[9462], Fresh[9461], Fresh[9460], Fresh[9459], Fresh[9458], Fresh[9457], Fresh[9456], Fresh[9455], Fresh[9454], Fresh[9453], Fresh[9452], Fresh[9451], Fresh[9450], Fresh[9449], Fresh[9448], Fresh[9447], Fresh[9446], Fresh[9445], Fresh[9444], Fresh[9443], Fresh[9442], Fresh[9441], Fresh[9440], Fresh[9439], Fresh[9438], Fresh[9437], Fresh[9436], Fresh[9435], Fresh[9434], Fresh[9433], Fresh[9432], Fresh[9431], Fresh[9430], Fresh[9429], Fresh[9428], Fresh[9427], Fresh[9426], Fresh[9425], Fresh[9424], Fresh[9423], Fresh[9422], Fresh[9421], Fresh[9420], Fresh[9419], Fresh[9418], Fresh[9417], Fresh[9416], Fresh[9415], Fresh[9414], Fresh[9413], Fresh[9412], Fresh[9411], Fresh[9410], Fresh[9409], Fresh[9408], Fresh[9407], Fresh[9406], Fresh[9405], Fresh[9404], Fresh[9403], Fresh[9402], Fresh[9401], Fresh[9400], Fresh[9399], Fresh[9398], Fresh[9397], Fresh[9396], Fresh[9395], Fresh[9394], Fresh[9393], Fresh[9392], Fresh[9391], Fresh[9390], Fresh[9389], Fresh[9388], Fresh[9387], Fresh[9386], Fresh[9385], Fresh[9384], Fresh[9383], Fresh[9382], Fresh[9381], Fresh[9380], Fresh[9379], Fresh[9378], Fresh[9377], Fresh[9376], Fresh[9375], Fresh[9374], Fresh[9373], Fresh[9372], Fresh[9371], Fresh[9370], Fresh[9369], Fresh[9368], Fresh[9367], Fresh[9366], Fresh[9365], Fresh[9364], Fresh[9363], Fresh[9362], Fresh[9361], Fresh[9360], Fresh[9359], Fresh[9358], Fresh[9357], Fresh[9356], Fresh[9355], Fresh[9354], Fresh[9353], Fresh[9352], Fresh[9351], Fresh[9350], Fresh[9349], Fresh[9348], Fresh[9347], Fresh[9346], Fresh[9345], Fresh[9344], Fresh[9343], Fresh[9342], Fresh[9341], Fresh[9340], Fresh[9339], Fresh[9338], Fresh[9337], Fresh[9336], Fresh[9335], Fresh[9334], Fresh[9333], Fresh[9332], Fresh[9331], Fresh[9330], Fresh[9329], Fresh[9328], Fresh[9327], Fresh[9326], Fresh[9325], Fresh[9324], Fresh[9323], Fresh[9322], Fresh[9321], Fresh[9320], Fresh[9319], Fresh[9318], Fresh[9317], Fresh[9316], Fresh[9315], Fresh[9314], Fresh[9313], Fresh[9312], Fresh[9311], Fresh[9310], Fresh[9309], Fresh[9308], Fresh[9307], Fresh[9306], Fresh[9305], Fresh[9304], Fresh[9303], Fresh[9302], Fresh[9301], Fresh[9300], Fresh[9299], Fresh[9298], Fresh[9297], Fresh[9296], Fresh[9295], Fresh[9294], Fresh[9293], Fresh[9292], Fresh[9291], Fresh[9290], Fresh[9289], Fresh[9288], Fresh[9287], Fresh[9286], Fresh[9285], Fresh[9284], Fresh[9283], Fresh[9282], Fresh[9281], Fresh[9280], Fresh[9279], Fresh[9278], Fresh[9277], Fresh[9276], Fresh[9275], Fresh[9274], Fresh[9273], Fresh[9272], Fresh[9271], Fresh[9270], Fresh[9269], Fresh[9268], Fresh[9267], Fresh[9266], Fresh[9265], Fresh[9264], Fresh[9263], Fresh[9262], Fresh[9261], Fresh[9260], Fresh[9259], Fresh[9258], Fresh[9257], Fresh[9256], Fresh[9255], Fresh[9254], Fresh[9253], Fresh[9252], Fresh[9251], Fresh[9250], Fresh[9249], Fresh[9248], Fresh[9247], Fresh[9246], Fresh[9245], Fresh[9244], Fresh[9243], Fresh[9242], Fresh[9241], Fresh[9240], Fresh[9239], Fresh[9238], Fresh[9237], Fresh[9236], Fresh[9235], Fresh[9234], Fresh[9233], Fresh[9232], Fresh[9231], Fresh[9230], Fresh[9229], Fresh[9228], Fresh[9227], Fresh[9226], Fresh[9225], Fresh[9224], Fresh[9223], Fresh[9222], Fresh[9221], Fresh[9220], Fresh[9219], Fresh[9218], Fresh[9217], Fresh[9216], Fresh[9215], Fresh[9214], Fresh[9213], Fresh[9212], Fresh[9211], Fresh[9210], Fresh[9209], Fresh[9208], Fresh[9207], Fresh[9206], Fresh[9205], Fresh[9204], Fresh[9203], Fresh[9202], Fresh[9201], Fresh[9200], Fresh[9199], Fresh[9198], Fresh[9197], Fresh[9196], Fresh[9195], Fresh[9194], Fresh[9193], Fresh[9192], Fresh[9191], Fresh[9190], Fresh[9189], Fresh[9188], Fresh[9187], Fresh[9186], Fresh[9185], Fresh[9184], Fresh[9183], Fresh[9182], Fresh[9181], Fresh[9180], Fresh[9179], Fresh[9178], Fresh[9177], Fresh[9176], Fresh[9175], Fresh[9174], Fresh[9173], Fresh[9172], Fresh[9171], Fresh[9170], Fresh[9169], Fresh[9168], Fresh[9167], Fresh[9166], Fresh[9165], Fresh[9164], Fresh[9163], Fresh[9162], Fresh[9161], Fresh[9160], Fresh[9159], Fresh[9158], Fresh[9157], Fresh[9156], Fresh[9155], Fresh[9154], Fresh[9153], Fresh[9152], Fresh[9151], Fresh[9150], Fresh[9149], Fresh[9148], Fresh[9147], Fresh[9146], Fresh[9145], Fresh[9144], Fresh[9143], Fresh[9142], Fresh[9141], Fresh[9140], Fresh[9139], Fresh[9138], Fresh[9137], Fresh[9136], Fresh[9135], Fresh[9134], Fresh[9133], Fresh[9132], Fresh[9131], Fresh[9130], Fresh[9129], Fresh[9128], Fresh[9127], Fresh[9126], Fresh[9125], Fresh[9124], Fresh[9123], Fresh[9122], Fresh[9121], Fresh[9120], Fresh[9119], Fresh[9118], Fresh[9117], Fresh[9116], Fresh[9115], Fresh[9114], Fresh[9113], Fresh[9112], Fresh[9111], Fresh[9110], Fresh[9109], Fresh[9108], Fresh[9107], Fresh[9106], Fresh[9105], Fresh[9104], Fresh[9103], Fresh[9102], Fresh[9101], Fresh[9100], Fresh[9099], Fresh[9098], Fresh[9097], Fresh[9096], Fresh[9095], Fresh[9094], Fresh[9093], Fresh[9092], Fresh[9091], Fresh[9090], Fresh[9089], Fresh[9088], Fresh[9087], Fresh[9086], Fresh[9085], Fresh[9084], Fresh[9083], Fresh[9082], Fresh[9081], Fresh[9080], Fresh[9079], Fresh[9078], Fresh[9077], Fresh[9076], Fresh[9075], Fresh[9074], Fresh[9073], Fresh[9072], Fresh[9071], Fresh[9070], Fresh[9069], Fresh[9068], Fresh[9067], Fresh[9066], Fresh[9065], Fresh[9064], Fresh[9063], Fresh[9062], Fresh[9061], Fresh[9060], Fresh[9059], Fresh[9058], Fresh[9057], Fresh[9056], Fresh[9055], Fresh[9054], Fresh[9053], Fresh[9052], Fresh[9051], Fresh[9050], Fresh[9049], Fresh[9048], Fresh[9047], Fresh[9046], Fresh[9045], Fresh[9044], Fresh[9043], Fresh[9042], Fresh[9041], Fresh[9040], Fresh[9039], Fresh[9038], Fresh[9037], Fresh[9036], Fresh[9035], Fresh[9034], Fresh[9033], Fresh[9032], Fresh[9031], Fresh[9030], Fresh[9029], Fresh[9028], Fresh[9027], Fresh[9026], Fresh[9025], Fresh[9024], Fresh[9023], Fresh[9022], Fresh[9021], Fresh[9020], Fresh[9019], Fresh[9018], Fresh[9017], Fresh[9016], Fresh[9015], Fresh[9014], Fresh[9013], Fresh[9012], Fresh[9011], Fresh[9010], Fresh[9009], Fresh[9008], Fresh[9007], Fresh[9006], Fresh[9005], Fresh[9004], Fresh[9003], Fresh[9002], Fresh[9001], Fresh[9000], Fresh[8999], Fresh[8998], Fresh[8997], Fresh[8996], Fresh[8995], Fresh[8994], Fresh[8993], Fresh[8992], Fresh[8991], Fresh[8990], Fresh[8989], Fresh[8988], Fresh[8987], Fresh[8986], Fresh[8985], Fresh[8984], Fresh[8983], Fresh[8982], Fresh[8981], Fresh[8980], Fresh[8979], Fresh[8978], Fresh[8977], Fresh[8976], Fresh[8975], Fresh[8974], Fresh[8973], Fresh[8972], Fresh[8971], Fresh[8970], Fresh[8969], Fresh[8968], Fresh[8967], Fresh[8966], Fresh[8965], Fresh[8964], Fresh[8963], Fresh[8962], Fresh[8961], Fresh[8960], Fresh[8959], Fresh[8958], Fresh[8957], Fresh[8956], Fresh[8955], Fresh[8954], Fresh[8953], Fresh[8952], Fresh[8951], Fresh[8950], Fresh[8949], Fresh[8948], Fresh[8947], Fresh[8946], Fresh[8945], Fresh[8944], Fresh[8943], Fresh[8942], Fresh[8941], Fresh[8940], Fresh[8939], Fresh[8938], Fresh[8937], Fresh[8936], Fresh[8935], Fresh[8934], Fresh[8933], Fresh[8932], Fresh[8931], Fresh[8930], Fresh[8929], Fresh[8928], Fresh[8927], Fresh[8926], Fresh[8925], Fresh[8924], Fresh[8923], Fresh[8922], Fresh[8921], Fresh[8920], Fresh[8919], Fresh[8918], Fresh[8917], Fresh[8916], Fresh[8915], Fresh[8914], Fresh[8913], Fresh[8912], Fresh[8911], Fresh[8910], Fresh[8909], Fresh[8908], Fresh[8907], Fresh[8906], Fresh[8905], Fresh[8904], Fresh[8903], Fresh[8902], Fresh[8901], Fresh[8900], Fresh[8899], Fresh[8898], Fresh[8897], Fresh[8896], Fresh[8895], Fresh[8894], Fresh[8893], Fresh[8892], Fresh[8891], Fresh[8890], Fresh[8889], Fresh[8888], Fresh[8887], Fresh[8886], Fresh[8885], Fresh[8884], Fresh[8883], Fresh[8882], Fresh[8881], Fresh[8880], Fresh[8879], Fresh[8878], Fresh[8877], Fresh[8876], Fresh[8875], Fresh[8874], Fresh[8873], Fresh[8872], Fresh[8871], Fresh[8870], Fresh[8869], Fresh[8868], Fresh[8867], Fresh[8866], Fresh[8865], Fresh[8864], Fresh[8863], Fresh[8862], Fresh[8861], Fresh[8860], Fresh[8859], Fresh[8858], Fresh[8857], Fresh[8856], Fresh[8855], Fresh[8854], Fresh[8853], Fresh[8852], Fresh[8851], Fresh[8850], Fresh[8849], Fresh[8848], Fresh[8847], Fresh[8846], Fresh[8845], Fresh[8844], Fresh[8843], Fresh[8842], Fresh[8841], Fresh[8840], Fresh[8839], Fresh[8838], Fresh[8837], Fresh[8836], Fresh[8835], Fresh[8834], Fresh[8833], Fresh[8832], Fresh[8831], Fresh[8830], Fresh[8829], Fresh[8828], Fresh[8827], Fresh[8826], Fresh[8825], Fresh[8824], Fresh[8823], Fresh[8822], Fresh[8821], Fresh[8820], Fresh[8819], Fresh[8818], Fresh[8817], Fresh[8816], Fresh[8815], Fresh[8814], Fresh[8813], Fresh[8812], Fresh[8811], Fresh[8810], Fresh[8809], Fresh[8808], Fresh[8807], Fresh[8806], Fresh[8805], Fresh[8804], Fresh[8803], Fresh[8802], Fresh[8801], Fresh[8800], Fresh[8799], Fresh[8798], Fresh[8797], Fresh[8796], Fresh[8795], Fresh[8794], Fresh[8793], Fresh[8792], Fresh[8791], Fresh[8790], Fresh[8789], Fresh[8788], Fresh[8787], Fresh[8786], Fresh[8785], Fresh[8784], Fresh[8783], Fresh[8782], Fresh[8781], Fresh[8780], Fresh[8779], Fresh[8778], Fresh[8777], Fresh[8776], Fresh[8775], Fresh[8774], Fresh[8773], Fresh[8772], Fresh[8771], Fresh[8770], Fresh[8769], Fresh[8768], Fresh[8767], Fresh[8766], Fresh[8765], Fresh[8764], Fresh[8763], Fresh[8762], Fresh[8761], Fresh[8760], Fresh[8759], Fresh[8758], Fresh[8757], Fresh[8756], Fresh[8755], Fresh[8754], Fresh[8753], Fresh[8752], Fresh[8751], Fresh[8750], Fresh[8749], Fresh[8748], Fresh[8747], Fresh[8746], Fresh[8745], Fresh[8744], Fresh[8743], Fresh[8742], Fresh[8741], Fresh[8740], Fresh[8739], Fresh[8738], Fresh[8737], Fresh[8736], Fresh[8735], Fresh[8734], Fresh[8733], Fresh[8732], Fresh[8731], Fresh[8730], Fresh[8729], Fresh[8728], Fresh[8727], Fresh[8726], Fresh[8725], Fresh[8724], Fresh[8723], Fresh[8722], Fresh[8721], Fresh[8720], Fresh[8719], Fresh[8718], Fresh[8717], Fresh[8716], Fresh[8715], Fresh[8714], Fresh[8713], Fresh[8712], Fresh[8711], Fresh[8710], Fresh[8709], Fresh[8708], Fresh[8707], Fresh[8706], Fresh[8705], Fresh[8704], Fresh[8703], Fresh[8702], Fresh[8701], Fresh[8700], Fresh[8699], Fresh[8698], Fresh[8697], Fresh[8696], Fresh[8695], Fresh[8694], Fresh[8693], Fresh[8692], Fresh[8691], Fresh[8690], Fresh[8689], Fresh[8688], Fresh[8687], Fresh[8686], Fresh[8685], Fresh[8684], Fresh[8683], Fresh[8682], Fresh[8681], Fresh[8680], Fresh[8679], Fresh[8678], Fresh[8677], Fresh[8676], Fresh[8675], Fresh[8674], Fresh[8673], Fresh[8672], Fresh[8671], Fresh[8670], Fresh[8669], Fresh[8668], Fresh[8667], Fresh[8666], Fresh[8665], Fresh[8664], Fresh[8663], Fresh[8662], Fresh[8661], Fresh[8660], Fresh[8659], Fresh[8658], Fresh[8657], Fresh[8656], Fresh[8655], Fresh[8654], Fresh[8653], Fresh[8652], Fresh[8651], Fresh[8650], Fresh[8649], Fresh[8648], Fresh[8647], Fresh[8646], Fresh[8645], Fresh[8644], Fresh[8643], Fresh[8642], Fresh[8641], Fresh[8640], Fresh[8639], Fresh[8638], Fresh[8637], Fresh[8636], Fresh[8635], Fresh[8634], Fresh[8633], Fresh[8632], Fresh[8631], Fresh[8630], Fresh[8629], Fresh[8628], Fresh[8627], Fresh[8626], Fresh[8625], Fresh[8624], Fresh[8623], Fresh[8622], Fresh[8621], Fresh[8620], Fresh[8619], Fresh[8618], Fresh[8617], Fresh[8616], Fresh[8615], Fresh[8614], Fresh[8613], Fresh[8612], Fresh[8611], Fresh[8610], Fresh[8609], Fresh[8608], Fresh[8607], Fresh[8606], Fresh[8605], Fresh[8604], Fresh[8603], Fresh[8602], Fresh[8601], Fresh[8600], Fresh[8599], Fresh[8598], Fresh[8597], Fresh[8596], Fresh[8595], Fresh[8594], Fresh[8593], Fresh[8592], Fresh[8591], Fresh[8590], Fresh[8589], Fresh[8588], Fresh[8587], Fresh[8586], Fresh[8585], Fresh[8584], Fresh[8583], Fresh[8582], Fresh[8581], Fresh[8580], Fresh[8579], Fresh[8578], Fresh[8577], Fresh[8576], Fresh[8575], Fresh[8574], Fresh[8573], Fresh[8572], Fresh[8571], Fresh[8570], Fresh[8569], Fresh[8568], Fresh[8567], Fresh[8566], Fresh[8565], Fresh[8564], Fresh[8563], Fresh[8562], Fresh[8561], Fresh[8560], Fresh[8559], Fresh[8558], Fresh[8557], Fresh[8556], Fresh[8555], Fresh[8554], Fresh[8553], Fresh[8552], Fresh[8551], Fresh[8550], Fresh[8549], Fresh[8548], Fresh[8547], Fresh[8546], Fresh[8545], Fresh[8544], Fresh[8543], Fresh[8542], Fresh[8541], Fresh[8540], Fresh[8539], Fresh[8538], Fresh[8537], Fresh[8536], Fresh[8535], Fresh[8534], Fresh[8533], Fresh[8532], Fresh[8531], Fresh[8530], Fresh[8529], Fresh[8528], Fresh[8527], Fresh[8526], Fresh[8525], Fresh[8524], Fresh[8523], Fresh[8522], Fresh[8521], Fresh[8520], Fresh[8519], Fresh[8518], Fresh[8517], Fresh[8516], Fresh[8515], Fresh[8514], Fresh[8513], Fresh[8512], Fresh[8511], Fresh[8510], Fresh[8509], Fresh[8508], Fresh[8507], Fresh[8506], Fresh[8505], Fresh[8504], Fresh[8503], Fresh[8502], Fresh[8501], Fresh[8500], Fresh[8499], Fresh[8498], Fresh[8497], Fresh[8496], Fresh[8495], Fresh[8494], Fresh[8493], Fresh[8492], Fresh[8491], Fresh[8490], Fresh[8489], Fresh[8488], Fresh[8487], Fresh[8486], Fresh[8485], Fresh[8484], Fresh[8483], Fresh[8482], Fresh[8481], Fresh[8480], Fresh[8479], Fresh[8478], Fresh[8477], Fresh[8476], Fresh[8475], Fresh[8474], Fresh[8473], Fresh[8472], Fresh[8471], Fresh[8470], Fresh[8469], Fresh[8468], Fresh[8467], Fresh[8466], Fresh[8465], Fresh[8464], Fresh[8463], Fresh[8462], Fresh[8461], Fresh[8460], Fresh[8459], Fresh[8458], Fresh[8457], Fresh[8456], Fresh[8455], Fresh[8454], Fresh[8453], Fresh[8452], Fresh[8451], Fresh[8450], Fresh[8449], Fresh[8448], Fresh[8447], Fresh[8446], Fresh[8445], Fresh[8444], Fresh[8443], Fresh[8442], Fresh[8441], Fresh[8440], Fresh[8439], Fresh[8438], Fresh[8437], Fresh[8436], Fresh[8435], Fresh[8434], Fresh[8433], Fresh[8432], Fresh[8431], Fresh[8430], Fresh[8429], Fresh[8428], Fresh[8427], Fresh[8426], Fresh[8425], Fresh[8424], Fresh[8423], Fresh[8422], Fresh[8421], Fresh[8420], Fresh[8419], Fresh[8418], Fresh[8417], Fresh[8416], Fresh[8415], Fresh[8414], Fresh[8413], Fresh[8412], Fresh[8411], Fresh[8410], Fresh[8409], Fresh[8408], Fresh[8407], Fresh[8406], Fresh[8405], Fresh[8404], Fresh[8403], Fresh[8402], Fresh[8401], Fresh[8400], Fresh[8399], Fresh[8398], Fresh[8397], Fresh[8396], Fresh[8395], Fresh[8394], Fresh[8393], Fresh[8392], Fresh[8391], Fresh[8390], Fresh[8389], Fresh[8388], Fresh[8387], Fresh[8386], Fresh[8385], Fresh[8384], Fresh[8383], Fresh[8382], Fresh[8381], Fresh[8380], Fresh[8379], Fresh[8378], Fresh[8377], Fresh[8376], Fresh[8375], Fresh[8374], Fresh[8373], Fresh[8372], Fresh[8371], Fresh[8370], Fresh[8369], Fresh[8368], Fresh[8367], Fresh[8366], Fresh[8365], Fresh[8364], Fresh[8363], Fresh[8362], Fresh[8361], Fresh[8360], Fresh[8359], Fresh[8358], Fresh[8357], Fresh[8356], Fresh[8355], Fresh[8354], Fresh[8353], Fresh[8352], Fresh[8351], Fresh[8350], Fresh[8349], Fresh[8348], Fresh[8347], Fresh[8346], Fresh[8345], Fresh[8344], Fresh[8343], Fresh[8342], Fresh[8341], Fresh[8340], Fresh[8339], Fresh[8338], Fresh[8337], Fresh[8336], Fresh[8335], Fresh[8334], Fresh[8333], Fresh[8332], Fresh[8331], Fresh[8330], Fresh[8329], Fresh[8328], Fresh[8327], Fresh[8326], Fresh[8325], Fresh[8324], Fresh[8323], Fresh[8322], Fresh[8321], Fresh[8320], Fresh[8319], Fresh[8318], Fresh[8317], Fresh[8316], Fresh[8315], Fresh[8314], Fresh[8313], Fresh[8312], Fresh[8311], Fresh[8310], Fresh[8309], Fresh[8308], Fresh[8307], Fresh[8306], Fresh[8305], Fresh[8304], Fresh[8303], Fresh[8302], Fresh[8301], Fresh[8300], Fresh[8299], Fresh[8298], Fresh[8297], Fresh[8296], Fresh[8295], Fresh[8294], Fresh[8293], Fresh[8292], Fresh[8291], Fresh[8290], Fresh[8289], Fresh[8288], Fresh[8287], Fresh[8286], Fresh[8285], Fresh[8284], Fresh[8283], Fresh[8282], Fresh[8281], Fresh[8280], Fresh[8279], Fresh[8278], Fresh[8277], Fresh[8276], Fresh[8275], Fresh[8274], Fresh[8273], Fresh[8272], Fresh[8271], Fresh[8270], Fresh[8269], Fresh[8268], Fresh[8267], Fresh[8266], Fresh[8265], Fresh[8264], Fresh[8263], Fresh[8262], Fresh[8261], Fresh[8260], Fresh[8259], Fresh[8258], Fresh[8257], Fresh[8256], Fresh[8255], Fresh[8254], Fresh[8253], Fresh[8252], Fresh[8251], Fresh[8250], Fresh[8249], Fresh[8248], Fresh[8247], Fresh[8246], Fresh[8245], Fresh[8244], Fresh[8243], Fresh[8242], Fresh[8241], Fresh[8240], Fresh[8239], Fresh[8238], Fresh[8237], Fresh[8236], Fresh[8235], Fresh[8234], Fresh[8233], Fresh[8232], Fresh[8231], Fresh[8230], Fresh[8229], Fresh[8228], Fresh[8227], Fresh[8226], Fresh[8225], Fresh[8224], Fresh[8223], Fresh[8222], Fresh[8221], Fresh[8220], Fresh[8219], Fresh[8218], Fresh[8217], Fresh[8216], Fresh[8215], Fresh[8214], Fresh[8213], Fresh[8212], Fresh[8211], Fresh[8210], Fresh[8209], Fresh[8208], Fresh[8207], Fresh[8206], Fresh[8205], Fresh[8204], Fresh[8203], Fresh[8202], Fresh[8201], Fresh[8200], Fresh[8199], Fresh[8198], Fresh[8197], Fresh[8196], Fresh[8195], Fresh[8194], Fresh[8193], Fresh[8192], Fresh[8191], Fresh[8190], Fresh[8189], Fresh[8188], Fresh[8187], Fresh[8186], Fresh[8185], Fresh[8184], Fresh[8183], Fresh[8182], Fresh[8181], Fresh[8180], Fresh[8179], Fresh[8178], Fresh[8177], Fresh[8176], Fresh[8175], Fresh[8174], Fresh[8173], Fresh[8172], Fresh[8171], Fresh[8170], Fresh[8169], Fresh[8168], Fresh[8167], Fresh[8166], Fresh[8165], Fresh[8164], Fresh[8163], Fresh[8162], Fresh[8161], Fresh[8160], Fresh[8159], Fresh[8158], Fresh[8157], Fresh[8156], Fresh[8155], Fresh[8154], Fresh[8153], Fresh[8152], Fresh[8151], Fresh[8150], Fresh[8149], Fresh[8148], Fresh[8147], Fresh[8146], Fresh[8145], Fresh[8144], Fresh[8143], Fresh[8142], Fresh[8141], Fresh[8140], Fresh[8139], Fresh[8138], Fresh[8137], Fresh[8136], Fresh[8135], Fresh[8134], Fresh[8133], Fresh[8132], Fresh[8131], Fresh[8130], Fresh[8129], Fresh[8128], Fresh[8127], Fresh[8126], Fresh[8125], Fresh[8124], Fresh[8123], Fresh[8122], Fresh[8121], Fresh[8120], Fresh[8119], Fresh[8118], Fresh[8117], Fresh[8116], Fresh[8115], Fresh[8114], Fresh[8113], Fresh[8112], Fresh[8111], Fresh[8110], Fresh[8109], Fresh[8108], Fresh[8107], Fresh[8106], Fresh[8105], Fresh[8104], Fresh[8103], Fresh[8102], Fresh[8101], Fresh[8100], Fresh[8099], Fresh[8098], Fresh[8097], Fresh[8096], Fresh[8095], Fresh[8094], Fresh[8093], Fresh[8092], Fresh[8091], Fresh[8090], Fresh[8089], Fresh[8088], Fresh[8087], Fresh[8086], Fresh[8085], Fresh[8084], Fresh[8083], Fresh[8082], Fresh[8081], Fresh[8080], Fresh[8079], Fresh[8078], Fresh[8077], Fresh[8076], Fresh[8075], Fresh[8074], Fresh[8073], Fresh[8072], Fresh[8071], Fresh[8070], Fresh[8069], Fresh[8068], Fresh[8067], Fresh[8066], Fresh[8065], Fresh[8064], Fresh[8063], Fresh[8062], Fresh[8061], Fresh[8060], Fresh[8059], Fresh[8058], Fresh[8057], Fresh[8056], Fresh[8055], Fresh[8054], Fresh[8053], Fresh[8052], Fresh[8051], Fresh[8050], Fresh[8049], Fresh[8048], Fresh[8047], Fresh[8046], Fresh[8045], Fresh[8044], Fresh[8043], Fresh[8042], Fresh[8041], Fresh[8040], Fresh[8039], Fresh[8038], Fresh[8037], Fresh[8036], Fresh[8035], Fresh[8034], Fresh[8033], Fresh[8032], Fresh[8031], Fresh[8030], Fresh[8029], Fresh[8028], Fresh[8027], Fresh[8026], Fresh[8025], Fresh[8024], Fresh[8023], Fresh[8022], Fresh[8021], Fresh[8020], Fresh[8019], Fresh[8018], Fresh[8017], Fresh[8016], Fresh[8015], Fresh[8014], Fresh[8013], Fresh[8012], Fresh[8011], Fresh[8010], Fresh[8009], Fresh[8008], Fresh[8007], Fresh[8006], Fresh[8005], Fresh[8004], Fresh[8003], Fresh[8002], Fresh[8001], Fresh[8000], Fresh[7999], Fresh[7998], Fresh[7997], Fresh[7996], Fresh[7995], Fresh[7994], Fresh[7993], Fresh[7992], Fresh[7991], Fresh[7990], Fresh[7989], Fresh[7988], Fresh[7987], Fresh[7986], Fresh[7985], Fresh[7984], Fresh[7983], Fresh[7982], Fresh[7981], Fresh[7980], Fresh[7979], Fresh[7978], Fresh[7977], Fresh[7976], Fresh[7975], Fresh[7974], Fresh[7973], Fresh[7972], Fresh[7971], Fresh[7970], Fresh[7969], Fresh[7968], Fresh[7967], Fresh[7966], Fresh[7965], Fresh[7964], Fresh[7963], Fresh[7962], Fresh[7961], Fresh[7960], Fresh[7959], Fresh[7958], Fresh[7957], Fresh[7956], Fresh[7955], Fresh[7954], Fresh[7953], Fresh[7952], Fresh[7951], Fresh[7950], Fresh[7949], Fresh[7948], Fresh[7947], Fresh[7946], Fresh[7945], Fresh[7944], Fresh[7943], Fresh[7942], Fresh[7941], Fresh[7940], Fresh[7939], Fresh[7938], Fresh[7937], Fresh[7936], Fresh[7935], Fresh[7934], Fresh[7933], Fresh[7932], Fresh[7931], Fresh[7930], Fresh[7929], Fresh[7928], Fresh[7927], Fresh[7926], Fresh[7925], Fresh[7924], Fresh[7923], Fresh[7922], Fresh[7921], Fresh[7920], Fresh[7919], Fresh[7918], Fresh[7917], Fresh[7916], Fresh[7915], Fresh[7914], Fresh[7913], Fresh[7912], Fresh[7911], Fresh[7910], Fresh[7909], Fresh[7908], Fresh[7907], Fresh[7906], Fresh[7905], Fresh[7904], Fresh[7903], Fresh[7902], Fresh[7901], Fresh[7900], Fresh[7899], Fresh[7898], Fresh[7897], Fresh[7896], Fresh[7895], Fresh[7894], Fresh[7893], Fresh[7892], Fresh[7891], Fresh[7890], Fresh[7889], Fresh[7888], Fresh[7887], Fresh[7886], Fresh[7885], Fresh[7884], Fresh[7883], Fresh[7882], Fresh[7881], Fresh[7880], Fresh[7879], Fresh[7878], Fresh[7877], Fresh[7876], Fresh[7875], Fresh[7874], Fresh[7873], Fresh[7872], Fresh[7871], Fresh[7870], Fresh[7869], Fresh[7868], Fresh[7867], Fresh[7866], Fresh[7865], Fresh[7864], Fresh[7863], Fresh[7862], Fresh[7861], Fresh[7860], Fresh[7859], Fresh[7858], Fresh[7857], Fresh[7856], Fresh[7855], Fresh[7854], Fresh[7853], Fresh[7852], Fresh[7851], Fresh[7850], Fresh[7849], Fresh[7848], Fresh[7847], Fresh[7846], Fresh[7845], Fresh[7844], Fresh[7843], Fresh[7842], Fresh[7841], Fresh[7840], Fresh[7839], Fresh[7838], Fresh[7837], Fresh[7836], Fresh[7835], Fresh[7834], Fresh[7833], Fresh[7832], Fresh[7831], Fresh[7830], Fresh[7829], Fresh[7828], Fresh[7827], Fresh[7826], Fresh[7825], Fresh[7824], Fresh[7823], Fresh[7822], Fresh[7821], Fresh[7820], Fresh[7819], Fresh[7818], Fresh[7817], Fresh[7816], Fresh[7815], Fresh[7814], Fresh[7813], Fresh[7812], Fresh[7811], Fresh[7810], Fresh[7809], Fresh[7808], Fresh[7807], Fresh[7806], Fresh[7805], Fresh[7804], Fresh[7803], Fresh[7802], Fresh[7801], Fresh[7800], Fresh[7799], Fresh[7798], Fresh[7797], Fresh[7796], Fresh[7795], Fresh[7794], Fresh[7793], Fresh[7792], Fresh[7791], Fresh[7790], Fresh[7789], Fresh[7788], Fresh[7787], Fresh[7786], Fresh[7785], Fresh[7784], Fresh[7783], Fresh[7782], Fresh[7781], Fresh[7780], Fresh[7779], Fresh[7778], Fresh[7777], Fresh[7776], Fresh[7775], Fresh[7774], Fresh[7773], Fresh[7772], Fresh[7771], Fresh[7770], Fresh[7769], Fresh[7768], Fresh[7767], Fresh[7766], Fresh[7765], Fresh[7764], Fresh[7763], Fresh[7762], Fresh[7761], Fresh[7760], Fresh[7759], Fresh[7758], Fresh[7757], Fresh[7756], Fresh[7755], Fresh[7754], Fresh[7753], Fresh[7752], Fresh[7751], Fresh[7750], Fresh[7749], Fresh[7748], Fresh[7747], Fresh[7746], Fresh[7745], Fresh[7744], Fresh[7743], Fresh[7742], Fresh[7741], Fresh[7740], Fresh[7739], Fresh[7738], Fresh[7737], Fresh[7736], Fresh[7735], Fresh[7734], Fresh[7733], Fresh[7732], Fresh[7731], Fresh[7730], Fresh[7729], Fresh[7728], Fresh[7727], Fresh[7726], Fresh[7725], Fresh[7724], Fresh[7723], Fresh[7722], Fresh[7721], Fresh[7720], Fresh[7719], Fresh[7718], Fresh[7717], Fresh[7716], Fresh[7715], Fresh[7714], Fresh[7713], Fresh[7712], Fresh[7711], Fresh[7710], Fresh[7709], Fresh[7708], Fresh[7707], Fresh[7706], Fresh[7705], Fresh[7704], Fresh[7703], Fresh[7702], Fresh[7701], Fresh[7700], Fresh[7699], Fresh[7698], Fresh[7697], Fresh[7696], Fresh[7695], Fresh[7694], Fresh[7693], Fresh[7692], Fresh[7691], Fresh[7690], Fresh[7689], Fresh[7688], Fresh[7687], Fresh[7686], Fresh[7685], Fresh[7684], Fresh[7683], Fresh[7682], Fresh[7681], Fresh[7680], Fresh[7679], Fresh[7678], Fresh[7677], Fresh[7676], Fresh[7675], Fresh[7674], Fresh[7673], Fresh[7672], Fresh[7671], Fresh[7670], Fresh[7669], Fresh[7668], Fresh[7667], Fresh[7666], Fresh[7665], Fresh[7664], Fresh[7663], Fresh[7662], Fresh[7661], Fresh[7660], Fresh[7659], Fresh[7658], Fresh[7657], Fresh[7656], Fresh[7655], Fresh[7654], Fresh[7653], Fresh[7652], Fresh[7651], Fresh[7650], Fresh[7649], Fresh[7648], Fresh[7647], Fresh[7646], Fresh[7645], Fresh[7644], Fresh[7643], Fresh[7642], Fresh[7641], Fresh[7640], Fresh[7639], Fresh[7638], Fresh[7637], Fresh[7636], Fresh[7635], Fresh[7634], Fresh[7633], Fresh[7632], Fresh[7631], Fresh[7630], Fresh[7629], Fresh[7628], Fresh[7627], Fresh[7626], Fresh[7625], Fresh[7624], Fresh[7623], Fresh[7622], Fresh[7621], Fresh[7620], Fresh[7619], Fresh[7618], Fresh[7617], Fresh[7616], Fresh[7615], Fresh[7614], Fresh[7613], Fresh[7612], Fresh[7611], Fresh[7610], Fresh[7609], Fresh[7608], Fresh[7607], Fresh[7606], Fresh[7605], Fresh[7604], Fresh[7603], Fresh[7602], Fresh[7601], Fresh[7600], Fresh[7599], Fresh[7598], Fresh[7597], Fresh[7596], Fresh[7595], Fresh[7594], Fresh[7593], Fresh[7592], Fresh[7591], Fresh[7590], Fresh[7589], Fresh[7588], Fresh[7587], Fresh[7586], Fresh[7585], Fresh[7584], Fresh[7583], Fresh[7582], Fresh[7581], Fresh[7580], Fresh[7579], Fresh[7578], Fresh[7577], Fresh[7576], Fresh[7575], Fresh[7574], Fresh[7573], Fresh[7572], Fresh[7571], Fresh[7570], Fresh[7569], Fresh[7568], Fresh[7567], Fresh[7566], Fresh[7565], Fresh[7564], Fresh[7563], Fresh[7562], Fresh[7561], Fresh[7560], Fresh[7559], Fresh[7558], Fresh[7557], Fresh[7556], Fresh[7555], Fresh[7554], Fresh[7553], Fresh[7552], Fresh[7551], Fresh[7550], Fresh[7549], Fresh[7548], Fresh[7547], Fresh[7546], Fresh[7545], Fresh[7544], Fresh[7543], Fresh[7542], Fresh[7541], Fresh[7540], Fresh[7539], Fresh[7538], Fresh[7537], Fresh[7536], Fresh[7535], Fresh[7534], Fresh[7533], Fresh[7532], Fresh[7531], Fresh[7530], Fresh[7529], Fresh[7528], Fresh[7527], Fresh[7526], Fresh[7525], Fresh[7524], Fresh[7523], Fresh[7522], Fresh[7521], Fresh[7520], Fresh[7519], Fresh[7518], Fresh[7517], Fresh[7516], Fresh[7515], Fresh[7514], Fresh[7513], Fresh[7512], Fresh[7511], Fresh[7510], Fresh[7509], Fresh[7508], Fresh[7507], Fresh[7506], Fresh[7505], Fresh[7504], Fresh[7503], Fresh[7502], Fresh[7501], Fresh[7500], Fresh[7499], Fresh[7498], Fresh[7497], Fresh[7496], Fresh[7495], Fresh[7494], Fresh[7493], Fresh[7492], Fresh[7491], Fresh[7490], Fresh[7489], Fresh[7488], Fresh[7487], Fresh[7486], Fresh[7485], Fresh[7484], Fresh[7483], Fresh[7482], Fresh[7481], Fresh[7480], Fresh[7479], Fresh[7478], Fresh[7477], Fresh[7476], Fresh[7475], Fresh[7474], Fresh[7473], Fresh[7472], Fresh[7471], Fresh[7470], Fresh[7469], Fresh[7468], Fresh[7467], Fresh[7466], Fresh[7465], Fresh[7464], Fresh[7463], Fresh[7462], Fresh[7461], Fresh[7460], Fresh[7459], Fresh[7458], Fresh[7457], Fresh[7456], Fresh[7455], Fresh[7454], Fresh[7453], Fresh[7452], Fresh[7451], Fresh[7450], Fresh[7449], Fresh[7448], Fresh[7447], Fresh[7446], Fresh[7445], Fresh[7444], Fresh[7443], Fresh[7442], Fresh[7441], Fresh[7440], Fresh[7439], Fresh[7438], Fresh[7437], Fresh[7436], Fresh[7435], Fresh[7434], Fresh[7433], Fresh[7432], Fresh[7431], Fresh[7430], Fresh[7429], Fresh[7428], Fresh[7427], Fresh[7426], Fresh[7425], Fresh[7424], Fresh[7423], Fresh[7422], Fresh[7421], Fresh[7420], Fresh[7419], Fresh[7418], Fresh[7417], Fresh[7416], Fresh[7415], Fresh[7414], Fresh[7413], Fresh[7412], Fresh[7411], Fresh[7410], Fresh[7409], Fresh[7408], Fresh[7407], Fresh[7406], Fresh[7405], Fresh[7404], Fresh[7403], Fresh[7402], Fresh[7401], Fresh[7400], Fresh[7399], Fresh[7398], Fresh[7397], Fresh[7396], Fresh[7395], Fresh[7394], Fresh[7393], Fresh[7392], Fresh[7391], Fresh[7390], Fresh[7389], Fresh[7388], Fresh[7387], Fresh[7386], Fresh[7385], Fresh[7384], Fresh[7383], Fresh[7382], Fresh[7381], Fresh[7380], Fresh[7379], Fresh[7378], Fresh[7377], Fresh[7376], Fresh[7375], Fresh[7374], Fresh[7373], Fresh[7372], Fresh[7371], Fresh[7370], Fresh[7369], Fresh[7368], Fresh[7367], Fresh[7366], Fresh[7365], Fresh[7364], Fresh[7363], Fresh[7362], Fresh[7361], Fresh[7360], Fresh[7359], Fresh[7358], Fresh[7357], Fresh[7356], Fresh[7355], Fresh[7354], Fresh[7353], Fresh[7352], Fresh[7351], Fresh[7350], Fresh[7349], Fresh[7348], Fresh[7347], Fresh[7346], Fresh[7345], Fresh[7344], Fresh[7343], Fresh[7342], Fresh[7341], Fresh[7340], Fresh[7339], Fresh[7338], Fresh[7337], Fresh[7336], Fresh[7335], Fresh[7334], Fresh[7333], Fresh[7332], Fresh[7331], Fresh[7330], Fresh[7329], Fresh[7328], Fresh[7327], Fresh[7326], Fresh[7325], Fresh[7324], Fresh[7323], Fresh[7322], Fresh[7321], Fresh[7320], Fresh[7319], Fresh[7318], Fresh[7317], Fresh[7316], Fresh[7315], Fresh[7314], Fresh[7313], Fresh[7312], Fresh[7311], Fresh[7310], Fresh[7309], Fresh[7308], Fresh[7307], Fresh[7306], Fresh[7305], Fresh[7304], Fresh[7303], Fresh[7302], Fresh[7301], Fresh[7300], Fresh[7299], Fresh[7298], Fresh[7297], Fresh[7296], Fresh[7295], Fresh[7294], Fresh[7293], Fresh[7292], Fresh[7291], Fresh[7290], Fresh[7289], Fresh[7288], Fresh[7287], Fresh[7286], Fresh[7285], Fresh[7284], Fresh[7283], Fresh[7282], Fresh[7281], Fresh[7280], Fresh[7279], Fresh[7278], Fresh[7277], Fresh[7276], Fresh[7275], Fresh[7274], Fresh[7273], Fresh[7272], Fresh[7271], Fresh[7270], Fresh[7269], Fresh[7268], Fresh[7267], Fresh[7266], Fresh[7265], Fresh[7264], Fresh[7263], Fresh[7262], Fresh[7261], Fresh[7260], Fresh[7259], Fresh[7258], Fresh[7257], Fresh[7256], Fresh[7255], Fresh[7254], Fresh[7253], Fresh[7252], Fresh[7251], Fresh[7250], Fresh[7249], Fresh[7248], Fresh[7247], Fresh[7246], Fresh[7245], Fresh[7244], Fresh[7243], Fresh[7242], Fresh[7241], Fresh[7240], Fresh[7239], Fresh[7238], Fresh[7237], Fresh[7236], Fresh[7235], Fresh[7234], Fresh[7233], Fresh[7232], Fresh[7231], Fresh[7230], Fresh[7229], Fresh[7228], Fresh[7227], Fresh[7226], Fresh[7225], Fresh[7224], Fresh[7223], Fresh[7222], Fresh[7221], Fresh[7220], Fresh[7219], Fresh[7218], Fresh[7217], Fresh[7216], Fresh[7215], Fresh[7214], Fresh[7213], Fresh[7212], Fresh[7211], Fresh[7210], Fresh[7209], Fresh[7208], Fresh[7207], Fresh[7206], Fresh[7205], Fresh[7204], Fresh[7203], Fresh[7202], Fresh[7201], Fresh[7200], Fresh[7199], Fresh[7198], Fresh[7197], Fresh[7196], Fresh[7195], Fresh[7194], Fresh[7193], Fresh[7192], Fresh[7191], Fresh[7190], Fresh[7189], Fresh[7188], Fresh[7187], Fresh[7186], Fresh[7185], Fresh[7184], Fresh[7183], Fresh[7182], Fresh[7181], Fresh[7180], Fresh[7179], Fresh[7178], Fresh[7177], Fresh[7176], Fresh[7175], Fresh[7174], Fresh[7173], Fresh[7172], Fresh[7171], Fresh[7170], Fresh[7169], Fresh[7168], Fresh[7167], Fresh[7166], Fresh[7165], Fresh[7164], Fresh[7163], Fresh[7162], Fresh[7161], Fresh[7160], Fresh[7159], Fresh[7158], Fresh[7157], Fresh[7156], Fresh[7155], Fresh[7154], Fresh[7153], Fresh[7152], Fresh[7151], Fresh[7150], Fresh[7149], Fresh[7148], Fresh[7147], Fresh[7146], Fresh[7145], Fresh[7144], Fresh[7143], Fresh[7142], Fresh[7141], Fresh[7140], Fresh[7139], Fresh[7138], Fresh[7137], Fresh[7136], Fresh[7135], Fresh[7134], Fresh[7133], Fresh[7132], Fresh[7131], Fresh[7130], Fresh[7129], Fresh[7128], Fresh[7127], Fresh[7126], Fresh[7125], Fresh[7124], Fresh[7123], Fresh[7122], Fresh[7121], Fresh[7120], Fresh[7119], Fresh[7118], Fresh[7117], Fresh[7116], Fresh[7115], Fresh[7114], Fresh[7113], Fresh[7112], Fresh[7111], Fresh[7110], Fresh[7109], Fresh[7108], Fresh[7107], Fresh[7106], Fresh[7105], Fresh[7104], Fresh[7103], Fresh[7102], Fresh[7101], Fresh[7100], Fresh[7099], Fresh[7098], Fresh[7097], Fresh[7096], Fresh[7095], Fresh[7094], Fresh[7093], Fresh[7092], Fresh[7091], Fresh[7090], Fresh[7089], Fresh[7088], Fresh[7087], Fresh[7086], Fresh[7085], Fresh[7084], Fresh[7083], Fresh[7082], Fresh[7081], Fresh[7080], Fresh[7079], Fresh[7078], Fresh[7077], Fresh[7076], Fresh[7075], Fresh[7074], Fresh[7073], Fresh[7072], Fresh[7071], Fresh[7070], Fresh[7069], Fresh[7068], Fresh[7067], Fresh[7066], Fresh[7065], Fresh[7064], Fresh[7063], Fresh[7062], Fresh[7061], Fresh[7060], Fresh[7059], Fresh[7058], Fresh[7057], Fresh[7056], Fresh[7055], Fresh[7054], Fresh[7053], Fresh[7052], Fresh[7051], Fresh[7050], Fresh[7049], Fresh[7048], Fresh[7047], Fresh[7046], Fresh[7045], Fresh[7044], Fresh[7043], Fresh[7042], Fresh[7041], Fresh[7040], Fresh[7039], Fresh[7038], Fresh[7037], Fresh[7036], Fresh[7035], Fresh[7034], Fresh[7033], Fresh[7032], Fresh[7031], Fresh[7030], Fresh[7029], Fresh[7028], Fresh[7027], Fresh[7026], Fresh[7025], Fresh[7024], Fresh[7023], Fresh[7022], Fresh[7021], Fresh[7020], Fresh[7019], Fresh[7018], Fresh[7017], Fresh[7016], Fresh[7015], Fresh[7014], Fresh[7013], Fresh[7012], Fresh[7011], Fresh[7010], Fresh[7009], Fresh[7008], Fresh[7007], Fresh[7006], Fresh[7005], Fresh[7004], Fresh[7003], Fresh[7002], Fresh[7001], Fresh[7000], Fresh[6999], Fresh[6998], Fresh[6997], Fresh[6996], Fresh[6995], Fresh[6994], Fresh[6993], Fresh[6992], Fresh[6991], Fresh[6990], Fresh[6989], Fresh[6988], Fresh[6987], Fresh[6986], Fresh[6985], Fresh[6984], Fresh[6983], Fresh[6982], Fresh[6981], Fresh[6980], Fresh[6979], Fresh[6978], Fresh[6977], Fresh[6976], Fresh[6975], Fresh[6974], Fresh[6973], Fresh[6972], Fresh[6971], Fresh[6970], Fresh[6969], Fresh[6968], Fresh[6967], Fresh[6966], Fresh[6965], Fresh[6964], Fresh[6963], Fresh[6962], Fresh[6961], Fresh[6960], Fresh[6959], Fresh[6958], Fresh[6957], Fresh[6956], Fresh[6955], Fresh[6954], Fresh[6953], Fresh[6952], Fresh[6951], Fresh[6950], Fresh[6949], Fresh[6948], Fresh[6947], Fresh[6946], Fresh[6945], Fresh[6944], Fresh[6943], Fresh[6942], Fresh[6941], Fresh[6940], Fresh[6939], Fresh[6938], Fresh[6937], Fresh[6936], Fresh[6935], Fresh[6934], Fresh[6933], Fresh[6932], Fresh[6931], Fresh[6930], Fresh[6929], Fresh[6928], Fresh[6927], Fresh[6926], Fresh[6925], Fresh[6924], Fresh[6923], Fresh[6922], Fresh[6921], Fresh[6920], Fresh[6919], Fresh[6918], Fresh[6917], Fresh[6916], Fresh[6915], Fresh[6914], Fresh[6913], Fresh[6912], Fresh[6911], Fresh[6910], Fresh[6909], Fresh[6908], Fresh[6907], Fresh[6906], Fresh[6905], Fresh[6904], Fresh[6903], Fresh[6902], Fresh[6901], Fresh[6900], Fresh[6899], Fresh[6898], Fresh[6897], Fresh[6896], Fresh[6895], Fresh[6894], Fresh[6893], Fresh[6892], Fresh[6891], Fresh[6890], Fresh[6889], Fresh[6888], Fresh[6887], Fresh[6886], Fresh[6885], Fresh[6884], Fresh[6883], Fresh[6882], Fresh[6881], Fresh[6880], Fresh[6879], Fresh[6878], Fresh[6877], Fresh[6876], Fresh[6875], Fresh[6874], Fresh[6873], Fresh[6872], Fresh[6871], Fresh[6870], Fresh[6869], Fresh[6868], Fresh[6867], Fresh[6866], Fresh[6865], Fresh[6864], Fresh[6863], Fresh[6862], Fresh[6861], Fresh[6860], Fresh[6859], Fresh[6858], Fresh[6857], Fresh[6856], Fresh[6855], Fresh[6854], Fresh[6853], Fresh[6852], Fresh[6851], Fresh[6850], Fresh[6849], Fresh[6848], Fresh[6847], Fresh[6846], Fresh[6845], Fresh[6844], Fresh[6843], Fresh[6842], Fresh[6841], Fresh[6840], Fresh[6839], Fresh[6838], Fresh[6837], Fresh[6836], Fresh[6835], Fresh[6834], Fresh[6833], Fresh[6832], Fresh[6831], Fresh[6830], Fresh[6829], Fresh[6828], Fresh[6827], Fresh[6826], Fresh[6825], Fresh[6824], Fresh[6823], Fresh[6822], Fresh[6821], Fresh[6820], Fresh[6819], Fresh[6818], Fresh[6817], Fresh[6816], Fresh[6815], Fresh[6814], Fresh[6813], Fresh[6812], Fresh[6811], Fresh[6810], Fresh[6809], Fresh[6808], Fresh[6807], Fresh[6806], Fresh[6805], Fresh[6804], Fresh[6803], Fresh[6802], Fresh[6801], Fresh[6800], Fresh[6799], Fresh[6798], Fresh[6797], Fresh[6796], Fresh[6795], Fresh[6794], Fresh[6793], Fresh[6792], Fresh[6791], Fresh[6790], Fresh[6789], Fresh[6788], Fresh[6787], Fresh[6786], Fresh[6785], Fresh[6784], Fresh[6783], Fresh[6782], Fresh[6781], Fresh[6780], Fresh[6779], Fresh[6778], Fresh[6777], Fresh[6776], Fresh[6775], Fresh[6774], Fresh[6773], Fresh[6772], Fresh[6771], Fresh[6770], Fresh[6769], Fresh[6768], Fresh[6767], Fresh[6766], Fresh[6765], Fresh[6764], Fresh[6763], Fresh[6762], Fresh[6761], Fresh[6760], Fresh[6759], Fresh[6758], Fresh[6757], Fresh[6756], Fresh[6755], Fresh[6754], Fresh[6753], Fresh[6752], Fresh[6751], Fresh[6750], Fresh[6749], Fresh[6748], Fresh[6747], Fresh[6746], Fresh[6745], Fresh[6744], Fresh[6743], Fresh[6742], Fresh[6741], Fresh[6740], Fresh[6739], Fresh[6738], Fresh[6737], Fresh[6736], Fresh[6735], Fresh[6734], Fresh[6733], Fresh[6732], Fresh[6731], Fresh[6730], Fresh[6729], Fresh[6728], Fresh[6727], Fresh[6726], Fresh[6725], Fresh[6724], Fresh[6723], Fresh[6722], Fresh[6721], Fresh[6720], Fresh[6719], Fresh[6718], Fresh[6717], Fresh[6716], Fresh[6715], Fresh[6714], Fresh[6713], Fresh[6712], Fresh[6711], Fresh[6710], Fresh[6709], Fresh[6708], Fresh[6707], Fresh[6706], Fresh[6705], Fresh[6704], Fresh[6703], Fresh[6702], Fresh[6701], Fresh[6700], Fresh[6699], Fresh[6698], Fresh[6697], Fresh[6696], Fresh[6695], Fresh[6694], Fresh[6693], Fresh[6692], Fresh[6691], Fresh[6690], Fresh[6689], Fresh[6688], Fresh[6687], Fresh[6686], Fresh[6685], Fresh[6684], Fresh[6683], Fresh[6682], Fresh[6681], Fresh[6680], Fresh[6679], Fresh[6678], Fresh[6677], Fresh[6676], Fresh[6675], Fresh[6674], Fresh[6673], Fresh[6672], Fresh[6671], Fresh[6670], Fresh[6669], Fresh[6668], Fresh[6667], Fresh[6666], Fresh[6665], Fresh[6664], Fresh[6663], Fresh[6662], Fresh[6661], Fresh[6660], Fresh[6659], Fresh[6658], Fresh[6657], Fresh[6656], Fresh[6655], Fresh[6654], Fresh[6653], Fresh[6652], Fresh[6651], Fresh[6650], Fresh[6649], Fresh[6648], Fresh[6647], Fresh[6646], Fresh[6645], Fresh[6644], Fresh[6643], Fresh[6642], Fresh[6641], Fresh[6640], Fresh[6639], Fresh[6638], Fresh[6637], Fresh[6636], Fresh[6635], Fresh[6634], Fresh[6633], Fresh[6632], Fresh[6631], Fresh[6630], Fresh[6629], Fresh[6628], Fresh[6627], Fresh[6626], Fresh[6625], Fresh[6624], Fresh[6623], Fresh[6622], Fresh[6621], Fresh[6620], Fresh[6619], Fresh[6618], Fresh[6617], Fresh[6616], Fresh[6615], Fresh[6614], Fresh[6613], Fresh[6612], Fresh[6611], Fresh[6610], Fresh[6609], Fresh[6608], Fresh[6607], Fresh[6606], Fresh[6605], Fresh[6604], Fresh[6603], Fresh[6602], Fresh[6601], Fresh[6600], Fresh[6599], Fresh[6598], Fresh[6597], Fresh[6596], Fresh[6595], Fresh[6594], Fresh[6593], Fresh[6592], Fresh[6591], Fresh[6590], Fresh[6589], Fresh[6588], Fresh[6587], Fresh[6586], Fresh[6585], Fresh[6584], Fresh[6583], Fresh[6582], Fresh[6581], Fresh[6580], Fresh[6579], Fresh[6578], Fresh[6577], Fresh[6576], Fresh[6575], Fresh[6574], Fresh[6573], Fresh[6572], Fresh[6571], Fresh[6570], Fresh[6569], Fresh[6568], Fresh[6567], Fresh[6566], Fresh[6565], Fresh[6564], Fresh[6563], Fresh[6562], Fresh[6561], Fresh[6560], Fresh[6559], Fresh[6558], Fresh[6557], Fresh[6556], Fresh[6555], Fresh[6554], Fresh[6553], Fresh[6552], Fresh[6551], Fresh[6550], Fresh[6549], Fresh[6548], Fresh[6547], Fresh[6546], Fresh[6545], Fresh[6544], Fresh[6543], Fresh[6542], Fresh[6541], Fresh[6540], Fresh[6539], Fresh[6538], Fresh[6537], Fresh[6536], Fresh[6535], Fresh[6534], Fresh[6533], Fresh[6532], Fresh[6531], Fresh[6530], Fresh[6529], Fresh[6528], Fresh[6527], Fresh[6526], Fresh[6525], Fresh[6524], Fresh[6523], Fresh[6522], Fresh[6521], Fresh[6520], Fresh[6519], Fresh[6518], Fresh[6517], Fresh[6516], Fresh[6515], Fresh[6514], Fresh[6513], Fresh[6512], Fresh[6511], Fresh[6510], Fresh[6509], Fresh[6508], Fresh[6507], Fresh[6506], Fresh[6505], Fresh[6504], Fresh[6503], Fresh[6502], Fresh[6501], Fresh[6500], Fresh[6499], Fresh[6498], Fresh[6497], Fresh[6496], Fresh[6495], Fresh[6494], Fresh[6493], Fresh[6492], Fresh[6491], Fresh[6490], Fresh[6489], Fresh[6488], Fresh[6487], Fresh[6486], Fresh[6485], Fresh[6484], Fresh[6483], Fresh[6482], Fresh[6481], Fresh[6480], Fresh[6479], Fresh[6478], Fresh[6477], Fresh[6476], Fresh[6475], Fresh[6474], Fresh[6473], Fresh[6472], Fresh[6471], Fresh[6470], Fresh[6469], Fresh[6468], Fresh[6467], Fresh[6466], Fresh[6465], Fresh[6464], Fresh[6463], Fresh[6462], Fresh[6461], Fresh[6460], Fresh[6459], Fresh[6458], Fresh[6457], Fresh[6456], Fresh[6455], Fresh[6454], Fresh[6453], Fresh[6452], Fresh[6451], Fresh[6450], Fresh[6449], Fresh[6448], Fresh[6447], Fresh[6446], Fresh[6445], Fresh[6444], Fresh[6443], Fresh[6442], Fresh[6441], Fresh[6440], Fresh[6439], Fresh[6438], Fresh[6437], Fresh[6436], Fresh[6435], Fresh[6434], Fresh[6433], Fresh[6432], Fresh[6431], Fresh[6430], Fresh[6429], Fresh[6428], Fresh[6427], Fresh[6426], Fresh[6425], Fresh[6424], Fresh[6423], Fresh[6422], Fresh[6421], Fresh[6420], Fresh[6419], Fresh[6418], Fresh[6417], Fresh[6416], Fresh[6415], Fresh[6414], Fresh[6413], Fresh[6412], Fresh[6411], Fresh[6410], Fresh[6409], Fresh[6408], Fresh[6407], Fresh[6406], Fresh[6405], Fresh[6404], Fresh[6403], Fresh[6402], Fresh[6401], Fresh[6400], Fresh[6399], Fresh[6398], Fresh[6397], Fresh[6396], Fresh[6395], Fresh[6394], Fresh[6393], Fresh[6392], Fresh[6391], Fresh[6390], Fresh[6389], Fresh[6388], Fresh[6387], Fresh[6386], Fresh[6385], Fresh[6384], Fresh[6383], Fresh[6382], Fresh[6381], Fresh[6380], Fresh[6379], Fresh[6378], Fresh[6377], Fresh[6376], Fresh[6375], Fresh[6374], Fresh[6373], Fresh[6372], Fresh[6371], Fresh[6370], Fresh[6369], Fresh[6368], Fresh[6367], Fresh[6366], Fresh[6365], Fresh[6364], Fresh[6363], Fresh[6362], Fresh[6361], Fresh[6360], Fresh[6359], Fresh[6358], Fresh[6357], Fresh[6356], Fresh[6355], Fresh[6354], Fresh[6353], Fresh[6352], Fresh[6351], Fresh[6350], Fresh[6349], Fresh[6348], Fresh[6347], Fresh[6346], Fresh[6345], Fresh[6344], Fresh[6343], Fresh[6342], Fresh[6341], Fresh[6340], Fresh[6339], Fresh[6338], Fresh[6337], Fresh[6336], Fresh[6335], Fresh[6334], Fresh[6333], Fresh[6332], Fresh[6331], Fresh[6330], Fresh[6329], Fresh[6328], Fresh[6327], Fresh[6326], Fresh[6325], Fresh[6324], Fresh[6323], Fresh[6322], Fresh[6321], Fresh[6320], Fresh[6319], Fresh[6318], Fresh[6317], Fresh[6316], Fresh[6315], Fresh[6314], Fresh[6313], Fresh[6312], Fresh[6311], Fresh[6310], Fresh[6309], Fresh[6308], Fresh[6307], Fresh[6306], Fresh[6305], Fresh[6304], Fresh[6303], Fresh[6302], Fresh[6301], Fresh[6300], Fresh[6299], Fresh[6298], Fresh[6297], Fresh[6296], Fresh[6295], Fresh[6294], Fresh[6293], Fresh[6292], Fresh[6291], Fresh[6290], Fresh[6289], Fresh[6288], Fresh[6287], Fresh[6286], Fresh[6285], Fresh[6284], Fresh[6283], Fresh[6282], Fresh[6281], Fresh[6280], Fresh[6279], Fresh[6278], Fresh[6277], Fresh[6276], Fresh[6275], Fresh[6274], Fresh[6273], Fresh[6272], Fresh[6271], Fresh[6270], Fresh[6269], Fresh[6268], Fresh[6267], Fresh[6266], Fresh[6265], Fresh[6264], Fresh[6263], Fresh[6262], Fresh[6261], Fresh[6260], Fresh[6259], Fresh[6258], Fresh[6257], Fresh[6256], Fresh[6255], Fresh[6254], Fresh[6253], Fresh[6252], Fresh[6251], Fresh[6250], Fresh[6249], Fresh[6248], Fresh[6247], Fresh[6246], Fresh[6245], Fresh[6244], Fresh[6243], Fresh[6242], Fresh[6241], Fresh[6240], Fresh[6239], Fresh[6238], Fresh[6237], Fresh[6236], Fresh[6235], Fresh[6234], Fresh[6233], Fresh[6232], Fresh[6231], Fresh[6230], Fresh[6229], Fresh[6228], Fresh[6227], Fresh[6226], Fresh[6225], Fresh[6224], Fresh[6223], Fresh[6222], Fresh[6221], Fresh[6220], Fresh[6219], Fresh[6218], Fresh[6217], Fresh[6216], Fresh[6215], Fresh[6214], Fresh[6213], Fresh[6212], Fresh[6211], Fresh[6210], Fresh[6209], Fresh[6208], Fresh[6207], Fresh[6206], Fresh[6205], Fresh[6204], Fresh[6203], Fresh[6202], Fresh[6201], Fresh[6200], Fresh[6199], Fresh[6198], Fresh[6197], Fresh[6196], Fresh[6195], Fresh[6194], Fresh[6193], Fresh[6192], Fresh[6191], Fresh[6190], Fresh[6189], Fresh[6188], Fresh[6187], Fresh[6186], Fresh[6185], Fresh[6184], Fresh[6183], Fresh[6182], Fresh[6181], Fresh[6180], Fresh[6179], Fresh[6178], Fresh[6177], Fresh[6176], Fresh[6175], Fresh[6174], Fresh[6173], Fresh[6172], Fresh[6171], Fresh[6170], Fresh[6169], Fresh[6168], Fresh[6167], Fresh[6166], Fresh[6165], Fresh[6164], Fresh[6163], Fresh[6162], Fresh[6161], Fresh[6160], Fresh[6159], Fresh[6158], Fresh[6157], Fresh[6156], Fresh[6155], Fresh[6154], Fresh[6153], Fresh[6152], Fresh[6151], Fresh[6150], Fresh[6149], Fresh[6148], Fresh[6147], Fresh[6146], Fresh[6145], Fresh[6144], Fresh[6143], Fresh[6142], Fresh[6141], Fresh[6140], Fresh[6139], Fresh[6138], Fresh[6137], Fresh[6136], Fresh[6135], Fresh[6134], Fresh[6133], Fresh[6132], Fresh[6131], Fresh[6130], Fresh[6129], Fresh[6128], Fresh[6127], Fresh[6126], Fresh[6125], Fresh[6124], Fresh[6123], Fresh[6122], Fresh[6121], Fresh[6120], Fresh[6119], Fresh[6118], Fresh[6117], Fresh[6116], Fresh[6115], Fresh[6114], Fresh[6113], Fresh[6112], Fresh[6111], Fresh[6110], Fresh[6109], Fresh[6108], Fresh[6107], Fresh[6106], Fresh[6105], Fresh[6104], Fresh[6103], Fresh[6102], Fresh[6101], Fresh[6100], Fresh[6099], Fresh[6098], Fresh[6097], Fresh[6096], Fresh[6095], Fresh[6094], Fresh[6093], Fresh[6092], Fresh[6091], Fresh[6090], Fresh[6089], Fresh[6088], Fresh[6087], Fresh[6086], Fresh[6085], Fresh[6084], Fresh[6083], Fresh[6082], Fresh[6081], Fresh[6080], Fresh[6079], Fresh[6078], Fresh[6077], Fresh[6076], Fresh[6075], Fresh[6074], Fresh[6073], Fresh[6072], Fresh[6071], Fresh[6070], Fresh[6069], Fresh[6068], Fresh[6067], Fresh[6066], Fresh[6065], Fresh[6064], Fresh[6063], Fresh[6062], Fresh[6061], Fresh[6060], Fresh[6059], Fresh[6058], Fresh[6057], Fresh[6056], Fresh[6055], Fresh[6054], Fresh[6053], Fresh[6052], Fresh[6051], Fresh[6050], Fresh[6049], Fresh[6048], Fresh[6047], Fresh[6046], Fresh[6045], Fresh[6044], Fresh[6043], Fresh[6042], Fresh[6041], Fresh[6040], Fresh[6039], Fresh[6038], Fresh[6037], Fresh[6036], Fresh[6035], Fresh[6034], Fresh[6033], Fresh[6032], Fresh[6031], Fresh[6030], Fresh[6029], Fresh[6028], Fresh[6027], Fresh[6026], Fresh[6025], Fresh[6024], Fresh[6023], Fresh[6022], Fresh[6021], Fresh[6020], Fresh[6019], Fresh[6018], Fresh[6017], Fresh[6016], Fresh[6015], Fresh[6014], Fresh[6013], Fresh[6012], Fresh[6011], Fresh[6010], Fresh[6009], Fresh[6008], Fresh[6007], Fresh[6006], Fresh[6005], Fresh[6004], Fresh[6003], Fresh[6002], Fresh[6001], Fresh[6000], Fresh[5999], Fresh[5998], Fresh[5997], Fresh[5996], Fresh[5995], Fresh[5994], Fresh[5993], Fresh[5992], Fresh[5991], Fresh[5990], Fresh[5989], Fresh[5988], Fresh[5987], Fresh[5986], Fresh[5985], Fresh[5984], Fresh[5983], Fresh[5982], Fresh[5981], Fresh[5980], Fresh[5979], Fresh[5978], Fresh[5977], Fresh[5976], Fresh[5975], Fresh[5974], Fresh[5973], Fresh[5972], Fresh[5971], Fresh[5970], Fresh[5969], Fresh[5968], Fresh[5967], Fresh[5966], Fresh[5965], Fresh[5964], Fresh[5963], Fresh[5962], Fresh[5961], Fresh[5960], Fresh[5959], Fresh[5958], Fresh[5957], Fresh[5956], Fresh[5955], Fresh[5954], Fresh[5953], Fresh[5952], Fresh[5951], Fresh[5950], Fresh[5949], Fresh[5948], Fresh[5947], Fresh[5946], Fresh[5945], Fresh[5944], Fresh[5943], Fresh[5942], Fresh[5941], Fresh[5940], Fresh[5939], Fresh[5938], Fresh[5937], Fresh[5936], Fresh[5935], Fresh[5934], Fresh[5933], Fresh[5932], Fresh[5931], Fresh[5930], Fresh[5929], Fresh[5928], Fresh[5927], Fresh[5926], Fresh[5925], Fresh[5924], Fresh[5923], Fresh[5922], Fresh[5921], Fresh[5920], Fresh[5919], Fresh[5918], Fresh[5917], Fresh[5916], Fresh[5915], Fresh[5914], Fresh[5913], Fresh[5912], Fresh[5911], Fresh[5910], Fresh[5909], Fresh[5908], Fresh[5907], Fresh[5906], Fresh[5905], Fresh[5904], Fresh[5903], Fresh[5902], Fresh[5901], Fresh[5900], Fresh[5899], Fresh[5898], Fresh[5897], Fresh[5896], Fresh[5895], Fresh[5894], Fresh[5893], Fresh[5892], Fresh[5891], Fresh[5890], Fresh[5889], Fresh[5888], Fresh[5887], Fresh[5886], Fresh[5885], Fresh[5884], Fresh[5883], Fresh[5882], Fresh[5881], Fresh[5880], Fresh[5879], Fresh[5878], Fresh[5877], Fresh[5876], Fresh[5875], Fresh[5874], Fresh[5873], Fresh[5872], Fresh[5871], Fresh[5870], Fresh[5869], Fresh[5868], Fresh[5867], Fresh[5866], Fresh[5865], Fresh[5864], Fresh[5863], Fresh[5862], Fresh[5861], Fresh[5860], Fresh[5859], Fresh[5858], Fresh[5857], Fresh[5856], Fresh[5855], Fresh[5854], Fresh[5853], Fresh[5852], Fresh[5851], Fresh[5850], Fresh[5849], Fresh[5848], Fresh[5847], Fresh[5846], Fresh[5845], Fresh[5844], Fresh[5843], Fresh[5842], Fresh[5841], Fresh[5840], Fresh[5839], Fresh[5838], Fresh[5837], Fresh[5836], Fresh[5835], Fresh[5834], Fresh[5833], Fresh[5832], Fresh[5831], Fresh[5830], Fresh[5829], Fresh[5828], Fresh[5827], Fresh[5826], Fresh[5825], Fresh[5824], Fresh[5823], Fresh[5822], Fresh[5821], Fresh[5820], Fresh[5819], Fresh[5818], Fresh[5817], Fresh[5816], Fresh[5815], Fresh[5814], Fresh[5813], Fresh[5812], Fresh[5811], Fresh[5810], Fresh[5809], Fresh[5808], Fresh[5807], Fresh[5806], Fresh[5805], Fresh[5804], Fresh[5803], Fresh[5802], Fresh[5801], Fresh[5800], Fresh[5799], Fresh[5798], Fresh[5797], Fresh[5796], Fresh[5795], Fresh[5794], Fresh[5793], Fresh[5792], Fresh[5791], Fresh[5790], Fresh[5789], Fresh[5788], Fresh[5787], Fresh[5786], Fresh[5785], Fresh[5784], Fresh[5783], Fresh[5782], Fresh[5781], Fresh[5780], Fresh[5779], Fresh[5778], Fresh[5777], Fresh[5776], Fresh[5775], Fresh[5774], Fresh[5773], Fresh[5772], Fresh[5771], Fresh[5770], Fresh[5769], Fresh[5768], Fresh[5767], Fresh[5766], Fresh[5765], Fresh[5764], Fresh[5763], Fresh[5762], Fresh[5761], Fresh[5760], Fresh[5759], Fresh[5758], Fresh[5757], Fresh[5756], Fresh[5755], Fresh[5754], Fresh[5753], Fresh[5752], Fresh[5751], Fresh[5750], Fresh[5749], Fresh[5748], Fresh[5747], Fresh[5746], Fresh[5745], Fresh[5744], Fresh[5743], Fresh[5742], Fresh[5741], Fresh[5740], Fresh[5739], Fresh[5738], Fresh[5737], Fresh[5736], Fresh[5735], Fresh[5734], Fresh[5733], Fresh[5732], Fresh[5731], Fresh[5730], Fresh[5729], Fresh[5728], Fresh[5727], Fresh[5726], Fresh[5725], Fresh[5724], Fresh[5723], Fresh[5722], Fresh[5721], Fresh[5720], Fresh[5719], Fresh[5718], Fresh[5717], Fresh[5716], Fresh[5715], Fresh[5714], Fresh[5713], Fresh[5712], Fresh[5711], Fresh[5710], Fresh[5709], Fresh[5708], Fresh[5707], Fresh[5706], Fresh[5705], Fresh[5704], Fresh[5703], Fresh[5702], Fresh[5701], Fresh[5700], Fresh[5699], Fresh[5698], Fresh[5697], Fresh[5696], Fresh[5695], Fresh[5694], Fresh[5693], Fresh[5692], Fresh[5691], Fresh[5690], Fresh[5689], Fresh[5688], Fresh[5687], Fresh[5686], Fresh[5685], Fresh[5684], Fresh[5683], Fresh[5682], Fresh[5681], Fresh[5680], Fresh[5679], Fresh[5678], Fresh[5677], Fresh[5676], Fresh[5675], Fresh[5674], Fresh[5673], Fresh[5672], Fresh[5671], Fresh[5670], Fresh[5669], Fresh[5668], Fresh[5667], Fresh[5666], Fresh[5665], Fresh[5664], Fresh[5663], Fresh[5662], Fresh[5661], Fresh[5660], Fresh[5659], Fresh[5658], Fresh[5657], Fresh[5656], Fresh[5655], Fresh[5654], Fresh[5653], Fresh[5652], Fresh[5651], Fresh[5650], Fresh[5649], Fresh[5648], Fresh[5647], Fresh[5646], Fresh[5645], Fresh[5644], Fresh[5643], Fresh[5642], Fresh[5641], Fresh[5640], Fresh[5639], Fresh[5638], Fresh[5637], Fresh[5636], Fresh[5635], Fresh[5634], Fresh[5633], Fresh[5632], Fresh[5631], Fresh[5630], Fresh[5629], Fresh[5628], Fresh[5627], Fresh[5626], Fresh[5625], Fresh[5624], Fresh[5623], Fresh[5622], Fresh[5621], Fresh[5620], Fresh[5619], Fresh[5618], Fresh[5617], Fresh[5616], Fresh[5615], Fresh[5614], Fresh[5613], Fresh[5612], Fresh[5611], Fresh[5610], Fresh[5609], Fresh[5608], Fresh[5607], Fresh[5606], Fresh[5605], Fresh[5604], Fresh[5603], Fresh[5602], Fresh[5601], Fresh[5600], Fresh[5599], Fresh[5598], Fresh[5597], Fresh[5596], Fresh[5595], Fresh[5594], Fresh[5593], Fresh[5592], Fresh[5591], Fresh[5590], Fresh[5589], Fresh[5588], Fresh[5587], Fresh[5586], Fresh[5585], Fresh[5584], Fresh[5583], Fresh[5582], Fresh[5581], Fresh[5580], Fresh[5579], Fresh[5578], Fresh[5577], Fresh[5576], Fresh[5575], Fresh[5574], Fresh[5573], Fresh[5572], Fresh[5571], Fresh[5570], Fresh[5569], Fresh[5568], Fresh[5567], Fresh[5566], Fresh[5565], Fresh[5564], Fresh[5563], Fresh[5562], Fresh[5561], Fresh[5560], Fresh[5559], Fresh[5558], Fresh[5557], Fresh[5556], Fresh[5555], Fresh[5554], Fresh[5553], Fresh[5552], Fresh[5551], Fresh[5550], Fresh[5549], Fresh[5548], Fresh[5547], Fresh[5546], Fresh[5545], Fresh[5544], Fresh[5543], Fresh[5542], Fresh[5541], Fresh[5540], Fresh[5539], Fresh[5538], Fresh[5537], Fresh[5536], Fresh[5535], Fresh[5534], Fresh[5533], Fresh[5532], Fresh[5531], Fresh[5530], Fresh[5529], Fresh[5528], Fresh[5527], Fresh[5526], Fresh[5525], Fresh[5524], Fresh[5523], Fresh[5522], Fresh[5521], Fresh[5520], Fresh[5519], Fresh[5518], Fresh[5517], Fresh[5516], Fresh[5515], Fresh[5514], Fresh[5513], Fresh[5512], Fresh[5511], Fresh[5510], Fresh[5509], Fresh[5508], Fresh[5507], Fresh[5506], Fresh[5505], Fresh[5504], Fresh[5503], Fresh[5502], Fresh[5501], Fresh[5500], Fresh[5499], Fresh[5498], Fresh[5497], Fresh[5496], Fresh[5495], Fresh[5494], Fresh[5493], Fresh[5492], Fresh[5491], Fresh[5490], Fresh[5489], Fresh[5488], Fresh[5487], Fresh[5486], Fresh[5485], Fresh[5484], Fresh[5483], Fresh[5482], Fresh[5481], Fresh[5480], Fresh[5479], Fresh[5478], Fresh[5477], Fresh[5476], Fresh[5475], Fresh[5474], Fresh[5473], Fresh[5472], Fresh[5471], Fresh[5470], Fresh[5469], Fresh[5468], Fresh[5467], Fresh[5466], Fresh[5465], Fresh[5464], Fresh[5463], Fresh[5462], Fresh[5461], Fresh[5460], Fresh[5459], Fresh[5458], Fresh[5457], Fresh[5456], Fresh[5455], Fresh[5454], Fresh[5453], Fresh[5452], Fresh[5451], Fresh[5450], Fresh[5449], Fresh[5448], Fresh[5447], Fresh[5446], Fresh[5445], Fresh[5444], Fresh[5443], Fresh[5442], Fresh[5441], Fresh[5440], Fresh[5439], Fresh[5438], Fresh[5437], Fresh[5436], Fresh[5435], Fresh[5434], Fresh[5433], Fresh[5432], Fresh[5431], Fresh[5430], Fresh[5429], Fresh[5428], Fresh[5427], Fresh[5426], Fresh[5425], Fresh[5424], Fresh[5423], Fresh[5422], Fresh[5421], Fresh[5420], Fresh[5419], Fresh[5418], Fresh[5417], Fresh[5416], Fresh[5415], Fresh[5414], Fresh[5413], Fresh[5412], Fresh[5411], Fresh[5410], Fresh[5409], Fresh[5408], Fresh[5407], Fresh[5406], Fresh[5405], Fresh[5404], Fresh[5403], Fresh[5402], Fresh[5401], Fresh[5400], Fresh[5399], Fresh[5398], Fresh[5397], Fresh[5396], Fresh[5395], Fresh[5394], Fresh[5393], Fresh[5392], Fresh[5391], Fresh[5390], Fresh[5389], Fresh[5388], Fresh[5387], Fresh[5386], Fresh[5385], Fresh[5384], Fresh[5383], Fresh[5382], Fresh[5381], Fresh[5380], Fresh[5379], Fresh[5378], Fresh[5377], Fresh[5376], Fresh[5375], Fresh[5374], Fresh[5373], Fresh[5372], Fresh[5371], Fresh[5370], Fresh[5369], Fresh[5368], Fresh[5367], Fresh[5366], Fresh[5365], Fresh[5364], Fresh[5363], Fresh[5362], Fresh[5361], Fresh[5360], Fresh[5359], Fresh[5358], Fresh[5357], Fresh[5356], Fresh[5355], Fresh[5354], Fresh[5353], Fresh[5352], Fresh[5351], Fresh[5350], Fresh[5349], Fresh[5348], Fresh[5347], Fresh[5346], Fresh[5345], Fresh[5344], Fresh[5343], Fresh[5342], Fresh[5341], Fresh[5340], Fresh[5339], Fresh[5338], Fresh[5337], Fresh[5336], Fresh[5335], Fresh[5334], Fresh[5333], Fresh[5332], Fresh[5331], Fresh[5330], Fresh[5329], Fresh[5328], Fresh[5327], Fresh[5326], Fresh[5325], Fresh[5324], Fresh[5323], Fresh[5322], Fresh[5321], Fresh[5320], Fresh[5319], Fresh[5318], Fresh[5317], Fresh[5316], Fresh[5315], Fresh[5314], Fresh[5313], Fresh[5312], Fresh[5311], Fresh[5310], Fresh[5309], Fresh[5308], Fresh[5307], Fresh[5306], Fresh[5305], Fresh[5304], Fresh[5303], Fresh[5302], Fresh[5301], Fresh[5300], Fresh[5299], Fresh[5298], Fresh[5297], Fresh[5296], Fresh[5295], Fresh[5294], Fresh[5293], Fresh[5292], Fresh[5291], Fresh[5290], Fresh[5289], Fresh[5288], Fresh[5287], Fresh[5286], Fresh[5285], Fresh[5284], Fresh[5283], Fresh[5282], Fresh[5281], Fresh[5280], Fresh[5279], Fresh[5278], Fresh[5277], Fresh[5276], Fresh[5275], Fresh[5274], Fresh[5273], Fresh[5272], Fresh[5271], Fresh[5270], Fresh[5269], Fresh[5268], Fresh[5267], Fresh[5266], Fresh[5265], Fresh[5264], Fresh[5263], Fresh[5262], Fresh[5261], Fresh[5260], Fresh[5259], Fresh[5258], Fresh[5257], Fresh[5256], Fresh[5255], Fresh[5254], Fresh[5253], Fresh[5252], Fresh[5251], Fresh[5250], Fresh[5249], Fresh[5248], Fresh[5247], Fresh[5246], Fresh[5245], Fresh[5244], Fresh[5243], Fresh[5242], Fresh[5241], Fresh[5240], Fresh[5239], Fresh[5238], Fresh[5237], Fresh[5236], Fresh[5235], Fresh[5234], Fresh[5233], Fresh[5232], Fresh[5231], Fresh[5230], Fresh[5229], Fresh[5228], Fresh[5227], Fresh[5226], Fresh[5225], Fresh[5224], Fresh[5223], Fresh[5222], Fresh[5221], Fresh[5220], Fresh[5219], Fresh[5218], Fresh[5217], Fresh[5216], Fresh[5215], Fresh[5214], Fresh[5213], Fresh[5212], Fresh[5211], Fresh[5210], Fresh[5209], Fresh[5208], Fresh[5207], Fresh[5206], Fresh[5205], Fresh[5204], Fresh[5203], Fresh[5202], Fresh[5201], Fresh[5200], Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196], Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190], Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184], Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180], Fresh[5179], Fresh[5178], Fresh[5177], Fresh[5176], Fresh[5175], Fresh[5174], Fresh[5173], Fresh[5172], Fresh[5171], Fresh[5170], Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166], Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160], Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154], Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150], Fresh[5149], Fresh[5148], Fresh[5147], Fresh[5146], Fresh[5145], Fresh[5144], Fresh[5143], Fresh[5142], Fresh[5141], Fresh[5140], Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136], Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130], Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124], Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120], Fresh[5119], Fresh[5118], Fresh[5117], Fresh[5116], Fresh[5115], Fresh[5114], Fresh[5113], Fresh[5112], Fresh[5111], Fresh[5110], Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106], Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100], Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094], Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090], Fresh[5089], Fresh[5088], Fresh[5087], Fresh[5086], Fresh[5085], Fresh[5084], Fresh[5083], Fresh[5082], Fresh[5081], Fresh[5080], Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076], Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070], Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064], Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060], Fresh[5059], Fresh[5058], Fresh[5057], Fresh[5056], Fresh[5055], Fresh[5054], Fresh[5053], Fresh[5052], Fresh[5051], Fresh[5050], Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046], Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040], Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034], Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030], Fresh[5029], Fresh[5028], Fresh[5027], Fresh[5026], Fresh[5025], Fresh[5024], Fresh[5023], Fresh[5022], Fresh[5021], Fresh[5020], Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016], Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010], Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004], Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000], Fresh[4999], Fresh[4998], Fresh[4997], Fresh[4996], Fresh[4995], Fresh[4994], Fresh[4993], Fresh[4992], Fresh[4991], Fresh[4990], Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986], Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980], Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974], Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970], Fresh[4969], Fresh[4968], Fresh[4967], Fresh[4966], Fresh[4965], Fresh[4964], Fresh[4963], Fresh[4962], Fresh[4961], Fresh[4960], Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956], Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950], Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944], Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940], Fresh[4939], Fresh[4938], Fresh[4937], Fresh[4936], Fresh[4935], Fresh[4934], Fresh[4933], Fresh[4932], Fresh[4931], Fresh[4930], Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926], Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920], Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914], Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910], Fresh[4909], Fresh[4908], Fresh[4907], Fresh[4906], Fresh[4905], Fresh[4904], Fresh[4903], Fresh[4902], Fresh[4901], Fresh[4900], Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896], Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890], Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884], Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880], Fresh[4879], Fresh[4878], Fresh[4877], Fresh[4876], Fresh[4875], Fresh[4874], Fresh[4873], Fresh[4872], Fresh[4871], Fresh[4870], Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866], Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860], Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854], Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850], Fresh[4849], Fresh[4848], Fresh[4847], Fresh[4846], Fresh[4845], Fresh[4844], Fresh[4843], Fresh[4842], Fresh[4841], Fresh[4840], Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836], Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830], Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824], Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820], Fresh[4819], Fresh[4818], Fresh[4817], Fresh[4816], Fresh[4815], Fresh[4814], Fresh[4813], Fresh[4812], Fresh[4811], Fresh[4810], Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806], Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800], Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794], Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790], Fresh[4789], Fresh[4788], Fresh[4787], Fresh[4786], Fresh[4785], Fresh[4784], Fresh[4783], Fresh[4782], Fresh[4781], Fresh[4780], Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776], Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770], Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764], Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760], Fresh[4759], Fresh[4758], Fresh[4757], Fresh[4756], Fresh[4755], Fresh[4754], Fresh[4753], Fresh[4752], Fresh[4751], Fresh[4750], Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746], Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740], Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734], Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730], Fresh[4729], Fresh[4728], Fresh[4727], Fresh[4726], Fresh[4725], Fresh[4724], Fresh[4723], Fresh[4722], Fresh[4721], Fresh[4720], Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716], Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710], Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704], Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700], Fresh[4699], Fresh[4698], Fresh[4697], Fresh[4696], Fresh[4695], Fresh[4694], Fresh[4693], Fresh[4692], Fresh[4691], Fresh[4690], Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686], Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680], Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674], Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670], Fresh[4669], Fresh[4668], Fresh[4667], Fresh[4666], Fresh[4665], Fresh[4664], Fresh[4663], Fresh[4662], Fresh[4661], Fresh[4660], Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656], Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650], Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644], Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640], Fresh[4639], Fresh[4638], Fresh[4637], Fresh[4636], Fresh[4635], Fresh[4634], Fresh[4633], Fresh[4632], Fresh[4631], Fresh[4630], Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626], Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620], Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614], Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610], Fresh[4609], Fresh[4608], Fresh[4607], Fresh[4606], Fresh[4605], Fresh[4604], Fresh[4603], Fresh[4602], Fresh[4601], Fresh[4600], Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596], Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590], Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584], Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580], Fresh[4579], Fresh[4578], Fresh[4577], Fresh[4576], Fresh[4575], Fresh[4574], Fresh[4573], Fresh[4572], Fresh[4571], Fresh[4570], Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566], Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560], Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554], Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550], Fresh[4549], Fresh[4548], Fresh[4547], Fresh[4546], Fresh[4545], Fresh[4544], Fresh[4543], Fresh[4542], Fresh[4541], Fresh[4540], Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536], Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530], Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524], Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520], Fresh[4519], Fresh[4518], Fresh[4517], Fresh[4516], Fresh[4515], Fresh[4514], Fresh[4513], Fresh[4512], Fresh[4511], Fresh[4510], Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506], Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500], Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494], Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490], Fresh[4489], Fresh[4488], Fresh[4487], Fresh[4486], Fresh[4485], Fresh[4484], Fresh[4483], Fresh[4482], Fresh[4481], Fresh[4480], Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476], Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470], Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464], Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460], Fresh[4459], Fresh[4458], Fresh[4457], Fresh[4456], Fresh[4455], Fresh[4454], Fresh[4453], Fresh[4452], Fresh[4451], Fresh[4450], Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446], Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440], Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434], Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430], Fresh[4429], Fresh[4428], Fresh[4427], Fresh[4426], Fresh[4425], Fresh[4424], Fresh[4423], Fresh[4422], Fresh[4421], Fresh[4420], Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416], Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410], Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404], Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400], Fresh[4399], Fresh[4398], Fresh[4397], Fresh[4396], Fresh[4395], Fresh[4394], Fresh[4393], Fresh[4392], Fresh[4391], Fresh[4390], Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386], Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380], Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374], Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370], Fresh[4369], Fresh[4368], Fresh[4367], Fresh[4366], Fresh[4365], Fresh[4364], Fresh[4363], Fresh[4362], Fresh[4361], Fresh[4360], Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356], Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350], Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344], Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340], Fresh[4339], Fresh[4338], Fresh[4337], Fresh[4336], Fresh[4335], Fresh[4334], Fresh[4333], Fresh[4332], Fresh[4331], Fresh[4330], Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326], Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320], Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314], Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310], Fresh[4309], Fresh[4308], Fresh[4307], Fresh[4306], Fresh[4305], Fresh[4304], Fresh[4303], Fresh[4302], Fresh[4301], Fresh[4300], Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296], Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290], Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284], Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280], Fresh[4279], Fresh[4278], Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272], Fresh[4271], Fresh[4270], Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266], Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260], Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254], Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250], Fresh[4249], Fresh[4248], Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242], Fresh[4241], Fresh[4240], Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236], Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230], Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224], Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220], Fresh[4219], Fresh[4218], Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212], Fresh[4211], Fresh[4210], Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206], Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200], Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194], Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190], Fresh[4189], Fresh[4188], Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182], Fresh[4181], Fresh[4180], Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176], Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170], Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164], Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160], Fresh[4159], Fresh[4158], Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152], Fresh[4151], Fresh[4150], Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146], Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140], Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134], Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130], Fresh[4129], Fresh[4128], Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122], Fresh[4121], Fresh[4120], Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116], Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110], Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104], Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100], Fresh[4099], Fresh[4098], Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092], Fresh[4091], Fresh[4090], Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086], Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080], Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074], Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068], Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062], Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056], Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050], Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044], Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038], Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032], Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026], Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020], Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014], Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008], Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002], Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996], Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990], Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984], Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978], Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972], Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966], Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960], Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954], Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948], Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942], Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936], Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930], Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924], Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918], Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912], Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906], Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900], Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894], Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888], Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882], Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876], Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870], Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864], Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858], Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852], Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846], Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840], Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834], Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828], Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822], Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816], Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810], Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804], Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798], Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792], Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786], Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780], Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774], Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768], Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762], Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756], Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750], Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744], Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738], Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732], Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726], Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720], Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714], Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708], Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702], Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696], Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690], Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684], Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678], Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672], Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666], Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660], Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654], Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648], Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642], Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636], Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630], Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624], Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618], Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612], Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606], Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600], Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594], Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588], Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582], Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576], Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570], Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564], Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558], Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552], Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546], Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540], Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534], Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528], Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522], Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516], Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510], Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504], Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498], Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492], Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486], Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480], Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474], Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468], Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462], Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456], Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450], Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444], Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438], Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432], Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426], Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420], Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414], Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408], Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402], Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396], Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390], Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384], Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378], Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372], Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366], Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360], Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354], Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348], Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342], Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336], Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330], Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324], Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318], Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312], Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306], Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300], Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294], Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288], Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282], Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276], Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270], Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264], Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258], Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252], Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246], Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240], Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234], Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228], Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222], Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216], Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210], Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204], Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198], Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192], Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186], Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180], Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174], Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168], Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162], Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156], Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150], Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144], Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138], Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132], Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126], Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120], Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114], Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108], Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102], Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096], Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090], Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084], Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078], Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072], Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066], Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060], Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054], Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048], Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042], Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036], Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030], Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024], Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018], Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012], Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006], Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000], Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994], Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988], Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982], Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976], Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970], Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964], Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958], Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952], Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946], Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940], Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934], Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928], Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922], Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916], Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910], Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904], Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898], Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892], Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886], Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880], Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874], Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868], Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862], Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856], Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850], Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844], Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838], Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832], Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826], Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820], Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814], Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808], Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802], Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796], Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790], Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784], Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778], Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772], Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766], Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760], Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754], Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748], Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742], Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736], Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730], Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724], Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718], Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712], Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706], Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700], Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694], Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688], Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682], Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676], Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670], Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664], Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658], Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652], Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646], Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640], Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634], Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628], Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622], Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616], Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610], Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604], Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598], Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592], Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586], Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580], Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574], Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568], Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562], Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556], Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550], Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544], Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532], Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520], Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508], Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496], Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490], Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484], Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472], Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460], Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448], Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436], Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430], Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424], Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412], Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400], Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388], Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376], Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370], Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364], Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352], Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340], Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328], Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316], Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310], Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304], Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292], Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280], Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268], Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256], Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250], Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244], Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232], Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220], Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208], Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196], Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190], Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184], Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172], Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160], Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148], Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136], Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130], Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124], Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112], Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100], Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088], Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076], Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070], Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064], Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052], Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040], Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028], Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016], Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010], Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004], Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992], Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980], Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968], Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956], Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950], Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944], Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932], Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920], Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908], Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896], Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890], Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884], Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872], Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860], Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848], Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836], Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830], Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824], Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812], Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800], Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788], Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776], Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770], Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764], Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752], Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740], Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728], Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716], Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710], Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704], Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692], Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680], Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668], Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656], Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650], Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644], Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632], Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620], Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608], Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596], Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590], Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584], Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572], Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560], Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548], Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536], Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530], Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524], Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512], Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500], Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488], Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476], Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470], Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464], Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452], Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440], Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428], Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416], Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410], Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404], Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392], Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380], Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368], Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356], Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350], Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344], Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332], Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320], Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308], Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296], Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290], Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284], Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272], Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260], Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248], Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236], Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230], Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224], Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212], Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200], Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188], Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176], Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170], Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164], Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152], Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140], Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128], Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116], Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110], Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104], Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092], Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080], Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068], Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056], Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050], Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044], Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032], Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020], Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960], Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900], Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840], Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780], Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720], Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660], Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600], Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540], Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480], Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420], Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360], Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300], Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240], Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180], Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_4548, signal_4547, signal_4546, signal_4545, signal_4544, signal_4543, signal_4542, signal_4541, signal_4540, signal_4539, signal_4538, signal_4537, signal_4536, signal_4535, signal_4534, signal_4533, signal_4532, signal_4531, signal_4530, signal_4529, signal_4528, signal_4527, signal_4526, signal_4525, signal_4516, signal_4514, signal_4511, signal_4510, signal_4509, signal_4508, signal_4506, signal_4503, signal_4502, signal_4501, signal_4500, signal_4498, signal_4495, signal_4494, signal_4493, signal_4492, signal_4490, signal_4487, signal_4486, signal_4485, signal_4484, signal_4482, signal_4479, signal_4478, signal_4477, signal_4476, signal_4474, signal_4471, signal_4470, signal_4469, signal_4468, signal_4466, signal_4463, signal_4462, signal_4461, signal_4460, signal_4458, signal_4455, signal_4454, signal_4453, signal_4452, signal_4450, signal_4447, signal_4446, signal_4445, signal_4444, signal_4442, signal_4439, signal_4438, signal_4437, signal_4436, signal_4434, signal_4431, signal_4430, signal_4429, signal_4428, signal_4426, signal_4423, signal_4422, signal_4421, signal_4420, signal_4418, signal_4415, signal_4414, signal_4413, signal_4412, signal_4410, signal_4407, signal_4406, signal_4405, signal_4404, signal_4402, signal_4399, signal_4398, signal_4397, signal_4396, signal_4394, signal_4391, signal_4390, signal_4389, signal_4121, signal_4120, signal_4119, signal_4118, signal_4117, signal_4116, signal_4115, signal_4114, signal_4112, signal_4111, signal_4110, signal_4109, signal_4108, signal_4107, signal_4106, signal_4105, signal_4104, signal_4103, signal_4102, signal_4101, signal_4100, signal_4099, signal_4098, signal_4097, signal_4096, signal_4095, signal_4094, signal_4093, signal_4092, signal_4091, signal_4089, signal_4088, signal_4087, signal_4086, signal_4085, signal_4084, signal_4083, signal_4082, signal_4080, signal_4079, signal_4078, signal_4077, signal_4076, signal_4075, signal_4074, signal_4073, signal_4072, signal_4071, signal_4070, signal_4069, signal_4068, signal_4067, signal_4066, signal_4065, signal_4064, signal_4063, signal_4062, signal_4061, signal_4060, signal_4059, signal_4057, signal_4056, signal_4055, signal_4054, signal_4053, signal_4052, signal_4051, signal_4050, signal_4048, signal_4047, signal_4046, signal_4045, signal_4044, signal_4043, signal_4042, signal_4041, signal_4040, signal_4039, signal_4038, signal_4037, signal_4036, signal_4035, signal_4034, signal_4033, signal_4032, signal_4031, signal_4030, signal_4029, signal_4028, signal_4027, signal_4025, signal_4024, signal_4023, signal_4022, signal_4021, signal_4020, signal_4019, signal_4018, signal_4016, signal_4015, signal_4014, signal_4013, signal_4012, signal_4011, signal_4010, signal_4009, signal_4008, signal_4007, signal_4006, signal_4005, signal_4004, signal_4003, signal_4002, signal_4001, signal_4000, signal_3999, signal_3998, signal_3997, signal_3996, signal_3995, signal_3994, signal_3992, signal_3991, signal_3986, signal_3984, signal_3983, signal_3978, signal_3976, signal_3975, signal_3970, signal_3968, signal_3967, signal_3962, signal_3960, signal_3959, signal_3954, signal_3952, signal_3951, signal_3946, signal_3944, signal_3943, signal_3938, signal_3936, signal_3935, signal_3930, signal_3928, signal_3927, signal_3922, signal_3920, signal_3919, signal_3914, signal_3912, signal_3911, signal_3906, signal_3904, signal_3903, signal_3898, signal_3896, signal_3895, signal_3890, signal_3888, signal_3887, signal_3882, signal_3880, signal_3879, signal_3874, signal_3872, signal_3871, signal_3116, signal_3115, signal_3114, signal_3113, signal_3112, signal_3111, signal_3110, signal_3109, signal_2852, signal_2789, signal_2788, signal_2725, signal_2724, signal_2661, signal_2660, signal_2597}), .out1 ({signal_5236, signal_5235, signal_5234, signal_5233, signal_5232, signal_5231, signal_5230, signal_5229, signal_5228, signal_5227, signal_5226, signal_5225, signal_5224, signal_5223, signal_5222, signal_5221, signal_5220, signal_5219, signal_5218, signal_5217, signal_5216, signal_5215, signal_5214, signal_5213, signal_5212, signal_5211, signal_5210, signal_5209, signal_5208, signal_5207, signal_5206, signal_5205, signal_5204, signal_5203, signal_5202, signal_5201, signal_5200, signal_5199, signal_5198, signal_5197, signal_5196, signal_5195, signal_5194, signal_5193, signal_5192, signal_5191, signal_5190, signal_5189, signal_5188, signal_5187, signal_5186, signal_5185, signal_5184, signal_5183, signal_5182, signal_5181, signal_5180, signal_5179, signal_5178, signal_5177, signal_5176, signal_5175, signal_5174, signal_5173, signal_5172, signal_5171, signal_5170, signal_5169, signal_5168, signal_5167, signal_5166, signal_5165, signal_5164, signal_5163, signal_5162, signal_5161, signal_5160, signal_5159, signal_5158, signal_5157, signal_5156, signal_5155, signal_5154, signal_5153, signal_5152, signal_5151, signal_5150, signal_5149, signal_5148, signal_5147, signal_5146, signal_5145, signal_5144, signal_5143, signal_5142, signal_5141, signal_5140, signal_5139, signal_5138, signal_5137, signal_5136, signal_5135, signal_5134, signal_5133, signal_5132, signal_5131, signal_5130, signal_5129, signal_5128, signal_5127, signal_5126, signal_5125, signal_5124, signal_5123, signal_5122, signal_5121, signal_5120, signal_5119, signal_5118, signal_5117, signal_5116, signal_5115, signal_5114, signal_5113, signal_5112, signal_5111, signal_5110, signal_5109, signal_5108, signal_5107, signal_5106, signal_5105, signal_5104, signal_5103, signal_5102, signal_5101, signal_5100, signal_5099, signal_5098, signal_5097, signal_5096, signal_5095, signal_5094, signal_5093, signal_5092, signal_5091, signal_5090, signal_5089, signal_5088, signal_5087, signal_5086, signal_5085, signal_5084, signal_5083, signal_5082, signal_5081, signal_5080, signal_5079, signal_5078, signal_5077, signal_5076, signal_5075, signal_5074, signal_5073, signal_5072, signal_5071, signal_5070, signal_5069, signal_5068, signal_5067, signal_5066, signal_5065, signal_5064, signal_5063, signal_5062, signal_5061, signal_5060, signal_5059, signal_5058, signal_5057, signal_5056, signal_5055, signal_5054, signal_5053, signal_5052, signal_5051, signal_5050, signal_5049, signal_5048, signal_5047, signal_5046, signal_5045, signal_5044, signal_5043, signal_5042, signal_5041, signal_5040, signal_5039, signal_5038, signal_5037, signal_5036, signal_5035, signal_5034, signal_5033, signal_5032, signal_5031, signal_5030, signal_5029, signal_5028, signal_5027, signal_5026, signal_5025, signal_5024, signal_5023, signal_5022, signal_5021, signal_5020, signal_5019, signal_5018, signal_5017, signal_5016, signal_5015, signal_5014, signal_5013, signal_5012, signal_5011, signal_5010, signal_5009, signal_5008, signal_5007, signal_5006, signal_5005, signal_5004, signal_5003, signal_5002, signal_5001, signal_5000, signal_4999, signal_4998, signal_4997, signal_4996, signal_4995, signal_4994, signal_4993, signal_4992, signal_4991, signal_4990, signal_4989, signal_4988, signal_4987, signal_4986, signal_4985, signal_4984, signal_4983, signal_4982, signal_4981, signal_4980, signal_4979, signal_4978, signal_4977, signal_4976, signal_4975, signal_4974, signal_4973, signal_4972, signal_4971, signal_4970, signal_4969, signal_4968, signal_4967, signal_4966, signal_4965, signal_4964, signal_4963, signal_4962, signal_4961, signal_4960, signal_4959, signal_4958, signal_4957, signal_4956, signal_4955, signal_4954, signal_4953, signal_4952, signal_4951, signal_4950, signal_4949}) ) ;

    /* register cells */
    reg_masked #(.low_latency(1), .pipeline(0)) cell_293 ( .clk (signal_46981), .D ({signal_5478, signal_421}), .Q ({signal_4549, signal_3870}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_296 ( .clk (signal_46981), .D ({signal_5480, signal_423}), .Q ({signal_4666, signal_3869}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_299 ( .clk (signal_46981), .D ({signal_5482, signal_425}), .Q ({signal_4699, signal_3868}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_302 ( .clk (signal_46981), .D ({signal_5484, signal_427}), .Q ({signal_4732, signal_3867}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_305 ( .clk (signal_46981), .D ({signal_5486, signal_429}), .Q ({signal_4765, signal_3866}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_308 ( .clk (signal_46981), .D ({signal_5488, signal_431}), .Q ({signal_4798, signal_3865}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_311 ( .clk (signal_46981), .D ({signal_5490, signal_433}), .Q ({signal_4831, signal_3864}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_314 ( .clk (signal_46981), .D ({signal_5492, signal_435}), .Q ({signal_4864, signal_3863}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_317 ( .clk (signal_46981), .D ({signal_5494, signal_437}), .Q ({signal_4897, signal_3862}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_320 ( .clk (signal_46981), .D ({signal_5496, signal_439}), .Q ({signal_4930, signal_3861}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_323 ( .clk (signal_46981), .D ({signal_5498, signal_441}), .Q ({signal_4582, signal_3860}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_326 ( .clk (signal_46981), .D ({signal_5500, signal_443}), .Q ({signal_4615, signal_3859}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_329 ( .clk (signal_46981), .D ({signal_5502, signal_445}), .Q ({signal_4642, signal_3858}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_332 ( .clk (signal_46981), .D ({signal_5504, signal_447}), .Q ({signal_4645, signal_3857}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_335 ( .clk (signal_46981), .D ({signal_5506, signal_449}), .Q ({signal_4648, signal_3856}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_338 ( .clk (signal_46981), .D ({signal_5508, signal_451}), .Q ({signal_4651, signal_3855}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_341 ( .clk (signal_46981), .D ({signal_5510, signal_453}), .Q ({signal_4654, signal_3854}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_344 ( .clk (signal_46981), .D ({signal_5512, signal_455}), .Q ({signal_4657, signal_3853}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_347 ( .clk (signal_46981), .D ({signal_5514, signal_457}), .Q ({signal_4660, signal_3852}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_350 ( .clk (signal_46981), .D ({signal_5516, signal_459}), .Q ({signal_4663, signal_3851}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_353 ( .clk (signal_46981), .D ({signal_5518, signal_461}), .Q ({signal_4669, signal_3850}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_356 ( .clk (signal_46981), .D ({signal_5520, signal_463}), .Q ({signal_4672, signal_3849}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_359 ( .clk (signal_46981), .D ({signal_5522, signal_465}), .Q ({signal_4675, signal_3848}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_362 ( .clk (signal_46981), .D ({signal_5524, signal_467}), .Q ({signal_4678, signal_3847}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_365 ( .clk (signal_46981), .D ({signal_5526, signal_469}), .Q ({signal_4681, signal_3846}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_368 ( .clk (signal_46981), .D ({signal_5528, signal_471}), .Q ({signal_4684, signal_3845}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_371 ( .clk (signal_46981), .D ({signal_5530, signal_473}), .Q ({signal_4687, signal_3844}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_374 ( .clk (signal_46981), .D ({signal_5532, signal_475}), .Q ({signal_4690, signal_3843}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_377 ( .clk (signal_46981), .D ({signal_5534, signal_477}), .Q ({signal_4693, signal_3842}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_380 ( .clk (signal_46981), .D ({signal_5536, signal_479}), .Q ({signal_4696, signal_3841}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_383 ( .clk (signal_46981), .D ({signal_5538, signal_481}), .Q ({signal_4702, signal_3840}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_386 ( .clk (signal_46981), .D ({signal_5540, signal_483}), .Q ({signal_4705, signal_3839}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_389 ( .clk (signal_46981), .D ({signal_5542, signal_485}), .Q ({signal_4708, signal_3838}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_392 ( .clk (signal_46981), .D ({signal_5544, signal_487}), .Q ({signal_4711, signal_3837}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_395 ( .clk (signal_46981), .D ({signal_5546, signal_489}), .Q ({signal_4714, signal_3836}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_398 ( .clk (signal_46981), .D ({signal_5548, signal_491}), .Q ({signal_4717, signal_3835}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_401 ( .clk (signal_46981), .D ({signal_5550, signal_493}), .Q ({signal_4720, signal_3834}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_404 ( .clk (signal_46981), .D ({signal_5552, signal_495}), .Q ({signal_4723, signal_3833}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_407 ( .clk (signal_46981), .D ({signal_5554, signal_497}), .Q ({signal_4726, signal_3832}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_410 ( .clk (signal_46981), .D ({signal_5556, signal_499}), .Q ({signal_4729, signal_3831}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_413 ( .clk (signal_46981), .D ({signal_5558, signal_501}), .Q ({signal_4735, signal_3830}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_416 ( .clk (signal_46981), .D ({signal_5560, signal_503}), .Q ({signal_4738, signal_3829}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_419 ( .clk (signal_46981), .D ({signal_5562, signal_505}), .Q ({signal_4741, signal_3828}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_422 ( .clk (signal_46981), .D ({signal_5564, signal_507}), .Q ({signal_4744, signal_3827}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_425 ( .clk (signal_46981), .D ({signal_5566, signal_509}), .Q ({signal_4747, signal_3826}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_428 ( .clk (signal_46981), .D ({signal_5568, signal_511}), .Q ({signal_4750, signal_3825}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_431 ( .clk (signal_46981), .D ({signal_5570, signal_513}), .Q ({signal_4753, signal_3824}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_434 ( .clk (signal_46981), .D ({signal_5572, signal_515}), .Q ({signal_4756, signal_3823}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_437 ( .clk (signal_46981), .D ({signal_5574, signal_517}), .Q ({signal_4759, signal_3822}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_440 ( .clk (signal_46981), .D ({signal_5576, signal_519}), .Q ({signal_4762, signal_3821}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_443 ( .clk (signal_46981), .D ({signal_5578, signal_521}), .Q ({signal_4768, signal_3820}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_446 ( .clk (signal_46981), .D ({signal_5580, signal_523}), .Q ({signal_4771, signal_3819}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_449 ( .clk (signal_46981), .D ({signal_5582, signal_525}), .Q ({signal_4774, signal_3818}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_452 ( .clk (signal_46981), .D ({signal_5584, signal_527}), .Q ({signal_4777, signal_3817}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_455 ( .clk (signal_46981), .D ({signal_5586, signal_529}), .Q ({signal_4780, signal_3816}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_458 ( .clk (signal_46981), .D ({signal_5588, signal_531}), .Q ({signal_4783, signal_3815}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_461 ( .clk (signal_46981), .D ({signal_5590, signal_533}), .Q ({signal_4786, signal_3814}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_464 ( .clk (signal_46981), .D ({signal_5592, signal_535}), .Q ({signal_4789, signal_3813}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_467 ( .clk (signal_46981), .D ({signal_5594, signal_537}), .Q ({signal_4792, signal_3812}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_470 ( .clk (signal_46981), .D ({signal_5596, signal_539}), .Q ({signal_4795, signal_3811}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_473 ( .clk (signal_46981), .D ({signal_5598, signal_541}), .Q ({signal_4801, signal_3810}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_476 ( .clk (signal_46981), .D ({signal_5600, signal_543}), .Q ({signal_4804, signal_3809}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_479 ( .clk (signal_46981), .D ({signal_5602, signal_545}), .Q ({signal_4807, signal_3808}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_482 ( .clk (signal_46981), .D ({signal_5604, signal_547}), .Q ({signal_4810, signal_3807}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_485 ( .clk (signal_46981), .D ({signal_5606, signal_549}), .Q ({signal_4813, signal_3806}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_488 ( .clk (signal_46981), .D ({signal_5608, signal_551}), .Q ({signal_4816, signal_3805}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_491 ( .clk (signal_46981), .D ({signal_5610, signal_553}), .Q ({signal_4819, signal_3804}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_494 ( .clk (signal_46981), .D ({signal_5612, signal_555}), .Q ({signal_4822, signal_3803}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_497 ( .clk (signal_46981), .D ({signal_5614, signal_557}), .Q ({signal_4825, signal_3802}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_500 ( .clk (signal_46981), .D ({signal_5616, signal_559}), .Q ({signal_4828, signal_3801}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_503 ( .clk (signal_46981), .D ({signal_5618, signal_561}), .Q ({signal_4834, signal_3800}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_506 ( .clk (signal_46981), .D ({signal_5620, signal_563}), .Q ({signal_4837, signal_3799}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_509 ( .clk (signal_46981), .D ({signal_5622, signal_565}), .Q ({signal_4840, signal_3798}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_512 ( .clk (signal_46981), .D ({signal_5624, signal_567}), .Q ({signal_4843, signal_3797}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_515 ( .clk (signal_46981), .D ({signal_5626, signal_569}), .Q ({signal_4846, signal_3796}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_518 ( .clk (signal_46981), .D ({signal_5628, signal_571}), .Q ({signal_4849, signal_3795}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_521 ( .clk (signal_46981), .D ({signal_5630, signal_573}), .Q ({signal_4852, signal_3794}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_524 ( .clk (signal_46981), .D ({signal_5632, signal_575}), .Q ({signal_4855, signal_3793}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_527 ( .clk (signal_46981), .D ({signal_5634, signal_577}), .Q ({signal_4858, signal_3792}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_530 ( .clk (signal_46981), .D ({signal_5636, signal_579}), .Q ({signal_4861, signal_3791}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_533 ( .clk (signal_46981), .D ({signal_5638, signal_581}), .Q ({signal_4867, signal_3790}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_536 ( .clk (signal_46981), .D ({signal_5640, signal_583}), .Q ({signal_4870, signal_3789}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_539 ( .clk (signal_46981), .D ({signal_5642, signal_585}), .Q ({signal_4873, signal_3788}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_542 ( .clk (signal_46981), .D ({signal_5644, signal_587}), .Q ({signal_4876, signal_3787}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_545 ( .clk (signal_46981), .D ({signal_5646, signal_589}), .Q ({signal_4879, signal_3786}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_548 ( .clk (signal_46981), .D ({signal_5648, signal_591}), .Q ({signal_4882, signal_3785}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_551 ( .clk (signal_46981), .D ({signal_5650, signal_593}), .Q ({signal_4885, signal_3784}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_554 ( .clk (signal_46981), .D ({signal_5652, signal_595}), .Q ({signal_4888, signal_3783}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_557 ( .clk (signal_46981), .D ({signal_5654, signal_597}), .Q ({signal_4891, signal_3782}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_560 ( .clk (signal_46981), .D ({signal_5656, signal_599}), .Q ({signal_4894, signal_3781}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_563 ( .clk (signal_46981), .D ({signal_5658, signal_601}), .Q ({signal_4900, signal_3780}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_566 ( .clk (signal_46981), .D ({signal_5660, signal_603}), .Q ({signal_4903, signal_3779}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_569 ( .clk (signal_46981), .D ({signal_5662, signal_605}), .Q ({signal_4906, signal_3778}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_572 ( .clk (signal_46981), .D ({signal_5664, signal_607}), .Q ({signal_4909, signal_3777}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_575 ( .clk (signal_46981), .D ({signal_5666, signal_609}), .Q ({signal_4912, signal_3776}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_578 ( .clk (signal_46981), .D ({signal_5668, signal_611}), .Q ({signal_4915, signal_3775}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_581 ( .clk (signal_46981), .D ({signal_5670, signal_613}), .Q ({signal_4918, signal_3774}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_584 ( .clk (signal_46981), .D ({signal_5672, signal_615}), .Q ({signal_4921, signal_3773}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_587 ( .clk (signal_46981), .D ({signal_5674, signal_617}), .Q ({signal_4924, signal_3772}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_590 ( .clk (signal_46981), .D ({signal_5676, signal_619}), .Q ({signal_4927, signal_3771}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_593 ( .clk (signal_46981), .D ({signal_5678, signal_621}), .Q ({signal_4552, signal_3770}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_596 ( .clk (signal_46981), .D ({signal_5680, signal_623}), .Q ({signal_4555, signal_3769}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_599 ( .clk (signal_46981), .D ({signal_5682, signal_625}), .Q ({signal_4558, signal_3768}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_602 ( .clk (signal_46981), .D ({signal_5684, signal_627}), .Q ({signal_4561, signal_3767}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_605 ( .clk (signal_46981), .D ({signal_5686, signal_629}), .Q ({signal_4564, signal_3766}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_608 ( .clk (signal_46981), .D ({signal_5688, signal_631}), .Q ({signal_4567, signal_3765}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_611 ( .clk (signal_46981), .D ({signal_5690, signal_633}), .Q ({signal_4570, signal_3764}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_614 ( .clk (signal_46981), .D ({signal_5692, signal_635}), .Q ({signal_4573, signal_3763}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_617 ( .clk (signal_46981), .D ({signal_5694, signal_637}), .Q ({signal_4576, signal_3762}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_620 ( .clk (signal_46981), .D ({signal_5696, signal_639}), .Q ({signal_4579, signal_3761}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_623 ( .clk (signal_46981), .D ({signal_5698, signal_641}), .Q ({signal_4585, signal_3760}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_626 ( .clk (signal_46981), .D ({signal_5700, signal_643}), .Q ({signal_4588, signal_3759}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_629 ( .clk (signal_46981), .D ({signal_5702, signal_645}), .Q ({signal_4591, signal_3758}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_632 ( .clk (signal_46981), .D ({signal_5704, signal_647}), .Q ({signal_4594, signal_3757}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_635 ( .clk (signal_46981), .D ({signal_5706, signal_649}), .Q ({signal_4597, signal_3756}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_638 ( .clk (signal_46981), .D ({signal_5708, signal_651}), .Q ({signal_4600, signal_3755}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_641 ( .clk (signal_46981), .D ({signal_5710, signal_653}), .Q ({signal_4603, signal_3754}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_644 ( .clk (signal_46981), .D ({signal_5712, signal_655}), .Q ({signal_4606, signal_3753}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_647 ( .clk (signal_46981), .D ({signal_5714, signal_657}), .Q ({signal_4609, signal_3752}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_650 ( .clk (signal_46981), .D ({signal_5716, signal_659}), .Q ({signal_4612, signal_3751}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_653 ( .clk (signal_46981), .D ({signal_5718, signal_661}), .Q ({signal_4618, signal_3750}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_656 ( .clk (signal_46981), .D ({signal_5720, signal_663}), .Q ({signal_4621, signal_3749}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_659 ( .clk (signal_46981), .D ({signal_5722, signal_665}), .Q ({signal_4624, signal_3748}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_662 ( .clk (signal_46981), .D ({signal_5724, signal_667}), .Q ({signal_4627, signal_3747}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_665 ( .clk (signal_46981), .D ({signal_5726, signal_669}), .Q ({signal_4630, signal_3746}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_668 ( .clk (signal_46981), .D ({signal_5728, signal_671}), .Q ({signal_4633, signal_3745}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_671 ( .clk (signal_46981), .D ({signal_5730, signal_673}), .Q ({signal_4636, signal_3744}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_674 ( .clk (signal_46981), .D ({signal_5732, signal_675}), .Q ({signal_4639, signal_3743}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3157 ( .clk (signal_46981), .D ({signal_5910, signal_2853}), .Q ({signal_4550, signal_4378}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3160 ( .clk (signal_46981), .D ({signal_5912, signal_2855}), .Q ({signal_4667, signal_4377}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3163 ( .clk (signal_46981), .D ({signal_5914, signal_2857}), .Q ({signal_4700, signal_4376}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3166 ( .clk (signal_46981), .D ({signal_5916, signal_2859}), .Q ({signal_4733, signal_4375}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3169 ( .clk (signal_46981), .D ({signal_5918, signal_2861}), .Q ({signal_4766, signal_4374}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3172 ( .clk (signal_46981), .D ({signal_5920, signal_2863}), .Q ({signal_4799, signal_4373}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3175 ( .clk (signal_46981), .D ({signal_5922, signal_2865}), .Q ({signal_4832, signal_4372}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3178 ( .clk (signal_46981), .D ({signal_5924, signal_2867}), .Q ({signal_4865, signal_4371}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3181 ( .clk (signal_46981), .D ({signal_5926, signal_2869}), .Q ({signal_4898, signal_4370}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3184 ( .clk (signal_46981), .D ({signal_5928, signal_2871}), .Q ({signal_4931, signal_4369}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3187 ( .clk (signal_46981), .D ({signal_5930, signal_2873}), .Q ({signal_4583, signal_4368}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3190 ( .clk (signal_46981), .D ({signal_5932, signal_2875}), .Q ({signal_4616, signal_4367}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3193 ( .clk (signal_46981), .D ({signal_5934, signal_2877}), .Q ({signal_4643, signal_4366}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3196 ( .clk (signal_46981), .D ({signal_5936, signal_2879}), .Q ({signal_4646, signal_4365}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3199 ( .clk (signal_46981), .D ({signal_5938, signal_2881}), .Q ({signal_4649, signal_4364}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3202 ( .clk (signal_46981), .D ({signal_5940, signal_2883}), .Q ({signal_4652, signal_4363}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3205 ( .clk (signal_46981), .D ({signal_5942, signal_2885}), .Q ({signal_4655, signal_4362}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3208 ( .clk (signal_46981), .D ({signal_5944, signal_2887}), .Q ({signal_4658, signal_4361}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3211 ( .clk (signal_46981), .D ({signal_5946, signal_2889}), .Q ({signal_4661, signal_4360}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3214 ( .clk (signal_46981), .D ({signal_5948, signal_2891}), .Q ({signal_4664, signal_4359}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3217 ( .clk (signal_46981), .D ({signal_5950, signal_2893}), .Q ({signal_4670, signal_4358}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3220 ( .clk (signal_46981), .D ({signal_5952, signal_2895}), .Q ({signal_4673, signal_4357}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3223 ( .clk (signal_46981), .D ({signal_5954, signal_2897}), .Q ({signal_4676, signal_4356}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3226 ( .clk (signal_46981), .D ({signal_5956, signal_2899}), .Q ({signal_4679, signal_4355}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3229 ( .clk (signal_46981), .D ({signal_5982, signal_2901}), .Q ({signal_4682, signal_4354}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3232 ( .clk (signal_46981), .D ({signal_5984, signal_2903}), .Q ({signal_4685, signal_4353}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3235 ( .clk (signal_46981), .D ({signal_6016, signal_2905}), .Q ({signal_4688, signal_4352}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3238 ( .clk (signal_46981), .D ({signal_6018, signal_2907}), .Q ({signal_4691, signal_4351}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3241 ( .clk (signal_46981), .D ({signal_6003, signal_2909}), .Q ({signal_4694, signal_4350}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3244 ( .clk (signal_46981), .D ({signal_6020, signal_2911}), .Q ({signal_4697, signal_4349}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3247 ( .clk (signal_46981), .D ({signal_5986, signal_2913}), .Q ({signal_4703, signal_4348}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3250 ( .clk (signal_46981), .D ({signal_6005, signal_2915}), .Q ({signal_4706, signal_4347}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3253 ( .clk (signal_46981), .D ({signal_5820, signal_2917}), .Q ({signal_4709, signal_4346}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3256 ( .clk (signal_46981), .D ({signal_5822, signal_2919}), .Q ({signal_4712, signal_4345}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3259 ( .clk (signal_46981), .D ({signal_5824, signal_2921}), .Q ({signal_4715, signal_4344}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3262 ( .clk (signal_46981), .D ({signal_5826, signal_2923}), .Q ({signal_4718, signal_4343}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3265 ( .clk (signal_46981), .D ({signal_5828, signal_2925}), .Q ({signal_4721, signal_4342}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3268 ( .clk (signal_46981), .D ({signal_5830, signal_2927}), .Q ({signal_4724, signal_4341}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3271 ( .clk (signal_46981), .D ({signal_5832, signal_2929}), .Q ({signal_4727, signal_4340}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3274 ( .clk (signal_46981), .D ({signal_5834, signal_2931}), .Q ({signal_4730, signal_4339}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3277 ( .clk (signal_46981), .D ({signal_5836, signal_2933}), .Q ({signal_4736, signal_4338}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3280 ( .clk (signal_46981), .D ({signal_5838, signal_2935}), .Q ({signal_4739, signal_4337}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3283 ( .clk (signal_46981), .D ({signal_5840, signal_2937}), .Q ({signal_4742, signal_4336}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3286 ( .clk (signal_46981), .D ({signal_5842, signal_2939}), .Q ({signal_4745, signal_4335}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3289 ( .clk (signal_46981), .D ({signal_5844, signal_2941}), .Q ({signal_4748, signal_4334}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3292 ( .clk (signal_46981), .D ({signal_5846, signal_2943}), .Q ({signal_4751, signal_4333}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3295 ( .clk (signal_46981), .D ({signal_5848, signal_2945}), .Q ({signal_4754, signal_4332}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3298 ( .clk (signal_46981), .D ({signal_5850, signal_2947}), .Q ({signal_4757, signal_4331}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3301 ( .clk (signal_46981), .D ({signal_5852, signal_2949}), .Q ({signal_4760, signal_4330}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3304 ( .clk (signal_46981), .D ({signal_5854, signal_2951}), .Q ({signal_4763, signal_4329}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3307 ( .clk (signal_46981), .D ({signal_5856, signal_2953}), .Q ({signal_4769, signal_4328}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3310 ( .clk (signal_46981), .D ({signal_5858, signal_2955}), .Q ({signal_4772, signal_4327}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3313 ( .clk (signal_46981), .D ({signal_5860, signal_2957}), .Q ({signal_4775, signal_4326}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3316 ( .clk (signal_46981), .D ({signal_5862, signal_2959}), .Q ({signal_4778, signal_4325}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3319 ( .clk (signal_46981), .D ({signal_5864, signal_2961}), .Q ({signal_4781, signal_4324}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3322 ( .clk (signal_46981), .D ({signal_5866, signal_2963}), .Q ({signal_4784, signal_4323}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3325 ( .clk (signal_46981), .D ({signal_5958, signal_2965}), .Q ({signal_4787, signal_4322}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3328 ( .clk (signal_46981), .D ({signal_5960, signal_2967}), .Q ({signal_4790, signal_4321}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3331 ( .clk (signal_46981), .D ({signal_6007, signal_2969}), .Q ({signal_4793, signal_4320}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3334 ( .clk (signal_46981), .D ({signal_6009, signal_2971}), .Q ({signal_4796, signal_4319}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3337 ( .clk (signal_46981), .D ({signal_5988, signal_2973}), .Q ({signal_4802, signal_4318}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3340 ( .clk (signal_46981), .D ({signal_6011, signal_2975}), .Q ({signal_4805, signal_4317}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3343 ( .clk (signal_46981), .D ({signal_5962, signal_2977}), .Q ({signal_4808, signal_4316}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3346 ( .clk (signal_46981), .D ({signal_5990, signal_2979}), .Q ({signal_4811, signal_4315}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3349 ( .clk (signal_46981), .D ({signal_5734, signal_2981}), .Q ({signal_4814, signal_4314}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3352 ( .clk (signal_46981), .D ({signal_5736, signal_2983}), .Q ({signal_4817, signal_4313}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3355 ( .clk (signal_46981), .D ({signal_5738, signal_2985}), .Q ({signal_4820, signal_4312}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3358 ( .clk (signal_46981), .D ({signal_5740, signal_2987}), .Q ({signal_4823, signal_4311}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3361 ( .clk (signal_46981), .D ({signal_5742, signal_2989}), .Q ({signal_4826, signal_4310}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3364 ( .clk (signal_46981), .D ({signal_5744, signal_2991}), .Q ({signal_4829, signal_4309}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3367 ( .clk (signal_46981), .D ({signal_5746, signal_2993}), .Q ({signal_4835, signal_4308}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3370 ( .clk (signal_46981), .D ({signal_5748, signal_2995}), .Q ({signal_4838, signal_4307}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3373 ( .clk (signal_46981), .D ({signal_5750, signal_2997}), .Q ({signal_4841, signal_4306}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3376 ( .clk (signal_46981), .D ({signal_5752, signal_2999}), .Q ({signal_4844, signal_4305}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3379 ( .clk (signal_46981), .D ({signal_5754, signal_3001}), .Q ({signal_4847, signal_4304}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3382 ( .clk (signal_46981), .D ({signal_5756, signal_3003}), .Q ({signal_4850, signal_4303}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3385 ( .clk (signal_46981), .D ({signal_5758, signal_3005}), .Q ({signal_4853, signal_4302}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3388 ( .clk (signal_46981), .D ({signal_5760, signal_3007}), .Q ({signal_4856, signal_4301}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3391 ( .clk (signal_46981), .D ({signal_5762, signal_3009}), .Q ({signal_4859, signal_4300}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3394 ( .clk (signal_46981), .D ({signal_5764, signal_3011}), .Q ({signal_4862, signal_4299}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3397 ( .clk (signal_46981), .D ({signal_5766, signal_3013}), .Q ({signal_4868, signal_4298}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3400 ( .clk (signal_46981), .D ({signal_5768, signal_3015}), .Q ({signal_4871, signal_4297}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3403 ( .clk (signal_46981), .D ({signal_5770, signal_3017}), .Q ({signal_4874, signal_4296}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3406 ( .clk (signal_46981), .D ({signal_5772, signal_3019}), .Q ({signal_4877, signal_4295}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3409 ( .clk (signal_46981), .D ({signal_5774, signal_3021}), .Q ({signal_4880, signal_4294}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3412 ( .clk (signal_46981), .D ({signal_5776, signal_3023}), .Q ({signal_4883, signal_4293}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3415 ( .clk (signal_46981), .D ({signal_5778, signal_3025}), .Q ({signal_4886, signal_4292}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3418 ( .clk (signal_46981), .D ({signal_5780, signal_3027}), .Q ({signal_4889, signal_4291}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3421 ( .clk (signal_46981), .D ({signal_5868, signal_3029}), .Q ({signal_4892, signal_4290}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3424 ( .clk (signal_46981), .D ({signal_5870, signal_3031}), .Q ({signal_4895, signal_4289}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3427 ( .clk (signal_46981), .D ({signal_5992, signal_3033}), .Q ({signal_4901, signal_4288}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3430 ( .clk (signal_46981), .D ({signal_5994, signal_3035}), .Q ({signal_4904, signal_4287}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3433 ( .clk (signal_46981), .D ({signal_5964, signal_3037}), .Q ({signal_4907, signal_4286}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3436 ( .clk (signal_46981), .D ({signal_5996, signal_3039}), .Q ({signal_4910, signal_4285}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3439 ( .clk (signal_46981), .D ({signal_5872, signal_3041}), .Q ({signal_4913, signal_4284}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3442 ( .clk (signal_46981), .D ({signal_5966, signal_3043}), .Q ({signal_4916, signal_4283}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3445 ( .clk (signal_46981), .D ({signal_5401, signal_3045}), .Q ({signal_4919, signal_4282}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3448 ( .clk (signal_46981), .D ({signal_5403, signal_3047}), .Q ({signal_4922, signal_4281}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3451 ( .clk (signal_46981), .D ({signal_5405, signal_3049}), .Q ({signal_4925, signal_4280}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3454 ( .clk (signal_46981), .D ({signal_5407, signal_3051}), .Q ({signal_4928, signal_4279}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3457 ( .clk (signal_46981), .D ({signal_5409, signal_3053}), .Q ({signal_4553, signal_4278}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3460 ( .clk (signal_46981), .D ({signal_5411, signal_3055}), .Q ({signal_4556, signal_4277}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3463 ( .clk (signal_46981), .D ({signal_5413, signal_3057}), .Q ({signal_4559, signal_4276}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3466 ( .clk (signal_46981), .D ({signal_5415, signal_3059}), .Q ({signal_4562, signal_4275}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3469 ( .clk (signal_46981), .D ({signal_5417, signal_3061}), .Q ({signal_4565, signal_4274}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3472 ( .clk (signal_46981), .D ({signal_5419, signal_3063}), .Q ({signal_4568, signal_4273}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3475 ( .clk (signal_46981), .D ({signal_5421, signal_3065}), .Q ({signal_4571, signal_4272}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3478 ( .clk (signal_46981), .D ({signal_5423, signal_3067}), .Q ({signal_4574, signal_4271}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3481 ( .clk (signal_46981), .D ({signal_5425, signal_3069}), .Q ({signal_4577, signal_4270}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3484 ( .clk (signal_46981), .D ({signal_5427, signal_3071}), .Q ({signal_4580, signal_4269}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3487 ( .clk (signal_46981), .D ({signal_5429, signal_3073}), .Q ({signal_4586, signal_4268}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3490 ( .clk (signal_46981), .D ({signal_5431, signal_3075}), .Q ({signal_4589, signal_4267}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3493 ( .clk (signal_46981), .D ({signal_5433, signal_3077}), .Q ({signal_4592, signal_4266}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3496 ( .clk (signal_46981), .D ({signal_5435, signal_3079}), .Q ({signal_4595, signal_4265}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3499 ( .clk (signal_46981), .D ({signal_5437, signal_3081}), .Q ({signal_4598, signal_4264}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3502 ( .clk (signal_46981), .D ({signal_5439, signal_3083}), .Q ({signal_4601, signal_4263}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3505 ( .clk (signal_46981), .D ({signal_5441, signal_3085}), .Q ({signal_4604, signal_4262}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3508 ( .clk (signal_46981), .D ({signal_5443, signal_3087}), .Q ({signal_4607, signal_4261}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3511 ( .clk (signal_46981), .D ({signal_5445, signal_3089}), .Q ({signal_4610, signal_4260}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3514 ( .clk (signal_46981), .D ({signal_5447, signal_3091}), .Q ({signal_4613, signal_4259}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3517 ( .clk (signal_46981), .D ({signal_5782, signal_3093}), .Q ({signal_4619, signal_4258}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3520 ( .clk (signal_46981), .D ({signal_5784, signal_3095}), .Q ({signal_4622, signal_4257}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3523 ( .clk (signal_46981), .D ({signal_5968, signal_3097}), .Q ({signal_4625, signal_4256}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3526 ( .clk (signal_46981), .D ({signal_5970, signal_3099}), .Q ({signal_4628, signal_4255}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3529 ( .clk (signal_46981), .D ({signal_5874, signal_3101}), .Q ({signal_4631, signal_4254}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3532 ( .clk (signal_46981), .D ({signal_5972, signal_3103}), .Q ({signal_4634, signal_4253}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3535 ( .clk (signal_46981), .D ({signal_5786, signal_3105}), .Q ({signal_4637, signal_4252}) ) ;
    reg_masked #(.low_latency(1), .pipeline(0)) cell_3538 ( .clk (signal_46981), .D ({signal_5876, signal_3107}), .Q ({signal_4640, signal_4251}) ) ;
    DFF_X1 cell_4202 ( .CK (signal_46981), .D (signal_3612), .Q (signal_4388), .QN () ) ;
    DFF_X1 cell_4204 ( .CK (signal_46981), .D (signal_3610), .Q (signal_4387), .QN () ) ;
    DFF_X1 cell_4206 ( .CK (signal_46981), .D (signal_3607), .Q (signal_4386), .QN () ) ;
    DFF_X1 cell_4208 ( .CK (signal_46981), .D (signal_3608), .Q (signal_4385), .QN () ) ;
endmodule
