/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* 16 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 17 register stage(s) in total */

module sbox_HPC2_BDDsylvan_Pipeline_d2 (SI_s0, clk, SI_s1, SI_s2, Fresh, SO_s0, SO_s1, SO_s2);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [1229:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    wire signal_23 ;
    wire signal_24 ;
    wire signal_25 ;
    wire signal_26 ;
    wire signal_27 ;
    wire signal_28 ;
    wire signal_29 ;
    wire signal_30 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;

    /* cells in depth 0 */

    /* cells in depth 1 */
    buf_clk cell_1337 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( signal_3426 ) ) ;
    buf_clk cell_1339 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( signal_3428 ) ) ;
    buf_clk cell_1341 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( signal_3430 ) ) ;
    buf_clk cell_1343 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( signal_3432 ) ) ;
    buf_clk cell_1345 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( signal_3434 ) ) ;
    buf_clk cell_1347 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( signal_3436 ) ) ;
    buf_clk cell_1379 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( signal_3468 ) ) ;
    buf_clk cell_1383 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( signal_3472 ) ) ;
    buf_clk cell_1387 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( signal_3476 ) ) ;
    buf_clk cell_1529 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( signal_3618 ) ) ;
    buf_clk cell_1537 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( signal_3626 ) ) ;
    buf_clk cell_1545 ( .C ( clk ), .D ( SI_s2[4] ), .Q ( signal_3634 ) ) ;
    buf_clk cell_1559 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( signal_3648 ) ) ;
    buf_clk cell_1569 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( signal_3658 ) ) ;
    buf_clk cell_1579 ( .C ( clk ), .D ( SI_s2[5] ), .Q ( signal_3668 ) ) ;
    buf_clk cell_1589 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( signal_3678 ) ) ;
    buf_clk cell_1601 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( signal_3690 ) ) ;
    buf_clk cell_1613 ( .C ( clk ), .D ( SI_s2[6] ), .Q ( signal_3702 ) ) ;
    buf_clk cell_1625 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( signal_3714 ) ) ;
    buf_clk cell_1639 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( signal_3728 ) ) ;
    buf_clk cell_1653 ( .C ( clk ), .D ( SI_s2[7] ), .Q ( signal_3742 ) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_927 ( .s ({SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_1347, signal_1346, signal_942}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_928 ( .s ({SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({signal_1349, signal_1348, signal_943}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_929 ( .s ({SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_1353, signal_1352, signal_944}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_930 ( .s ({SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({signal_1355, signal_1354, signal_945}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_931 ( .s ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_1359, signal_1358, signal_946}) ) ;
    buf_clk cell_1338 ( .C ( clk ), .D ( signal_3426 ), .Q ( signal_3427 ) ) ;
    buf_clk cell_1340 ( .C ( clk ), .D ( signal_3428 ), .Q ( signal_3429 ) ) ;
    buf_clk cell_1342 ( .C ( clk ), .D ( signal_3430 ), .Q ( signal_3431 ) ) ;
    buf_clk cell_1344 ( .C ( clk ), .D ( signal_3432 ), .Q ( signal_3433 ) ) ;
    buf_clk cell_1346 ( .C ( clk ), .D ( signal_3434 ), .Q ( signal_3435 ) ) ;
    buf_clk cell_1348 ( .C ( clk ), .D ( signal_3436 ), .Q ( signal_3437 ) ) ;
    buf_clk cell_1380 ( .C ( clk ), .D ( signal_3468 ), .Q ( signal_3469 ) ) ;
    buf_clk cell_1384 ( .C ( clk ), .D ( signal_3472 ), .Q ( signal_3473 ) ) ;
    buf_clk cell_1388 ( .C ( clk ), .D ( signal_3476 ), .Q ( signal_3477 ) ) ;
    buf_clk cell_1530 ( .C ( clk ), .D ( signal_3618 ), .Q ( signal_3619 ) ) ;
    buf_clk cell_1538 ( .C ( clk ), .D ( signal_3626 ), .Q ( signal_3627 ) ) ;
    buf_clk cell_1546 ( .C ( clk ), .D ( signal_3634 ), .Q ( signal_3635 ) ) ;
    buf_clk cell_1560 ( .C ( clk ), .D ( signal_3648 ), .Q ( signal_3649 ) ) ;
    buf_clk cell_1570 ( .C ( clk ), .D ( signal_3658 ), .Q ( signal_3659 ) ) ;
    buf_clk cell_1580 ( .C ( clk ), .D ( signal_3668 ), .Q ( signal_3669 ) ) ;
    buf_clk cell_1590 ( .C ( clk ), .D ( signal_3678 ), .Q ( signal_3679 ) ) ;
    buf_clk cell_1602 ( .C ( clk ), .D ( signal_3690 ), .Q ( signal_3691 ) ) ;
    buf_clk cell_1614 ( .C ( clk ), .D ( signal_3702 ), .Q ( signal_3703 ) ) ;
    buf_clk cell_1626 ( .C ( clk ), .D ( signal_3714 ), .Q ( signal_3715 ) ) ;
    buf_clk cell_1640 ( .C ( clk ), .D ( signal_3728 ), .Q ( signal_3729 ) ) ;
    buf_clk cell_1654 ( .C ( clk ), .D ( signal_3742 ), .Q ( signal_3743 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_1349 ( .C ( clk ), .D ( signal_3433 ), .Q ( signal_3438 ) ) ;
    buf_clk cell_1351 ( .C ( clk ), .D ( signal_3435 ), .Q ( signal_3440 ) ) ;
    buf_clk cell_1353 ( .C ( clk ), .D ( signal_3437 ), .Q ( signal_3442 ) ) ;
    buf_clk cell_1355 ( .C ( clk ), .D ( signal_943 ), .Q ( signal_3444 ) ) ;
    buf_clk cell_1357 ( .C ( clk ), .D ( signal_1348 ), .Q ( signal_3446 ) ) ;
    buf_clk cell_1359 ( .C ( clk ), .D ( signal_1349 ), .Q ( signal_3448 ) ) ;
    buf_clk cell_1361 ( .C ( clk ), .D ( signal_944 ), .Q ( signal_3450 ) ) ;
    buf_clk cell_1363 ( .C ( clk ), .D ( signal_1352 ), .Q ( signal_3452 ) ) ;
    buf_clk cell_1365 ( .C ( clk ), .D ( signal_1353 ), .Q ( signal_3454 ) ) ;
    buf_clk cell_1367 ( .C ( clk ), .D ( signal_942 ), .Q ( signal_3456 ) ) ;
    buf_clk cell_1369 ( .C ( clk ), .D ( signal_1346 ), .Q ( signal_3458 ) ) ;
    buf_clk cell_1371 ( .C ( clk ), .D ( signal_1347 ), .Q ( signal_3460 ) ) ;
    buf_clk cell_1373 ( .C ( clk ), .D ( signal_945 ), .Q ( signal_3462 ) ) ;
    buf_clk cell_1375 ( .C ( clk ), .D ( signal_1354 ), .Q ( signal_3464 ) ) ;
    buf_clk cell_1377 ( .C ( clk ), .D ( signal_1355 ), .Q ( signal_3466 ) ) ;
    buf_clk cell_1381 ( .C ( clk ), .D ( signal_3469 ), .Q ( signal_3470 ) ) ;
    buf_clk cell_1385 ( .C ( clk ), .D ( signal_3473 ), .Q ( signal_3474 ) ) ;
    buf_clk cell_1389 ( .C ( clk ), .D ( signal_3477 ), .Q ( signal_3478 ) ) ;
    buf_clk cell_1451 ( .C ( clk ), .D ( signal_946 ), .Q ( signal_3540 ) ) ;
    buf_clk cell_1455 ( .C ( clk ), .D ( signal_1358 ), .Q ( signal_3544 ) ) ;
    buf_clk cell_1459 ( .C ( clk ), .D ( signal_1359 ), .Q ( signal_3548 ) ) ;
    buf_clk cell_1531 ( .C ( clk ), .D ( signal_3619 ), .Q ( signal_3620 ) ) ;
    buf_clk cell_1539 ( .C ( clk ), .D ( signal_3627 ), .Q ( signal_3628 ) ) ;
    buf_clk cell_1547 ( .C ( clk ), .D ( signal_3635 ), .Q ( signal_3636 ) ) ;
    buf_clk cell_1561 ( .C ( clk ), .D ( signal_3649 ), .Q ( signal_3650 ) ) ;
    buf_clk cell_1571 ( .C ( clk ), .D ( signal_3659 ), .Q ( signal_3660 ) ) ;
    buf_clk cell_1581 ( .C ( clk ), .D ( signal_3669 ), .Q ( signal_3670 ) ) ;
    buf_clk cell_1591 ( .C ( clk ), .D ( signal_3679 ), .Q ( signal_3680 ) ) ;
    buf_clk cell_1603 ( .C ( clk ), .D ( signal_3691 ), .Q ( signal_3692 ) ) ;
    buf_clk cell_1615 ( .C ( clk ), .D ( signal_3703 ), .Q ( signal_3704 ) ) ;
    buf_clk cell_1627 ( .C ( clk ), .D ( signal_3715 ), .Q ( signal_3716 ) ) ;
    buf_clk cell_1641 ( .C ( clk ), .D ( signal_3729 ), .Q ( signal_3730 ) ) ;
    buf_clk cell_1655 ( .C ( clk ), .D ( signal_3743 ), .Q ( signal_3744 ) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_932 ( .s ({signal_3431, signal_3429, signal_3427}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1347, signal_1346, signal_942}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({signal_1361, signal_1360, signal_947}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_933 ( .s ({signal_3431, signal_3429, signal_3427}), .b ({signal_1347, signal_1346, signal_942}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_1363, signal_1362, signal_948}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_934 ( .s ({signal_3431, signal_3429, signal_3427}), .b ({signal_1349, signal_1348, signal_943}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({signal_1365, signal_1364, signal_949}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_935 ( .s ({signal_3431, signal_3429, signal_3427}), .b ({signal_1347, signal_1346, signal_942}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_1367, signal_1366, signal_950}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_936 ( .s ({signal_3431, signal_3429, signal_3427}), .b ({signal_1347, signal_1346, signal_942}), .a ({signal_1349, signal_1348, signal_943}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({signal_1369, signal_1368, signal_951}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_937 ( .s ({signal_3431, signal_3429, signal_3427}), .b ({signal_1349, signal_1348, signal_943}), .a ({signal_1347, signal_1346, signal_942}), .clk ( clk ), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_1371, signal_1370, signal_952}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_938 ( .s ({signal_3431, signal_3429, signal_3427}), .b ({signal_1349, signal_1348, signal_943}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({signal_1373, signal_1372, signal_953}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_939 ( .s ({signal_3431, signal_3429, signal_3427}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_1347, signal_1346, signal_942}), .clk ( clk ), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_1375, signal_1374, signal_954}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_940 ( .s ({signal_3431, signal_3429, signal_3427}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_1349, signal_1348, signal_943}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({signal_1377, signal_1376, signal_955}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_941 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1355, signal_1354, signal_945}), .clk ( clk ), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_1379, signal_1378, signal_956}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_942 ( .s ({signal_3431, signal_3429, signal_3427}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1349, signal_1348, signal_943}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({signal_1381, signal_1380, signal_957}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_943 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1349, signal_1348, signal_943}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_1383, signal_1382, signal_958}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_944 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1353, signal_1352, signal_944}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({signal_1385, signal_1384, signal_959}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_945 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1353, signal_1352, signal_944}), .a ({signal_1347, signal_1346, signal_942}), .clk ( clk ), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_1387, signal_1386, signal_960}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_946 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1355, signal_1354, signal_945}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({signal_1389, signal_1388, signal_961}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_947 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1355, signal_1354, signal_945}), .a ({signal_1349, signal_1348, signal_943}), .clk ( clk ), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_1391, signal_1390, signal_962}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_948 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1355, signal_1354, signal_945}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({signal_1393, signal_1392, signal_963}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_949 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_1353, signal_1352, signal_944}), .clk ( clk ), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_1395, signal_1394, signal_964}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_950 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1353, signal_1352, signal_944}), .a ({signal_1349, signal_1348, signal_943}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({signal_1397, signal_1396, signal_965}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_951 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_1347, signal_1346, signal_942}), .clk ( clk ), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_1399, signal_1398, signal_966}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_952 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1349, signal_1348, signal_943}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({signal_1401, signal_1400, signal_967}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_953 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1355, signal_1354, signal_945}), .a ({signal_1353, signal_1352, signal_944}), .clk ( clk ), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_1403, signal_1402, signal_968}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_954 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1349, signal_1348, signal_943}), .a ({signal_1355, signal_1354, signal_945}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({signal_1405, signal_1404, signal_969}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_955 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1353, signal_1352, signal_944}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_1407, signal_1406, signal_970}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_956 ( .s ({signal_3437, signal_3435, signal_3433}), .b ({signal_1355, signal_1354, signal_945}), .a ({signal_1347, signal_1346, signal_942}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({signal_1409, signal_1408, signal_971}) ) ;
    buf_clk cell_1350 ( .C ( clk ), .D ( signal_3438 ), .Q ( signal_3439 ) ) ;
    buf_clk cell_1352 ( .C ( clk ), .D ( signal_3440 ), .Q ( signal_3441 ) ) ;
    buf_clk cell_1354 ( .C ( clk ), .D ( signal_3442 ), .Q ( signal_3443 ) ) ;
    buf_clk cell_1356 ( .C ( clk ), .D ( signal_3444 ), .Q ( signal_3445 ) ) ;
    buf_clk cell_1358 ( .C ( clk ), .D ( signal_3446 ), .Q ( signal_3447 ) ) ;
    buf_clk cell_1360 ( .C ( clk ), .D ( signal_3448 ), .Q ( signal_3449 ) ) ;
    buf_clk cell_1362 ( .C ( clk ), .D ( signal_3450 ), .Q ( signal_3451 ) ) ;
    buf_clk cell_1364 ( .C ( clk ), .D ( signal_3452 ), .Q ( signal_3453 ) ) ;
    buf_clk cell_1366 ( .C ( clk ), .D ( signal_3454 ), .Q ( signal_3455 ) ) ;
    buf_clk cell_1368 ( .C ( clk ), .D ( signal_3456 ), .Q ( signal_3457 ) ) ;
    buf_clk cell_1370 ( .C ( clk ), .D ( signal_3458 ), .Q ( signal_3459 ) ) ;
    buf_clk cell_1372 ( .C ( clk ), .D ( signal_3460 ), .Q ( signal_3461 ) ) ;
    buf_clk cell_1374 ( .C ( clk ), .D ( signal_3462 ), .Q ( signal_3463 ) ) ;
    buf_clk cell_1376 ( .C ( clk ), .D ( signal_3464 ), .Q ( signal_3465 ) ) ;
    buf_clk cell_1378 ( .C ( clk ), .D ( signal_3466 ), .Q ( signal_3467 ) ) ;
    buf_clk cell_1382 ( .C ( clk ), .D ( signal_3470 ), .Q ( signal_3471 ) ) ;
    buf_clk cell_1386 ( .C ( clk ), .D ( signal_3474 ), .Q ( signal_3475 ) ) ;
    buf_clk cell_1390 ( .C ( clk ), .D ( signal_3478 ), .Q ( signal_3479 ) ) ;
    buf_clk cell_1452 ( .C ( clk ), .D ( signal_3540 ), .Q ( signal_3541 ) ) ;
    buf_clk cell_1456 ( .C ( clk ), .D ( signal_3544 ), .Q ( signal_3545 ) ) ;
    buf_clk cell_1460 ( .C ( clk ), .D ( signal_3548 ), .Q ( signal_3549 ) ) ;
    buf_clk cell_1532 ( .C ( clk ), .D ( signal_3620 ), .Q ( signal_3621 ) ) ;
    buf_clk cell_1540 ( .C ( clk ), .D ( signal_3628 ), .Q ( signal_3629 ) ) ;
    buf_clk cell_1548 ( .C ( clk ), .D ( signal_3636 ), .Q ( signal_3637 ) ) ;
    buf_clk cell_1562 ( .C ( clk ), .D ( signal_3650 ), .Q ( signal_3651 ) ) ;
    buf_clk cell_1572 ( .C ( clk ), .D ( signal_3660 ), .Q ( signal_3661 ) ) ;
    buf_clk cell_1582 ( .C ( clk ), .D ( signal_3670 ), .Q ( signal_3671 ) ) ;
    buf_clk cell_1592 ( .C ( clk ), .D ( signal_3680 ), .Q ( signal_3681 ) ) ;
    buf_clk cell_1604 ( .C ( clk ), .D ( signal_3692 ), .Q ( signal_3693 ) ) ;
    buf_clk cell_1616 ( .C ( clk ), .D ( signal_3704 ), .Q ( signal_3705 ) ) ;
    buf_clk cell_1628 ( .C ( clk ), .D ( signal_3716 ), .Q ( signal_3717 ) ) ;
    buf_clk cell_1642 ( .C ( clk ), .D ( signal_3730 ), .Q ( signal_3731 ) ) ;
    buf_clk cell_1656 ( .C ( clk ), .D ( signal_3744 ), .Q ( signal_3745 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_1391 ( .C ( clk ), .D ( signal_3471 ), .Q ( signal_3480 ) ) ;
    buf_clk cell_1393 ( .C ( clk ), .D ( signal_3475 ), .Q ( signal_3482 ) ) ;
    buf_clk cell_1395 ( .C ( clk ), .D ( signal_3479 ), .Q ( signal_3484 ) ) ;
    buf_clk cell_1397 ( .C ( clk ), .D ( signal_956 ), .Q ( signal_3486 ) ) ;
    buf_clk cell_1399 ( .C ( clk ), .D ( signal_1378 ), .Q ( signal_3488 ) ) ;
    buf_clk cell_1401 ( .C ( clk ), .D ( signal_1379 ), .Q ( signal_3490 ) ) ;
    buf_clk cell_1403 ( .C ( clk ), .D ( signal_958 ), .Q ( signal_3492 ) ) ;
    buf_clk cell_1405 ( .C ( clk ), .D ( signal_1382 ), .Q ( signal_3494 ) ) ;
    buf_clk cell_1407 ( .C ( clk ), .D ( signal_1383 ), .Q ( signal_3496 ) ) ;
    buf_clk cell_1409 ( .C ( clk ), .D ( signal_959 ), .Q ( signal_3498 ) ) ;
    buf_clk cell_1411 ( .C ( clk ), .D ( signal_1384 ), .Q ( signal_3500 ) ) ;
    buf_clk cell_1413 ( .C ( clk ), .D ( signal_1385 ), .Q ( signal_3502 ) ) ;
    buf_clk cell_1415 ( .C ( clk ), .D ( signal_960 ), .Q ( signal_3504 ) ) ;
    buf_clk cell_1417 ( .C ( clk ), .D ( signal_1386 ), .Q ( signal_3506 ) ) ;
    buf_clk cell_1419 ( .C ( clk ), .D ( signal_1387 ), .Q ( signal_3508 ) ) ;
    buf_clk cell_1421 ( .C ( clk ), .D ( signal_961 ), .Q ( signal_3510 ) ) ;
    buf_clk cell_1423 ( .C ( clk ), .D ( signal_1388 ), .Q ( signal_3512 ) ) ;
    buf_clk cell_1425 ( .C ( clk ), .D ( signal_1389 ), .Q ( signal_3514 ) ) ;
    buf_clk cell_1427 ( .C ( clk ), .D ( signal_962 ), .Q ( signal_3516 ) ) ;
    buf_clk cell_1429 ( .C ( clk ), .D ( signal_1390 ), .Q ( signal_3518 ) ) ;
    buf_clk cell_1431 ( .C ( clk ), .D ( signal_1391 ), .Q ( signal_3520 ) ) ;
    buf_clk cell_1433 ( .C ( clk ), .D ( signal_963 ), .Q ( signal_3522 ) ) ;
    buf_clk cell_1435 ( .C ( clk ), .D ( signal_1392 ), .Q ( signal_3524 ) ) ;
    buf_clk cell_1437 ( .C ( clk ), .D ( signal_1393 ), .Q ( signal_3526 ) ) ;
    buf_clk cell_1439 ( .C ( clk ), .D ( signal_964 ), .Q ( signal_3528 ) ) ;
    buf_clk cell_1441 ( .C ( clk ), .D ( signal_1394 ), .Q ( signal_3530 ) ) ;
    buf_clk cell_1443 ( .C ( clk ), .D ( signal_1395 ), .Q ( signal_3532 ) ) ;
    buf_clk cell_1445 ( .C ( clk ), .D ( signal_965 ), .Q ( signal_3534 ) ) ;
    buf_clk cell_1447 ( .C ( clk ), .D ( signal_1396 ), .Q ( signal_3536 ) ) ;
    buf_clk cell_1449 ( .C ( clk ), .D ( signal_1397 ), .Q ( signal_3538 ) ) ;
    buf_clk cell_1453 ( .C ( clk ), .D ( signal_3541 ), .Q ( signal_3542 ) ) ;
    buf_clk cell_1457 ( .C ( clk ), .D ( signal_3545 ), .Q ( signal_3546 ) ) ;
    buf_clk cell_1461 ( .C ( clk ), .D ( signal_3549 ), .Q ( signal_3550 ) ) ;
    buf_clk cell_1463 ( .C ( clk ), .D ( signal_954 ), .Q ( signal_3552 ) ) ;
    buf_clk cell_1465 ( .C ( clk ), .D ( signal_1374 ), .Q ( signal_3554 ) ) ;
    buf_clk cell_1467 ( .C ( clk ), .D ( signal_1375 ), .Q ( signal_3556 ) ) ;
    buf_clk cell_1469 ( .C ( clk ), .D ( signal_3463 ), .Q ( signal_3558 ) ) ;
    buf_clk cell_1471 ( .C ( clk ), .D ( signal_3465 ), .Q ( signal_3560 ) ) ;
    buf_clk cell_1473 ( .C ( clk ), .D ( signal_3467 ), .Q ( signal_3562 ) ) ;
    buf_clk cell_1475 ( .C ( clk ), .D ( signal_3445 ), .Q ( signal_3564 ) ) ;
    buf_clk cell_1477 ( .C ( clk ), .D ( signal_3447 ), .Q ( signal_3566 ) ) ;
    buf_clk cell_1479 ( .C ( clk ), .D ( signal_3449 ), .Q ( signal_3568 ) ) ;
    buf_clk cell_1481 ( .C ( clk ), .D ( signal_966 ), .Q ( signal_3570 ) ) ;
    buf_clk cell_1483 ( .C ( clk ), .D ( signal_1398 ), .Q ( signal_3572 ) ) ;
    buf_clk cell_1485 ( .C ( clk ), .D ( signal_1399 ), .Q ( signal_3574 ) ) ;
    buf_clk cell_1487 ( .C ( clk ), .D ( signal_950 ), .Q ( signal_3576 ) ) ;
    buf_clk cell_1489 ( .C ( clk ), .D ( signal_1366 ), .Q ( signal_3578 ) ) ;
    buf_clk cell_1491 ( .C ( clk ), .D ( signal_1367 ), .Q ( signal_3580 ) ) ;
    buf_clk cell_1493 ( .C ( clk ), .D ( signal_3451 ), .Q ( signal_3582 ) ) ;
    buf_clk cell_1495 ( .C ( clk ), .D ( signal_3453 ), .Q ( signal_3584 ) ) ;
    buf_clk cell_1497 ( .C ( clk ), .D ( signal_3455 ), .Q ( signal_3586 ) ) ;
    buf_clk cell_1499 ( .C ( clk ), .D ( signal_967 ), .Q ( signal_3588 ) ) ;
    buf_clk cell_1501 ( .C ( clk ), .D ( signal_1400 ), .Q ( signal_3590 ) ) ;
    buf_clk cell_1503 ( .C ( clk ), .D ( signal_1401 ), .Q ( signal_3592 ) ) ;
    buf_clk cell_1505 ( .C ( clk ), .D ( signal_968 ), .Q ( signal_3594 ) ) ;
    buf_clk cell_1507 ( .C ( clk ), .D ( signal_1402 ), .Q ( signal_3596 ) ) ;
    buf_clk cell_1509 ( .C ( clk ), .D ( signal_1403 ), .Q ( signal_3598 ) ) ;
    buf_clk cell_1511 ( .C ( clk ), .D ( signal_947 ), .Q ( signal_3600 ) ) ;
    buf_clk cell_1513 ( .C ( clk ), .D ( signal_1360 ), .Q ( signal_3602 ) ) ;
    buf_clk cell_1515 ( .C ( clk ), .D ( signal_1361 ), .Q ( signal_3604 ) ) ;
    buf_clk cell_1517 ( .C ( clk ), .D ( signal_969 ), .Q ( signal_3606 ) ) ;
    buf_clk cell_1519 ( .C ( clk ), .D ( signal_1404 ), .Q ( signal_3608 ) ) ;
    buf_clk cell_1521 ( .C ( clk ), .D ( signal_1405 ), .Q ( signal_3610 ) ) ;
    buf_clk cell_1523 ( .C ( clk ), .D ( signal_970 ), .Q ( signal_3612 ) ) ;
    buf_clk cell_1525 ( .C ( clk ), .D ( signal_1406 ), .Q ( signal_3614 ) ) ;
    buf_clk cell_1527 ( .C ( clk ), .D ( signal_1407 ), .Q ( signal_3616 ) ) ;
    buf_clk cell_1533 ( .C ( clk ), .D ( signal_3621 ), .Q ( signal_3622 ) ) ;
    buf_clk cell_1541 ( .C ( clk ), .D ( signal_3629 ), .Q ( signal_3630 ) ) ;
    buf_clk cell_1549 ( .C ( clk ), .D ( signal_3637 ), .Q ( signal_3638 ) ) ;
    buf_clk cell_1563 ( .C ( clk ), .D ( signal_3651 ), .Q ( signal_3652 ) ) ;
    buf_clk cell_1573 ( .C ( clk ), .D ( signal_3661 ), .Q ( signal_3662 ) ) ;
    buf_clk cell_1583 ( .C ( clk ), .D ( signal_3671 ), .Q ( signal_3672 ) ) ;
    buf_clk cell_1593 ( .C ( clk ), .D ( signal_3681 ), .Q ( signal_3682 ) ) ;
    buf_clk cell_1605 ( .C ( clk ), .D ( signal_3693 ), .Q ( signal_3694 ) ) ;
    buf_clk cell_1617 ( .C ( clk ), .D ( signal_3705 ), .Q ( signal_3706 ) ) ;
    buf_clk cell_1629 ( .C ( clk ), .D ( signal_3717 ), .Q ( signal_3718 ) ) ;
    buf_clk cell_1643 ( .C ( clk ), .D ( signal_3731 ), .Q ( signal_3732 ) ) ;
    buf_clk cell_1657 ( .C ( clk ), .D ( signal_3745 ), .Q ( signal_3746 ) ) ;

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_957 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_1361, signal_1360, signal_947}), .clk ( clk ), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_1411, signal_1410, signal_972}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_958 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1365, signal_1364, signal_949}), .a ({signal_1363, signal_1362, signal_948}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({signal_1413, signal_1412, signal_973}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_959 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1367, signal_1366, signal_950}), .a ({signal_3449, signal_3447, signal_3445}), .clk ( clk ), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_1415, signal_1414, signal_974}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_960 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1369, signal_1368, signal_951}), .a ({signal_3455, signal_3453, signal_3451}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({signal_1417, signal_1416, signal_975}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_961 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_1419, signal_1418, signal_976}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_962 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({signal_1373, signal_1372, signal_953}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({signal_1421, signal_1420, signal_977}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_963 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3449, signal_3447, signal_3445}), .a ({signal_1375, signal_1374, signal_954}), .clk ( clk ), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_1423, signal_1422, signal_978}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_964 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({signal_1425, signal_1424, signal_979}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_965 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1363, signal_1362, signal_948}), .clk ( clk ), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_1427, signal_1426, signal_980}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_966 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1367, signal_1366, signal_950}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({signal_1429, signal_1428, signal_981}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_967 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1373, signal_1372, signal_953}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_1431, signal_1430, signal_982}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_968 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1371, signal_1370, signal_952}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({signal_1433, signal_1432, signal_983}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_969 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3449, signal_3447, signal_3445}), .a ({signal_1365, signal_1364, signal_949}), .clk ( clk ), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_1435, signal_1434, signal_984}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_970 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3461, signal_3459, signal_3457}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({signal_1437, signal_1436, signal_985}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_971 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_1439, signal_1438, signal_986}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_972 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1377, signal_1376, signal_955}), .a ({signal_3449, signal_3447, signal_3445}), .clk ( clk ), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({signal_1441, signal_1440, signal_987}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_973 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1377, signal_1376, signal_955}), .a ({signal_1361, signal_1360, signal_947}), .clk ( clk ), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_1443, signal_1442, signal_988}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_974 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3449, signal_3447, signal_3445}), .a ({signal_1381, signal_1380, signal_957}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({signal_1445, signal_1444, signal_989}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_975 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1377, signal_1376, signal_955}), .a ({signal_3467, signal_3465, signal_3463}), .clk ( clk ), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_1447, signal_1446, signal_990}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_976 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3455, signal_3453, signal_3451}), .a ({signal_1363, signal_1362, signal_948}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({signal_1449, signal_1448, signal_991}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_977 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1363, signal_1362, signal_948}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_1451, signal_1450, signal_992}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_978 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1365, signal_1364, signal_949}), .a ({signal_1361, signal_1360, signal_947}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({signal_1453, signal_1452, signal_993}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_979 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1365, signal_1364, signal_949}), .a ({signal_1367, signal_1366, signal_950}), .clk ( clk ), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_1455, signal_1454, signal_994}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_980 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1375, signal_1374, signal_954}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({signal_1457, signal_1456, signal_995}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_981 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1369, signal_1368, signal_951}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_1459, signal_1458, signal_996}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_982 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3467, signal_3465, signal_3463}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({signal_1461, signal_1460, signal_997}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_983 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1365, signal_1364, signal_949}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_1463, signal_1462, signal_998}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_984 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1367, signal_1366, signal_950}), .a ({signal_1365, signal_1364, signal_949}), .clk ( clk ), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({signal_1465, signal_1464, signal_999}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_985 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({signal_3467, signal_3465, signal_3463}), .clk ( clk ), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_1467, signal_1466, signal_1000}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_986 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1375, signal_1374, signal_954}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({signal_1469, signal_1468, signal_1001}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_987 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1375, signal_1374, signal_954}), .a ({signal_1369, signal_1368, signal_951}), .clk ( clk ), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_1471, signal_1470, signal_1002}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_988 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1361, signal_1360, signal_947}), .clk ( clk ), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({signal_1473, signal_1472, signal_1003}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_989 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({signal_1369, signal_1368, signal_951}), .clk ( clk ), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_1475, signal_1474, signal_1004}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_990 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({signal_1367, signal_1366, signal_950}), .clk ( clk ), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({signal_1477, signal_1476, signal_1005}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_991 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1369, signal_1368, signal_951}), .a ({signal_3449, signal_3447, signal_3445}), .clk ( clk ), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_1479, signal_1478, signal_1006}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_992 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3449, signal_3447, signal_3445}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({signal_1481, signal_1480, signal_1007}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_993 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3461, signal_3459, signal_3457}), .a ({signal_1361, signal_1360, signal_947}), .clk ( clk ), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_1483, signal_1482, signal_1008}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_994 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1377, signal_1376, signal_955}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({signal_1485, signal_1484, signal_1009}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_995 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1365, signal_1364, signal_949}), .a ({signal_1373, signal_1372, signal_953}), .clk ( clk ), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({signal_1487, signal_1486, signal_1010}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_996 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({signal_3455, signal_3453, signal_3451}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({signal_1489, signal_1488, signal_1011}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_997 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1371, signal_1370, signal_952}), .a ({signal_1381, signal_1380, signal_957}), .clk ( clk ), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_1491, signal_1490, signal_1012}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_998 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({signal_1493, signal_1492, signal_1013}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_999 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1371, signal_1370, signal_952}), .a ({signal_1365, signal_1364, signal_949}), .clk ( clk ), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({signal_1495, signal_1494, signal_1014}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1000 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3449, signal_3447, signal_3445}), .a ({signal_1363, signal_1362, signal_948}), .clk ( clk ), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({signal_1497, signal_1496, signal_1015}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1001 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3467, signal_3465, signal_3463}), .a ({signal_1361, signal_1360, signal_947}), .clk ( clk ), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({signal_1499, signal_1498, signal_1016}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1002 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1365, signal_1364, signal_949}), .a ({signal_3461, signal_3459, signal_3457}), .clk ( clk ), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({signal_1501, signal_1500, signal_1017}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1003 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1363, signal_1362, signal_948}), .a ({signal_1381, signal_1380, signal_957}), .clk ( clk ), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({signal_1503, signal_1502, signal_1018}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1004 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1377, signal_1376, signal_955}), .a ({signal_1375, signal_1374, signal_954}), .clk ( clk ), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({signal_1505, signal_1504, signal_1019}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1005 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1365, signal_1364, signal_949}), .a ({signal_3449, signal_3447, signal_3445}), .clk ( clk ), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({signal_1507, signal_1506, signal_1020}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1006 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1367, signal_1366, signal_950}), .a ({signal_1375, signal_1374, signal_954}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({signal_1509, signal_1508, signal_1021}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1007 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1371, signal_1370, signal_952}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_1511, signal_1510, signal_1022}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1008 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1371, signal_1370, signal_952}), .a ({signal_1367, signal_1366, signal_950}), .clk ( clk ), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({signal_1513, signal_1512, signal_1023}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1009 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1365, signal_1364, signal_949}), .a ({signal_3467, signal_3465, signal_3463}), .clk ( clk ), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({signal_1515, signal_1514, signal_1024}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1010 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1375, signal_1374, signal_954}), .a ({signal_3461, signal_3459, signal_3457}), .clk ( clk ), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({signal_1517, signal_1516, signal_1025}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1011 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({signal_1519, signal_1518, signal_1026}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1012 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1365, signal_1364, signal_949}), .clk ( clk ), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({signal_1521, signal_1520, signal_1027}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1013 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1377, signal_1376, signal_955}), .a ({signal_3455, signal_3453, signal_3451}), .clk ( clk ), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({signal_1523, signal_1522, signal_1028}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1014 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1377, signal_1376, signal_955}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({signal_1525, signal_1524, signal_1029}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1015 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3455, signal_3453, signal_3451}), .a ({signal_1373, signal_1372, signal_953}), .clk ( clk ), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({signal_1527, signal_1526, signal_1030}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1016 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({signal_3449, signal_3447, signal_3445}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({signal_1529, signal_1528, signal_1031}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1017 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1369, signal_1368, signal_951}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_1531, signal_1530, signal_1032}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1018 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1373, signal_1372, signal_953}), .a ({signal_3449, signal_3447, signal_3445}), .clk ( clk ), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({signal_1533, signal_1532, signal_1033}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1019 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({signal_3449, signal_3447, signal_3445}), .clk ( clk ), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({signal_1535, signal_1534, signal_1034}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1020 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({signal_1373, signal_1372, signal_953}), .clk ( clk ), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({signal_1537, signal_1536, signal_1035}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1021 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({signal_3467, signal_3465, signal_3463}), .clk ( clk ), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({signal_1539, signal_1538, signal_1036}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1022 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1363, signal_1362, signal_948}), .a ({signal_3449, signal_3447, signal_3445}), .clk ( clk ), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({signal_1541, signal_1540, signal_1037}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1023 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3455, signal_3453, signal_3451}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({signal_1543, signal_1542, signal_1038}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1024 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1375, signal_1374, signal_954}), .a ({signal_1381, signal_1380, signal_957}), .clk ( clk ), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({signal_1545, signal_1544, signal_1039}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1025 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({signal_1361, signal_1360, signal_947}), .clk ( clk ), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({signal_1547, signal_1546, signal_1040}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1026 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1371, signal_1370, signal_952}), .a ({signal_3467, signal_3465, signal_3463}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({signal_1549, signal_1548, signal_1041}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1027 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1367, signal_1366, signal_950}), .a ({signal_1369, signal_1368, signal_951}), .clk ( clk ), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_1551, signal_1550, signal_1042}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1028 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1377, signal_1376, signal_955}), .a ({signal_1367, signal_1366, signal_950}), .clk ( clk ), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({signal_1553, signal_1552, signal_1043}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1029 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1371, signal_1370, signal_952}), .a ({signal_1375, signal_1374, signal_954}), .clk ( clk ), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({signal_1555, signal_1554, signal_1044}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1030 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1373, signal_1372, signal_953}), .a ({signal_1369, signal_1368, signal_951}), .clk ( clk ), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({signal_1557, signal_1556, signal_1045}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1031 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1377, signal_1376, signal_955}), .a ({signal_1363, signal_1362, signal_948}), .clk ( clk ), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({signal_1559, signal_1558, signal_1046}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1032 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1369, signal_1368, signal_951}), .a ({signal_1365, signal_1364, signal_949}), .clk ( clk ), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({signal_1561, signal_1560, signal_1047}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1033 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3449, signal_3447, signal_3445}), .a ({signal_1367, signal_1366, signal_950}), .clk ( clk ), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({signal_1563, signal_1562, signal_1048}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1034 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({signal_1381, signal_1380, signal_957}), .clk ( clk ), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({signal_1565, signal_1564, signal_1049}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1035 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3467, signal_3465, signal_3463}), .a ({signal_1369, signal_1368, signal_951}), .clk ( clk ), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({signal_1567, signal_1566, signal_1050}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1036 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1371, signal_1370, signal_952}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({signal_1569, signal_1568, signal_1051}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1037 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3461, signal_3459, signal_3457}), .a ({signal_1373, signal_1372, signal_953}), .clk ( clk ), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_1571, signal_1570, signal_1052}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1038 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1373, signal_1372, signal_953}), .a ({signal_3461, signal_3459, signal_3457}), .clk ( clk ), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({signal_1573, signal_1572, signal_1053}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1039 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1369, signal_1368, signal_951}), .clk ( clk ), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({signal_1575, signal_1574, signal_1054}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1040 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1373, signal_1372, signal_953}), .clk ( clk ), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({signal_1577, signal_1576, signal_1055}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1041 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1369, signal_1368, signal_951}), .a ({signal_1363, signal_1362, signal_948}), .clk ( clk ), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({signal_1579, signal_1578, signal_1056}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1042 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1367, signal_1366, signal_950}), .a ({signal_3455, signal_3453, signal_3451}), .clk ( clk ), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({signal_1581, signal_1580, signal_1057}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1043 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({signal_3461, signal_3459, signal_3457}), .clk ( clk ), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({signal_1583, signal_1582, signal_1058}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1044 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1373, signal_1372, signal_953}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({signal_1585, signal_1584, signal_1059}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1045 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1375, signal_1374, signal_954}), .a ({signal_1361, signal_1360, signal_947}), .clk ( clk ), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({signal_1587, signal_1586, signal_1060}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1046 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1371, signal_1370, signal_952}), .a ({signal_1373, signal_1372, signal_953}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({signal_1589, signal_1588, signal_1061}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1047 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3467, signal_3465, signal_3463}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_1591, signal_1590, signal_1062}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1048 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3467, signal_3465, signal_3463}), .a ({signal_1365, signal_1364, signal_949}), .clk ( clk ), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({signal_1593, signal_1592, signal_1063}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1049 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1375, signal_1374, signal_954}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({signal_1595, signal_1594, signal_1064}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1050 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1363, signal_1362, signal_948}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({signal_1597, signal_1596, signal_1065}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1051 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1369, signal_1368, signal_951}), .a ({signal_1361, signal_1360, signal_947}), .clk ( clk ), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({signal_1599, signal_1598, signal_1066}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1052 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3455, signal_3453, signal_3451}), .a ({signal_1365, signal_1364, signal_949}), .clk ( clk ), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({signal_1601, signal_1600, signal_1067}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1053 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1373, signal_1372, signal_953}), .a ({signal_3467, signal_3465, signal_3463}), .clk ( clk ), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({signal_1603, signal_1602, signal_1068}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1054 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({signal_1605, signal_1604, signal_1069}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1055 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1369, signal_1368, signal_951}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({signal_1607, signal_1606, signal_1070}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1056 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({signal_1609, signal_1608, signal_1071}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1057 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({signal_3461, signal_3459, signal_3457}), .clk ( clk ), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_1611, signal_1610, signal_1072}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1058 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1367, signal_1366, signal_950}), .a ({signal_1381, signal_1380, signal_957}), .clk ( clk ), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({signal_1613, signal_1612, signal_1073}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1059 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1363, signal_1362, signal_948}), .a ({signal_3455, signal_3453, signal_3451}), .clk ( clk ), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({signal_1615, signal_1614, signal_1074}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1060 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1365, signal_1364, signal_949}), .a ({signal_1369, signal_1368, signal_951}), .clk ( clk ), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({signal_1617, signal_1616, signal_1075}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1061 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({signal_1619, signal_1618, signal_1076}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1062 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1377, signal_1376, signal_955}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({signal_1621, signal_1620, signal_1077}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1063 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1367, signal_1366, signal_950}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({signal_1623, signal_1622, signal_1078}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1064 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({signal_1375, signal_1374, signal_954}), .clk ( clk ), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({signal_1625, signal_1624, signal_1079}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1065 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({signal_1627, signal_1626, signal_1080}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1066 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1367, signal_1366, signal_950}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({signal_1629, signal_1628, signal_1081}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1067 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1381, signal_1380, signal_957}), .a ({signal_1369, signal_1368, signal_951}), .clk ( clk ), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_1631, signal_1630, signal_1082}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1068 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_1375, signal_1374, signal_954}), .clk ( clk ), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({signal_1633, signal_1632, signal_1083}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1069 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1363, signal_1362, signal_948}), .a ({signal_1373, signal_1372, signal_953}), .clk ( clk ), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({signal_1635, signal_1634, signal_1084}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1070 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1369, signal_1368, signal_951}), .a ({signal_3461, signal_3459, signal_3457}), .clk ( clk ), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({signal_1637, signal_1636, signal_1085}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1071 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1375, signal_1374, signal_954}), .a ({signal_1363, signal_1362, signal_948}), .clk ( clk ), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({signal_1639, signal_1638, signal_1086}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1072 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1373, signal_1372, signal_953}), .a ({signal_1381, signal_1380, signal_957}), .clk ( clk ), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({signal_1641, signal_1640, signal_1087}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1073 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1363, signal_1362, signal_948}), .a ({signal_1369, signal_1368, signal_951}), .clk ( clk ), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({signal_1643, signal_1642, signal_1088}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1074 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3455, signal_3453, signal_3451}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({signal_1645, signal_1644, signal_1089}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1075 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1361, signal_1360, signal_947}), .a ({signal_1365, signal_1364, signal_949}), .clk ( clk ), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({signal_1647, signal_1646, signal_1090}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1076 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3461, signal_3459, signal_3457}), .a ({signal_1381, signal_1380, signal_957}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({signal_1649, signal_1648, signal_1091}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1077 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_1371, signal_1370, signal_952}), .clk ( clk ), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_1651, signal_1650, signal_1092}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1078 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1367, signal_1366, signal_950}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({signal_1653, signal_1652, signal_1093}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1079 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1375, signal_1374, signal_954}), .a ({signal_3455, signal_3453, signal_3451}), .clk ( clk ), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({signal_1655, signal_1654, signal_1094}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1080 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1375, signal_1374, signal_954}), .a ({signal_1365, signal_1364, signal_949}), .clk ( clk ), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({signal_1657, signal_1656, signal_1095}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1081 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1363, signal_1362, signal_948}), .a ({signal_1365, signal_1364, signal_949}), .clk ( clk ), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({signal_1659, signal_1658, signal_1096}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1082 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1363, signal_1362, signal_948}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({signal_1661, signal_1660, signal_1097}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1083 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1371, signal_1370, signal_952}), .a ({signal_1369, signal_1368, signal_951}), .clk ( clk ), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({signal_1663, signal_1662, signal_1098}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1084 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1369, signal_1368, signal_951}), .a ({signal_1373, signal_1372, signal_953}), .clk ( clk ), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({signal_1665, signal_1664, signal_1099}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1085 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_3449, signal_3447, signal_3445}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({signal_1667, signal_1666, signal_1100}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1086 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_1381, signal_1380, signal_957}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({signal_1669, signal_1668, signal_1101}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1087 ( .s ({signal_3479, signal_3475, signal_3471}), .b ({signal_3449, signal_3447, signal_3445}), .a ({signal_1409, signal_1408, signal_971}), .clk ( clk ), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_1673, signal_1672, signal_1102}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1088 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({signal_1375, signal_1374, signal_954}), .a ({signal_3467, signal_3465, signal_3463}), .clk ( clk ), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({signal_1675, signal_1674, signal_1103}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1089 ( .s ({signal_3443, signal_3441, signal_3439}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_1377, signal_1376, signal_955}), .clk ( clk ), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({signal_1677, signal_1676, signal_1104}) ) ;
    buf_clk cell_1392 ( .C ( clk ), .D ( signal_3480 ), .Q ( signal_3481 ) ) ;
    buf_clk cell_1394 ( .C ( clk ), .D ( signal_3482 ), .Q ( signal_3483 ) ) ;
    buf_clk cell_1396 ( .C ( clk ), .D ( signal_3484 ), .Q ( signal_3485 ) ) ;
    buf_clk cell_1398 ( .C ( clk ), .D ( signal_3486 ), .Q ( signal_3487 ) ) ;
    buf_clk cell_1400 ( .C ( clk ), .D ( signal_3488 ), .Q ( signal_3489 ) ) ;
    buf_clk cell_1402 ( .C ( clk ), .D ( signal_3490 ), .Q ( signal_3491 ) ) ;
    buf_clk cell_1404 ( .C ( clk ), .D ( signal_3492 ), .Q ( signal_3493 ) ) ;
    buf_clk cell_1406 ( .C ( clk ), .D ( signal_3494 ), .Q ( signal_3495 ) ) ;
    buf_clk cell_1408 ( .C ( clk ), .D ( signal_3496 ), .Q ( signal_3497 ) ) ;
    buf_clk cell_1410 ( .C ( clk ), .D ( signal_3498 ), .Q ( signal_3499 ) ) ;
    buf_clk cell_1412 ( .C ( clk ), .D ( signal_3500 ), .Q ( signal_3501 ) ) ;
    buf_clk cell_1414 ( .C ( clk ), .D ( signal_3502 ), .Q ( signal_3503 ) ) ;
    buf_clk cell_1416 ( .C ( clk ), .D ( signal_3504 ), .Q ( signal_3505 ) ) ;
    buf_clk cell_1418 ( .C ( clk ), .D ( signal_3506 ), .Q ( signal_3507 ) ) ;
    buf_clk cell_1420 ( .C ( clk ), .D ( signal_3508 ), .Q ( signal_3509 ) ) ;
    buf_clk cell_1422 ( .C ( clk ), .D ( signal_3510 ), .Q ( signal_3511 ) ) ;
    buf_clk cell_1424 ( .C ( clk ), .D ( signal_3512 ), .Q ( signal_3513 ) ) ;
    buf_clk cell_1426 ( .C ( clk ), .D ( signal_3514 ), .Q ( signal_3515 ) ) ;
    buf_clk cell_1428 ( .C ( clk ), .D ( signal_3516 ), .Q ( signal_3517 ) ) ;
    buf_clk cell_1430 ( .C ( clk ), .D ( signal_3518 ), .Q ( signal_3519 ) ) ;
    buf_clk cell_1432 ( .C ( clk ), .D ( signal_3520 ), .Q ( signal_3521 ) ) ;
    buf_clk cell_1434 ( .C ( clk ), .D ( signal_3522 ), .Q ( signal_3523 ) ) ;
    buf_clk cell_1436 ( .C ( clk ), .D ( signal_3524 ), .Q ( signal_3525 ) ) ;
    buf_clk cell_1438 ( .C ( clk ), .D ( signal_3526 ), .Q ( signal_3527 ) ) ;
    buf_clk cell_1440 ( .C ( clk ), .D ( signal_3528 ), .Q ( signal_3529 ) ) ;
    buf_clk cell_1442 ( .C ( clk ), .D ( signal_3530 ), .Q ( signal_3531 ) ) ;
    buf_clk cell_1444 ( .C ( clk ), .D ( signal_3532 ), .Q ( signal_3533 ) ) ;
    buf_clk cell_1446 ( .C ( clk ), .D ( signal_3534 ), .Q ( signal_3535 ) ) ;
    buf_clk cell_1448 ( .C ( clk ), .D ( signal_3536 ), .Q ( signal_3537 ) ) ;
    buf_clk cell_1450 ( .C ( clk ), .D ( signal_3538 ), .Q ( signal_3539 ) ) ;
    buf_clk cell_1454 ( .C ( clk ), .D ( signal_3542 ), .Q ( signal_3543 ) ) ;
    buf_clk cell_1458 ( .C ( clk ), .D ( signal_3546 ), .Q ( signal_3547 ) ) ;
    buf_clk cell_1462 ( .C ( clk ), .D ( signal_3550 ), .Q ( signal_3551 ) ) ;
    buf_clk cell_1464 ( .C ( clk ), .D ( signal_3552 ), .Q ( signal_3553 ) ) ;
    buf_clk cell_1466 ( .C ( clk ), .D ( signal_3554 ), .Q ( signal_3555 ) ) ;
    buf_clk cell_1468 ( .C ( clk ), .D ( signal_3556 ), .Q ( signal_3557 ) ) ;
    buf_clk cell_1470 ( .C ( clk ), .D ( signal_3558 ), .Q ( signal_3559 ) ) ;
    buf_clk cell_1472 ( .C ( clk ), .D ( signal_3560 ), .Q ( signal_3561 ) ) ;
    buf_clk cell_1474 ( .C ( clk ), .D ( signal_3562 ), .Q ( signal_3563 ) ) ;
    buf_clk cell_1476 ( .C ( clk ), .D ( signal_3564 ), .Q ( signal_3565 ) ) ;
    buf_clk cell_1478 ( .C ( clk ), .D ( signal_3566 ), .Q ( signal_3567 ) ) ;
    buf_clk cell_1480 ( .C ( clk ), .D ( signal_3568 ), .Q ( signal_3569 ) ) ;
    buf_clk cell_1482 ( .C ( clk ), .D ( signal_3570 ), .Q ( signal_3571 ) ) ;
    buf_clk cell_1484 ( .C ( clk ), .D ( signal_3572 ), .Q ( signal_3573 ) ) ;
    buf_clk cell_1486 ( .C ( clk ), .D ( signal_3574 ), .Q ( signal_3575 ) ) ;
    buf_clk cell_1488 ( .C ( clk ), .D ( signal_3576 ), .Q ( signal_3577 ) ) ;
    buf_clk cell_1490 ( .C ( clk ), .D ( signal_3578 ), .Q ( signal_3579 ) ) ;
    buf_clk cell_1492 ( .C ( clk ), .D ( signal_3580 ), .Q ( signal_3581 ) ) ;
    buf_clk cell_1494 ( .C ( clk ), .D ( signal_3582 ), .Q ( signal_3583 ) ) ;
    buf_clk cell_1496 ( .C ( clk ), .D ( signal_3584 ), .Q ( signal_3585 ) ) ;
    buf_clk cell_1498 ( .C ( clk ), .D ( signal_3586 ), .Q ( signal_3587 ) ) ;
    buf_clk cell_1500 ( .C ( clk ), .D ( signal_3588 ), .Q ( signal_3589 ) ) ;
    buf_clk cell_1502 ( .C ( clk ), .D ( signal_3590 ), .Q ( signal_3591 ) ) ;
    buf_clk cell_1504 ( .C ( clk ), .D ( signal_3592 ), .Q ( signal_3593 ) ) ;
    buf_clk cell_1506 ( .C ( clk ), .D ( signal_3594 ), .Q ( signal_3595 ) ) ;
    buf_clk cell_1508 ( .C ( clk ), .D ( signal_3596 ), .Q ( signal_3597 ) ) ;
    buf_clk cell_1510 ( .C ( clk ), .D ( signal_3598 ), .Q ( signal_3599 ) ) ;
    buf_clk cell_1512 ( .C ( clk ), .D ( signal_3600 ), .Q ( signal_3601 ) ) ;
    buf_clk cell_1514 ( .C ( clk ), .D ( signal_3602 ), .Q ( signal_3603 ) ) ;
    buf_clk cell_1516 ( .C ( clk ), .D ( signal_3604 ), .Q ( signal_3605 ) ) ;
    buf_clk cell_1518 ( .C ( clk ), .D ( signal_3606 ), .Q ( signal_3607 ) ) ;
    buf_clk cell_1520 ( .C ( clk ), .D ( signal_3608 ), .Q ( signal_3609 ) ) ;
    buf_clk cell_1522 ( .C ( clk ), .D ( signal_3610 ), .Q ( signal_3611 ) ) ;
    buf_clk cell_1524 ( .C ( clk ), .D ( signal_3612 ), .Q ( signal_3613 ) ) ;
    buf_clk cell_1526 ( .C ( clk ), .D ( signal_3614 ), .Q ( signal_3615 ) ) ;
    buf_clk cell_1528 ( .C ( clk ), .D ( signal_3616 ), .Q ( signal_3617 ) ) ;
    buf_clk cell_1534 ( .C ( clk ), .D ( signal_3622 ), .Q ( signal_3623 ) ) ;
    buf_clk cell_1542 ( .C ( clk ), .D ( signal_3630 ), .Q ( signal_3631 ) ) ;
    buf_clk cell_1550 ( .C ( clk ), .D ( signal_3638 ), .Q ( signal_3639 ) ) ;
    buf_clk cell_1564 ( .C ( clk ), .D ( signal_3652 ), .Q ( signal_3653 ) ) ;
    buf_clk cell_1574 ( .C ( clk ), .D ( signal_3662 ), .Q ( signal_3663 ) ) ;
    buf_clk cell_1584 ( .C ( clk ), .D ( signal_3672 ), .Q ( signal_3673 ) ) ;
    buf_clk cell_1594 ( .C ( clk ), .D ( signal_3682 ), .Q ( signal_3683 ) ) ;
    buf_clk cell_1606 ( .C ( clk ), .D ( signal_3694 ), .Q ( signal_3695 ) ) ;
    buf_clk cell_1618 ( .C ( clk ), .D ( signal_3706 ), .Q ( signal_3707 ) ) ;
    buf_clk cell_1630 ( .C ( clk ), .D ( signal_3718 ), .Q ( signal_3719 ) ) ;
    buf_clk cell_1644 ( .C ( clk ), .D ( signal_3732 ), .Q ( signal_3733 ) ) ;
    buf_clk cell_1658 ( .C ( clk ), .D ( signal_3746 ), .Q ( signal_3747 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_1535 ( .C ( clk ), .D ( signal_3623 ), .Q ( signal_3624 ) ) ;
    buf_clk cell_1543 ( .C ( clk ), .D ( signal_3631 ), .Q ( signal_3632 ) ) ;
    buf_clk cell_1551 ( .C ( clk ), .D ( signal_3639 ), .Q ( signal_3640 ) ) ;
    buf_clk cell_1553 ( .C ( clk ), .D ( signal_1102 ), .Q ( signal_3642 ) ) ;
    buf_clk cell_1555 ( .C ( clk ), .D ( signal_1672 ), .Q ( signal_3644 ) ) ;
    buf_clk cell_1557 ( .C ( clk ), .D ( signal_1673 ), .Q ( signal_3646 ) ) ;
    buf_clk cell_1565 ( .C ( clk ), .D ( signal_3653 ), .Q ( signal_3654 ) ) ;
    buf_clk cell_1575 ( .C ( clk ), .D ( signal_3663 ), .Q ( signal_3664 ) ) ;
    buf_clk cell_1585 ( .C ( clk ), .D ( signal_3673 ), .Q ( signal_3674 ) ) ;
    buf_clk cell_1595 ( .C ( clk ), .D ( signal_3683 ), .Q ( signal_3684 ) ) ;
    buf_clk cell_1607 ( .C ( clk ), .D ( signal_3695 ), .Q ( signal_3696 ) ) ;
    buf_clk cell_1619 ( .C ( clk ), .D ( signal_3707 ), .Q ( signal_3708 ) ) ;
    buf_clk cell_1631 ( .C ( clk ), .D ( signal_3719 ), .Q ( signal_3720 ) ) ;
    buf_clk cell_1645 ( .C ( clk ), .D ( signal_3733 ), .Q ( signal_3734 ) ) ;
    buf_clk cell_1659 ( .C ( clk ), .D ( signal_3747 ), .Q ( signal_3748 ) ) ;

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1090 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1413, signal_1412, signal_973}), .a ({signal_1411, signal_1410, signal_972}), .clk ( clk ), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({signal_1679, signal_1678, signal_1105}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1091 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1417, signal_1416, signal_975}), .a ({signal_1415, signal_1414, signal_974}), .clk ( clk ), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({signal_1681, signal_1680, signal_1106}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1092 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1421, signal_1420, signal_977}), .a ({signal_1419, signal_1418, signal_976}), .clk ( clk ), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({signal_1683, signal_1682, signal_1107}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1093 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1425, signal_1424, signal_979}), .a ({signal_1423, signal_1422, signal_978}), .clk ( clk ), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({signal_1685, signal_1684, signal_1108}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1094 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1429, signal_1428, signal_981}), .a ({signal_1427, signal_1426, signal_980}), .clk ( clk ), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({signal_1687, signal_1686, signal_1109}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1095 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1427, signal_1426, signal_980}), .a ({signal_1431, signal_1430, signal_982}), .clk ( clk ), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({signal_1689, signal_1688, signal_1110}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1096 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1433, signal_1432, signal_983}), .a ({signal_3491, signal_3489, signal_3487}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({signal_1691, signal_1690, signal_1111}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1097 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1437, signal_1436, signal_985}), .a ({signal_1435, signal_1434, signal_984}), .clk ( clk ), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_1693, signal_1692, signal_1112}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1098 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1441, signal_1440, signal_987}), .a ({signal_1439, signal_1438, signal_986}), .clk ( clk ), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({signal_1695, signal_1694, signal_1113}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1099 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3497, signal_3495, signal_3493}), .a ({signal_1443, signal_1442, signal_988}), .clk ( clk ), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({signal_1697, signal_1696, signal_1114}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1100 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1447, signal_1446, signal_990}), .a ({signal_1445, signal_1444, signal_989}), .clk ( clk ), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({signal_1699, signal_1698, signal_1115}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1101 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1449, signal_1448, signal_991}), .a ({signal_1423, signal_1422, signal_978}), .clk ( clk ), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({signal_1701, signal_1700, signal_1116}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1102 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1453, signal_1452, signal_993}), .a ({signal_1451, signal_1450, signal_992}), .clk ( clk ), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({signal_1703, signal_1702, signal_1117}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1103 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1457, signal_1456, signal_995}), .a ({signal_1455, signal_1454, signal_994}), .clk ( clk ), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({signal_1705, signal_1704, signal_1118}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1104 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1461, signal_1460, signal_997}), .a ({signal_1459, signal_1458, signal_996}), .clk ( clk ), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({signal_1707, signal_1706, signal_1119}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1105 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1465, signal_1464, signal_999}), .a ({signal_1463, signal_1462, signal_998}), .clk ( clk ), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({signal_1709, signal_1708, signal_1120}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1106 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1469, signal_1468, signal_1001}), .a ({signal_1467, signal_1466, signal_1000}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({signal_1711, signal_1710, signal_1121}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1107 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1473, signal_1472, signal_1003}), .a ({signal_1471, signal_1470, signal_1002}), .clk ( clk ), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_1713, signal_1712, signal_1122}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1108 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1435, signal_1434, signal_984}), .a ({signal_1475, signal_1474, signal_1004}), .clk ( clk ), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({signal_1715, signal_1714, signal_1123}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1109 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1479, signal_1478, signal_1006}), .a ({signal_1477, signal_1476, signal_1005}), .clk ( clk ), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({signal_1717, signal_1716, signal_1124}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1110 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1483, signal_1482, signal_1008}), .a ({signal_1481, signal_1480, signal_1007}), .clk ( clk ), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({signal_1719, signal_1718, signal_1125}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1111 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1487, signal_1486, signal_1010}), .a ({signal_1485, signal_1484, signal_1009}), .clk ( clk ), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({signal_1721, signal_1720, signal_1126}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1112 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1489, signal_1488, signal_1011}), .a ({signal_3503, signal_3501, signal_3499}), .clk ( clk ), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({signal_1723, signal_1722, signal_1127}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1113 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1493, signal_1492, signal_1013}), .a ({signal_1491, signal_1490, signal_1012}), .clk ( clk ), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({signal_1725, signal_1724, signal_1128}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1114 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1497, signal_1496, signal_1015}), .a ({signal_1495, signal_1494, signal_1014}), .clk ( clk ), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({signal_1727, signal_1726, signal_1129}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1115 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1501, signal_1500, signal_1017}), .a ({signal_1499, signal_1498, signal_1016}), .clk ( clk ), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({signal_1729, signal_1728, signal_1130}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1116 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1503, signal_1502, signal_1018}), .a ({signal_1471, signal_1470, signal_1002}), .clk ( clk ), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({signal_1731, signal_1730, signal_1131}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1117 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1423, signal_1422, signal_978}), .a ({signal_1419, signal_1418, signal_976}), .clk ( clk ), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_1733, signal_1732, signal_1132}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1118 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1507, signal_1506, signal_1020}), .a ({signal_1505, signal_1504, signal_1019}), .clk ( clk ), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({signal_1735, signal_1734, signal_1133}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1119 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1509, signal_1508, signal_1021}), .a ({1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({signal_1737, signal_1736, signal_1134}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1120 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3509, signal_3507, signal_3505}), .a ({signal_1499, signal_1498, signal_1016}), .clk ( clk ), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({signal_1739, signal_1738, signal_1135}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1121 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1509, signal_1508, signal_1021}), .a ({signal_3515, signal_3513, signal_3511}), .clk ( clk ), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({signal_1741, signal_1740, signal_1136}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1122 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1417, signal_1416, signal_975}), .a ({signal_3521, signal_3519, signal_3517}), .clk ( clk ), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({signal_1743, signal_1742, signal_1137}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1123 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3491, signal_3489, signal_3487}), .a ({signal_1511, signal_1510, signal_1022}), .clk ( clk ), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({signal_1745, signal_1744, signal_1138}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1124 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1515, signal_1514, signal_1024}), .a ({signal_1513, signal_1512, signal_1023}), .clk ( clk ), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({signal_1747, signal_1746, signal_1139}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1125 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3515, signal_3513, signal_3511}), .a ({signal_1487, signal_1486, signal_1010}), .clk ( clk ), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({signal_1749, signal_1748, signal_1140}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1126 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1509, signal_1508, signal_1021}), .a ({signal_1517, signal_1516, signal_1025}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({signal_1751, signal_1750, signal_1141}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1127 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1521, signal_1520, signal_1027}), .a ({signal_1519, signal_1518, signal_1026}), .clk ( clk ), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_1753, signal_1752, signal_1142}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1128 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3527, signal_3525, signal_3523}), .a ({signal_1523, signal_1522, signal_1028}), .clk ( clk ), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({signal_1755, signal_1754, signal_1143}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1129 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1525, signal_1524, signal_1029}), .a ({signal_3533, signal_3531, signal_3529}), .clk ( clk ), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({signal_1757, signal_1756, signal_1144}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1130 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1529, signal_1528, signal_1031}), .a ({signal_1527, signal_1526, signal_1030}), .clk ( clk ), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({signal_1759, signal_1758, signal_1145}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1131 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1533, signal_1532, signal_1033}), .a ({signal_1531, signal_1530, signal_1032}), .clk ( clk ), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({signal_1761, signal_1760, signal_1146}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1132 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1537, signal_1536, signal_1035}), .a ({signal_1535, signal_1534, signal_1034}), .clk ( clk ), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({signal_1763, signal_1762, signal_1147}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1133 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1421, signal_1420, signal_977}), .a ({signal_1539, signal_1538, signal_1036}), .clk ( clk ), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({signal_1765, signal_1764, signal_1148}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1134 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1543, signal_1542, signal_1038}), .a ({signal_1541, signal_1540, signal_1037}), .clk ( clk ), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({signal_1767, signal_1766, signal_1149}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1135 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1525, signal_1524, signal_1029}), .a ({signal_1545, signal_1544, signal_1039}), .clk ( clk ), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({signal_1769, signal_1768, signal_1150}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1136 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1547, signal_1546, signal_1040}), .a ({signal_1523, signal_1522, signal_1028}), .clk ( clk ), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({signal_1771, signal_1770, signal_1151}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1137 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1549, signal_1548, signal_1041}), .a ({signal_1493, signal_1492, signal_1013}), .clk ( clk ), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_1773, signal_1772, signal_1152}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1138 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1551, signal_1550, signal_1042}), .a ({signal_1453, signal_1452, signal_993}), .clk ( clk ), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({signal_1775, signal_1774, signal_1153}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1139 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1555, signal_1554, signal_1044}), .a ({signal_1553, signal_1552, signal_1043}), .clk ( clk ), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({signal_1777, signal_1776, signal_1154}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1140 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1557, signal_1556, signal_1045}), .a ({signal_1467, signal_1466, signal_1000}), .clk ( clk ), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({signal_1779, signal_1778, signal_1155}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1141 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1559, signal_1558, signal_1046}), .a ({signal_1525, signal_1524, signal_1029}), .clk ( clk ), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({signal_1781, signal_1780, signal_1156}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1142 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1563, signal_1562, signal_1048}), .a ({signal_1561, signal_1560, signal_1047}), .clk ( clk ), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({signal_1783, signal_1782, signal_1157}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1143 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1567, signal_1566, signal_1050}), .a ({signal_1565, signal_1564, signal_1049}), .clk ( clk ), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({signal_1785, signal_1784, signal_1158}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1144 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3521, signal_3519, signal_3517}), .a ({signal_1569, signal_1568, signal_1051}), .clk ( clk ), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({signal_1787, signal_1786, signal_1159}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1145 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1559, signal_1558, signal_1046}), .a ({signal_1461, signal_1460, signal_997}), .clk ( clk ), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({signal_1789, signal_1788, signal_1160}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1146 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1439, signal_1438, signal_986}), .a ({signal_1571, signal_1570, signal_1052}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({signal_1791, signal_1790, signal_1161}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1147 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1487, signal_1486, signal_1010}), .a ({signal_1435, signal_1434, signal_984}), .clk ( clk ), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_1793, signal_1792, signal_1162}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1148 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1529, signal_1528, signal_1031}), .a ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({signal_1795, signal_1794, signal_1163}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1149 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1509, signal_1508, signal_1021}), .a ({signal_1573, signal_1572, signal_1053}), .clk ( clk ), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({signal_1797, signal_1796, signal_1164}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1150 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1575, signal_1574, signal_1054}), .a ({signal_1427, signal_1426, signal_980}), .clk ( clk ), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({signal_1799, signal_1798, signal_1165}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1151 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1533, signal_1532, signal_1033}), .a ({signal_1577, signal_1576, signal_1055}), .clk ( clk ), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({signal_1801, signal_1800, signal_1166}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1152 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1581, signal_1580, signal_1057}), .a ({signal_1579, signal_1578, signal_1056}), .clk ( clk ), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({signal_1803, signal_1802, signal_1167}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1153 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1481, signal_1480, signal_1007}), .a ({signal_1583, signal_1582, signal_1058}), .clk ( clk ), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({signal_1805, signal_1804, signal_1168}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1154 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1427, signal_1426, signal_980}), .a ({signal_1585, signal_1584, signal_1059}), .clk ( clk ), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({signal_1807, signal_1806, signal_1169}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1155 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1507, signal_1506, signal_1020}), .a ({signal_3539, signal_3537, signal_3535}), .clk ( clk ), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({signal_1809, signal_1808, signal_1170}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1156 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1587, signal_1586, signal_1060}), .a ({signal_1515, signal_1514, signal_1024}), .clk ( clk ), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({signal_1811, signal_1810, signal_1171}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1157 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3509, signal_3507, signal_3505}), .a ({signal_1487, signal_1486, signal_1010}), .clk ( clk ), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_1813, signal_1812, signal_1172}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1158 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1421, signal_1420, signal_977}), .a ({signal_1589, signal_1588, signal_1061}), .clk ( clk ), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({signal_1815, signal_1814, signal_1173}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1159 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1491, signal_1490, signal_1012}), .a ({signal_1431, signal_1430, signal_982}), .clk ( clk ), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({signal_1817, signal_1816, signal_1174}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1160 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1547, signal_1546, signal_1040}), .a ({signal_1591, signal_1590, signal_1062}), .clk ( clk ), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({signal_1819, signal_1818, signal_1175}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1161 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1493, signal_1492, signal_1013}), .a ({signal_1593, signal_1592, signal_1063}), .clk ( clk ), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({signal_1821, signal_1820, signal_1176}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1162 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1597, signal_1596, signal_1065}), .a ({signal_1595, signal_1594, signal_1064}), .clk ( clk ), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({signal_1823, signal_1822, signal_1177}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1163 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1599, signal_1598, signal_1066}), .a ({signal_1423, signal_1422, signal_978}), .clk ( clk ), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({signal_1825, signal_1824, signal_1178}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1164 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1601, signal_1600, signal_1067}), .a ({signal_1499, signal_1498, signal_1016}), .clk ( clk ), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({signal_1827, signal_1826, signal_1179}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1165 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1583, signal_1582, signal_1058}), .a ({signal_3551, signal_3547, signal_3543}), .clk ( clk ), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({signal_1829, signal_1828, signal_1180}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1166 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1605, signal_1604, signal_1069}), .a ({signal_1603, signal_1602, signal_1068}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({signal_1831, signal_1830, signal_1181}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1167 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3557, signal_3555, signal_3553}), .a ({signal_1607, signal_1606, signal_1070}), .clk ( clk ), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_1833, signal_1832, signal_1182}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1168 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1609, signal_1608, signal_1071}), .a ({signal_1573, signal_1572, signal_1053}), .clk ( clk ), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({signal_1835, signal_1834, signal_1183}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1169 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1413, signal_1412, signal_973}), .a ({signal_1451, signal_1450, signal_992}), .clk ( clk ), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({signal_1837, signal_1836, signal_1184}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1170 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1431, signal_1430, signal_982}), .a ({signal_1611, signal_1610, signal_1072}), .clk ( clk ), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({signal_1839, signal_1838, signal_1185}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1171 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1449, signal_1448, signal_991}), .a ({signal_1547, signal_1546, signal_1040}), .clk ( clk ), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({signal_1841, signal_1840, signal_1186}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1172 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1411, signal_1410, signal_972}), .a ({signal_1485, signal_1484, signal_1009}), .clk ( clk ), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({signal_1843, signal_1842, signal_1187}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1173 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1419, signal_1418, signal_976}), .a ({signal_1571, signal_1570, signal_1052}), .clk ( clk ), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({signal_1845, signal_1844, signal_1188}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1174 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1613, signal_1612, signal_1073}), .a ({signal_1509, signal_1508, signal_1021}), .clk ( clk ), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({signal_1847, signal_1846, signal_1189}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1175 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1587, signal_1586, signal_1060}), .a ({signal_3563, signal_3561, signal_3559}), .clk ( clk ), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({signal_1849, signal_1848, signal_1190}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1176 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1615, signal_1614, signal_1074}), .a ({signal_1433, signal_1432, signal_983}), .clk ( clk ), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({signal_1851, signal_1850, signal_1191}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1177 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1619, signal_1618, signal_1076}), .a ({signal_1617, signal_1616, signal_1075}), .clk ( clk ), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_1853, signal_1852, signal_1192}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1178 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1603, signal_1602, signal_1068}), .a ({signal_1621, signal_1620, signal_1077}), .clk ( clk ), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({signal_1855, signal_1854, signal_1193}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1179 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1453, signal_1452, signal_993}), .a ({signal_3569, signal_3567, signal_3565}), .clk ( clk ), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({signal_1857, signal_1856, signal_1194}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1180 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1625, signal_1624, signal_1079}), .a ({signal_1623, signal_1622, signal_1078}), .clk ( clk ), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({signal_1859, signal_1858, signal_1195}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1181 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1535, signal_1534, signal_1034}), .a ({signal_1423, signal_1422, signal_978}), .clk ( clk ), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({signal_1861, signal_1860, signal_1196}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1182 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1425, signal_1424, signal_979}), .a ({signal_1627, signal_1626, signal_1080}), .clk ( clk ), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({signal_1863, signal_1862, signal_1197}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1183 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1505, signal_1504, signal_1019}), .a ({signal_3575, signal_3573, signal_3571}), .clk ( clk ), .r ({Fresh[770], Fresh[769], Fresh[768]}), .c ({signal_1865, signal_1864, signal_1198}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1184 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1631, signal_1630, signal_1082}), .a ({signal_1629, signal_1628, signal_1081}), .clk ( clk ), .r ({Fresh[773], Fresh[772], Fresh[771]}), .c ({signal_1867, signal_1866, signal_1199}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1185 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1633, signal_1632, signal_1083}), .a ({signal_3581, signal_3579, signal_3577}), .clk ( clk ), .r ({Fresh[776], Fresh[775], Fresh[774]}), .c ({signal_1869, signal_1868, signal_1200}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1186 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1521, signal_1520, signal_1027}), .a ({signal_1635, signal_1634, signal_1084}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777]}), .c ({signal_1871, signal_1870, signal_1201}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1187 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3587, signal_3585, signal_3583}), .a ({signal_1609, signal_1608, signal_1071}), .clk ( clk ), .r ({Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_1873, signal_1872, signal_1202}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1188 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1637, signal_1636, signal_1085}), .a ({signal_1571, signal_1570, signal_1052}), .clk ( clk ), .r ({Fresh[785], Fresh[784], Fresh[783]}), .c ({signal_1875, signal_1874, signal_1203}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1189 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1641, signal_1640, signal_1087}), .a ({signal_1639, signal_1638, signal_1086}), .clk ( clk ), .r ({Fresh[788], Fresh[787], Fresh[786]}), .c ({signal_1877, signal_1876, signal_1204}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1190 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1621, signal_1620, signal_1077}), .a ({signal_3533, signal_3531, signal_3529}), .clk ( clk ), .r ({Fresh[791], Fresh[790], Fresh[789]}), .c ({signal_1879, signal_1878, signal_1205}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1191 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1643, signal_1642, signal_1088}), .a ({signal_1447, signal_1446, signal_990}), .clk ( clk ), .r ({Fresh[794], Fresh[793], Fresh[792]}), .c ({signal_1881, signal_1880, signal_1206}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1192 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1623, signal_1622, signal_1078}), .a ({signal_1645, signal_1644, signal_1089}), .clk ( clk ), .r ({Fresh[797], Fresh[796], Fresh[795]}), .c ({signal_1883, signal_1882, signal_1207}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1193 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1637, signal_1636, signal_1085}), .a ({signal_1437, signal_1436, signal_985}), .clk ( clk ), .r ({Fresh[800], Fresh[799], Fresh[798]}), .c ({signal_1885, signal_1884, signal_1208}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1194 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1649, signal_1648, signal_1091}), .a ({signal_1647, signal_1646, signal_1090}), .clk ( clk ), .r ({Fresh[803], Fresh[802], Fresh[801]}), .c ({signal_1887, signal_1886, signal_1209}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1195 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1523, signal_1522, signal_1028}), .a ({signal_1559, signal_1558, signal_1046}), .clk ( clk ), .r ({Fresh[806], Fresh[805], Fresh[804]}), .c ({signal_1889, signal_1888, signal_1210}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1196 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1441, signal_1440, signal_987}), .a ({signal_3503, signal_3501, signal_3499}), .clk ( clk ), .r ({Fresh[809], Fresh[808], Fresh[807]}), .c ({signal_1891, signal_1890, signal_1211}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1197 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1651, signal_1650, signal_1092}), .a ({signal_1571, signal_1570, signal_1052}), .clk ( clk ), .r ({Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_1893, signal_1892, signal_1212}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1198 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3593, signal_3591, signal_3589}), .a ({signal_1631, signal_1630, signal_1082}), .clk ( clk ), .r ({Fresh[815], Fresh[814], Fresh[813]}), .c ({signal_1895, signal_1894, signal_1213}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1199 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1603, signal_1602, signal_1068}), .a ({signal_3599, signal_3597, signal_3595}), .clk ( clk ), .r ({Fresh[818], Fresh[817], Fresh[816]}), .c ({signal_1897, signal_1896, signal_1214}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1200 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1653, signal_1652, signal_1093}), .a ({signal_1603, signal_1602, signal_1068}), .clk ( clk ), .r ({Fresh[821], Fresh[820], Fresh[819]}), .c ({signal_1899, signal_1898, signal_1215}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1201 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_1493, signal_1492, signal_1013}), .clk ( clk ), .r ({Fresh[824], Fresh[823], Fresh[822]}), .c ({signal_1901, signal_1900, signal_1216}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1202 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1655, signal_1654, signal_1094}), .a ({signal_1573, signal_1572, signal_1053}), .clk ( clk ), .r ({Fresh[827], Fresh[826], Fresh[825]}), .c ({signal_1903, signal_1902, signal_1217}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1203 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1657, signal_1656, signal_1095}), .a ({signal_1551, signal_1550, signal_1042}), .clk ( clk ), .r ({Fresh[830], Fresh[829], Fresh[828]}), .c ({signal_1905, signal_1904, signal_1218}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1204 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3605, signal_3603, signal_3601}), .a ({signal_1609, signal_1608, signal_1071}), .clk ( clk ), .r ({Fresh[833], Fresh[832], Fresh[831]}), .c ({signal_1907, signal_1906, signal_1219}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1205 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1659, signal_1658, signal_1096}), .a ({signal_1601, signal_1600, signal_1067}), .clk ( clk ), .r ({Fresh[836], Fresh[835], Fresh[834]}), .c ({signal_1909, signal_1908, signal_1220}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1206 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1645, signal_1644, signal_1089}), .a ({signal_1499, signal_1498, signal_1016}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837]}), .c ({signal_1911, signal_1910, signal_1221}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1207 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1661, signal_1660, signal_1097}), .a ({signal_3557, signal_3555, signal_3553}), .clk ( clk ), .r ({Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_1913, signal_1912, signal_1222}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1208 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_3611, signal_3609, signal_3607}), .a ({signal_1663, signal_1662, signal_1098}), .clk ( clk ), .r ({Fresh[845], Fresh[844], Fresh[843]}), .c ({signal_1915, signal_1914, signal_1223}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1209 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1665, signal_1664, signal_1099}), .a ({signal_3617, signal_3615, signal_3613}), .clk ( clk ), .r ({Fresh[848], Fresh[847], Fresh[846]}), .c ({signal_1917, signal_1916, signal_1224}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1210 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1667, signal_1666, signal_1100}), .a ({signal_1657, signal_1656, signal_1095}), .clk ( clk ), .r ({Fresh[851], Fresh[850], Fresh[849]}), .c ({signal_1919, signal_1918, signal_1225}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1211 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1669, signal_1668, signal_1101}), .a ({signal_1603, signal_1602, signal_1068}), .clk ( clk ), .r ({Fresh[854], Fresh[853], Fresh[852]}), .c ({signal_1921, signal_1920, signal_1226}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1212 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1481, signal_1480, signal_1007}), .a ({signal_1491, signal_1490, signal_1012}), .clk ( clk ), .r ({Fresh[857], Fresh[856], Fresh[855]}), .c ({signal_1923, signal_1922, signal_1227}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1213 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1641, signal_1640, signal_1087}), .a ({signal_3521, signal_3519, signal_3517}), .clk ( clk ), .r ({Fresh[860], Fresh[859], Fresh[858]}), .c ({signal_1925, signal_1924, signal_1228}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1214 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1675, signal_1674, signal_1103}), .a ({signal_1487, signal_1486, signal_1010}), .clk ( clk ), .r ({Fresh[863], Fresh[862], Fresh[861]}), .c ({signal_1927, signal_1926, signal_1229}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1215 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1471, signal_1470, signal_1002}), .a ({signal_1677, signal_1676, signal_1104}), .clk ( clk ), .r ({Fresh[866], Fresh[865], Fresh[864]}), .c ({signal_1929, signal_1928, signal_1230}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1216 ( .s ({signal_3485, signal_3483, signal_3481}), .b ({signal_1575, signal_1574, signal_1054}), .a ({signal_1469, signal_1468, signal_1001}), .clk ( clk ), .r ({Fresh[869], Fresh[868], Fresh[867]}), .c ({signal_1931, signal_1930, signal_1231}) ) ;
    buf_clk cell_1536 ( .C ( clk ), .D ( signal_3624 ), .Q ( signal_3625 ) ) ;
    buf_clk cell_1544 ( .C ( clk ), .D ( signal_3632 ), .Q ( signal_3633 ) ) ;
    buf_clk cell_1552 ( .C ( clk ), .D ( signal_3640 ), .Q ( signal_3641 ) ) ;
    buf_clk cell_1554 ( .C ( clk ), .D ( signal_3642 ), .Q ( signal_3643 ) ) ;
    buf_clk cell_1556 ( .C ( clk ), .D ( signal_3644 ), .Q ( signal_3645 ) ) ;
    buf_clk cell_1558 ( .C ( clk ), .D ( signal_3646 ), .Q ( signal_3647 ) ) ;
    buf_clk cell_1566 ( .C ( clk ), .D ( signal_3654 ), .Q ( signal_3655 ) ) ;
    buf_clk cell_1576 ( .C ( clk ), .D ( signal_3664 ), .Q ( signal_3665 ) ) ;
    buf_clk cell_1586 ( .C ( clk ), .D ( signal_3674 ), .Q ( signal_3675 ) ) ;
    buf_clk cell_1596 ( .C ( clk ), .D ( signal_3684 ), .Q ( signal_3685 ) ) ;
    buf_clk cell_1608 ( .C ( clk ), .D ( signal_3696 ), .Q ( signal_3697 ) ) ;
    buf_clk cell_1620 ( .C ( clk ), .D ( signal_3708 ), .Q ( signal_3709 ) ) ;
    buf_clk cell_1632 ( .C ( clk ), .D ( signal_3720 ), .Q ( signal_3721 ) ) ;
    buf_clk cell_1646 ( .C ( clk ), .D ( signal_3734 ), .Q ( signal_3735 ) ) ;
    buf_clk cell_1660 ( .C ( clk ), .D ( signal_3748 ), .Q ( signal_3749 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_1567 ( .C ( clk ), .D ( signal_3655 ), .Q ( signal_3656 ) ) ;
    buf_clk cell_1577 ( .C ( clk ), .D ( signal_3665 ), .Q ( signal_3666 ) ) ;
    buf_clk cell_1587 ( .C ( clk ), .D ( signal_3675 ), .Q ( signal_3676 ) ) ;
    buf_clk cell_1597 ( .C ( clk ), .D ( signal_3685 ), .Q ( signal_3686 ) ) ;
    buf_clk cell_1609 ( .C ( clk ), .D ( signal_3697 ), .Q ( signal_3698 ) ) ;
    buf_clk cell_1621 ( .C ( clk ), .D ( signal_3709 ), .Q ( signal_3710 ) ) ;
    buf_clk cell_1633 ( .C ( clk ), .D ( signal_3721 ), .Q ( signal_3722 ) ) ;
    buf_clk cell_1647 ( .C ( clk ), .D ( signal_3735 ), .Q ( signal_3736 ) ) ;
    buf_clk cell_1661 ( .C ( clk ), .D ( signal_3749 ), .Q ( signal_3750 ) ) ;

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1217 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1681, signal_1680, signal_1106}), .a ({signal_1679, signal_1678, signal_1105}), .clk ( clk ), .r ({Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_1935, signal_1934, signal_1232}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1218 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1685, signal_1684, signal_1108}), .a ({signal_1683, signal_1682, signal_1107}), .clk ( clk ), .r ({Fresh[875], Fresh[874], Fresh[873]}), .c ({signal_1937, signal_1936, signal_1233}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1219 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1689, signal_1688, signal_1110}), .a ({signal_1687, signal_1686, signal_1109}), .clk ( clk ), .r ({Fresh[878], Fresh[877], Fresh[876]}), .c ({signal_1939, signal_1938, signal_1234}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1220 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1693, signal_1692, signal_1112}), .a ({signal_1691, signal_1690, signal_1111}), .clk ( clk ), .r ({Fresh[881], Fresh[880], Fresh[879]}), .c ({signal_1941, signal_1940, signal_1235}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1221 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1697, signal_1696, signal_1114}), .a ({signal_1695, signal_1694, signal_1113}), .clk ( clk ), .r ({Fresh[884], Fresh[883], Fresh[882]}), .c ({signal_1943, signal_1942, signal_1236}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1222 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1701, signal_1700, signal_1116}), .a ({signal_1699, signal_1698, signal_1115}), .clk ( clk ), .r ({Fresh[887], Fresh[886], Fresh[885]}), .c ({signal_1945, signal_1944, signal_1237}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1223 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1705, signal_1704, signal_1118}), .a ({signal_1703, signal_1702, signal_1117}), .clk ( clk ), .r ({Fresh[890], Fresh[889], Fresh[888]}), .c ({signal_1947, signal_1946, signal_1238}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1224 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1709, signal_1708, signal_1120}), .a ({signal_1707, signal_1706, signal_1119}), .clk ( clk ), .r ({Fresh[893], Fresh[892], Fresh[891]}), .c ({signal_1949, signal_1948, signal_1239}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1225 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1713, signal_1712, signal_1122}), .a ({signal_1711, signal_1710, signal_1121}), .clk ( clk ), .r ({Fresh[896], Fresh[895], Fresh[894]}), .c ({signal_1951, signal_1950, signal_1240}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1226 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1717, signal_1716, signal_1124}), .a ({signal_1715, signal_1714, signal_1123}), .clk ( clk ), .r ({Fresh[899], Fresh[898], Fresh[897]}), .c ({signal_1953, signal_1952, signal_1241}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1227 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1721, signal_1720, signal_1126}), .a ({signal_1719, signal_1718, signal_1125}), .clk ( clk ), .r ({Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_1955, signal_1954, signal_1242}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1228 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1725, signal_1724, signal_1128}), .a ({signal_1723, signal_1722, signal_1127}), .clk ( clk ), .r ({Fresh[905], Fresh[904], Fresh[903]}), .c ({signal_1957, signal_1956, signal_1243}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1229 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1729, signal_1728, signal_1130}), .a ({signal_1727, signal_1726, signal_1129}), .clk ( clk ), .r ({Fresh[908], Fresh[907], Fresh[906]}), .c ({signal_1959, signal_1958, signal_1244}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1230 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1733, signal_1732, signal_1132}), .a ({signal_1731, signal_1730, signal_1131}), .clk ( clk ), .r ({Fresh[911], Fresh[910], Fresh[909]}), .c ({signal_1961, signal_1960, signal_1245}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1231 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1737, signal_1736, signal_1134}), .a ({signal_1735, signal_1734, signal_1133}), .clk ( clk ), .r ({Fresh[914], Fresh[913], Fresh[912]}), .c ({signal_1963, signal_1962, signal_1246}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1232 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1741, signal_1740, signal_1136}), .a ({signal_1739, signal_1738, signal_1135}), .clk ( clk ), .r ({Fresh[917], Fresh[916], Fresh[915]}), .c ({signal_1965, signal_1964, signal_1247}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1233 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1745, signal_1744, signal_1138}), .a ({signal_1743, signal_1742, signal_1137}), .clk ( clk ), .r ({Fresh[920], Fresh[919], Fresh[918]}), .c ({signal_1967, signal_1966, signal_1248}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1234 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1749, signal_1748, signal_1140}), .a ({signal_1747, signal_1746, signal_1139}), .clk ( clk ), .r ({Fresh[923], Fresh[922], Fresh[921]}), .c ({signal_1969, signal_1968, signal_1249}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1235 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1753, signal_1752, signal_1142}), .a ({signal_1751, signal_1750, signal_1141}), .clk ( clk ), .r ({Fresh[926], Fresh[925], Fresh[924]}), .c ({signal_1971, signal_1970, signal_1250}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1236 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1757, signal_1756, signal_1144}), .a ({signal_1755, signal_1754, signal_1143}), .clk ( clk ), .r ({Fresh[929], Fresh[928], Fresh[927]}), .c ({signal_1973, signal_1972, signal_1251}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1237 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1761, signal_1760, signal_1146}), .a ({signal_1759, signal_1758, signal_1145}), .clk ( clk ), .r ({Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_1975, signal_1974, signal_1252}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1238 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1765, signal_1764, signal_1148}), .a ({signal_1763, signal_1762, signal_1147}), .clk ( clk ), .r ({Fresh[935], Fresh[934], Fresh[933]}), .c ({signal_1977, signal_1976, signal_1253}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1239 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1769, signal_1768, signal_1150}), .a ({signal_1767, signal_1766, signal_1149}), .clk ( clk ), .r ({Fresh[938], Fresh[937], Fresh[936]}), .c ({signal_1979, signal_1978, signal_1254}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1240 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1773, signal_1772, signal_1152}), .a ({signal_1771, signal_1770, signal_1151}), .clk ( clk ), .r ({Fresh[941], Fresh[940], Fresh[939]}), .c ({signal_1981, signal_1980, signal_1255}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1241 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1777, signal_1776, signal_1154}), .a ({signal_1775, signal_1774, signal_1153}), .clk ( clk ), .r ({Fresh[944], Fresh[943], Fresh[942]}), .c ({signal_1983, signal_1982, signal_1256}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1242 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1781, signal_1780, signal_1156}), .a ({signal_1779, signal_1778, signal_1155}), .clk ( clk ), .r ({Fresh[947], Fresh[946], Fresh[945]}), .c ({signal_1985, signal_1984, signal_1257}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1243 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1785, signal_1784, signal_1158}), .a ({signal_1783, signal_1782, signal_1157}), .clk ( clk ), .r ({Fresh[950], Fresh[949], Fresh[948]}), .c ({signal_1987, signal_1986, signal_1258}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1244 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1789, signal_1788, signal_1160}), .a ({signal_1787, signal_1786, signal_1159}), .clk ( clk ), .r ({Fresh[953], Fresh[952], Fresh[951]}), .c ({signal_1989, signal_1988, signal_1259}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1245 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1793, signal_1792, signal_1162}), .a ({signal_1791, signal_1790, signal_1161}), .clk ( clk ), .r ({Fresh[956], Fresh[955], Fresh[954]}), .c ({signal_1991, signal_1990, signal_1260}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1246 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1797, signal_1796, signal_1164}), .a ({signal_1795, signal_1794, signal_1163}), .clk ( clk ), .r ({Fresh[959], Fresh[958], Fresh[957]}), .c ({signal_1993, signal_1992, signal_1261}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1247 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1801, signal_1800, signal_1166}), .a ({signal_1799, signal_1798, signal_1165}), .clk ( clk ), .r ({Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_1995, signal_1994, signal_1262}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1248 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1805, signal_1804, signal_1168}), .a ({signal_1803, signal_1802, signal_1167}), .clk ( clk ), .r ({Fresh[965], Fresh[964], Fresh[963]}), .c ({signal_1997, signal_1996, signal_1263}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1249 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1809, signal_1808, signal_1170}), .a ({signal_1807, signal_1806, signal_1169}), .clk ( clk ), .r ({Fresh[968], Fresh[967], Fresh[966]}), .c ({signal_1999, signal_1998, signal_1264}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1250 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1813, signal_1812, signal_1172}), .a ({signal_1811, signal_1810, signal_1171}), .clk ( clk ), .r ({Fresh[971], Fresh[970], Fresh[969]}), .c ({signal_2001, signal_2000, signal_1265}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1251 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1817, signal_1816, signal_1174}), .a ({signal_1815, signal_1814, signal_1173}), .clk ( clk ), .r ({Fresh[974], Fresh[973], Fresh[972]}), .c ({signal_2003, signal_2002, signal_1266}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1252 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1821, signal_1820, signal_1176}), .a ({signal_1819, signal_1818, signal_1175}), .clk ( clk ), .r ({Fresh[977], Fresh[976], Fresh[975]}), .c ({signal_2005, signal_2004, signal_1267}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1253 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1825, signal_1824, signal_1178}), .a ({signal_1823, signal_1822, signal_1177}), .clk ( clk ), .r ({Fresh[980], Fresh[979], Fresh[978]}), .c ({signal_2007, signal_2006, signal_1268}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1254 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1829, signal_1828, signal_1180}), .a ({signal_1827, signal_1826, signal_1179}), .clk ( clk ), .r ({Fresh[983], Fresh[982], Fresh[981]}), .c ({signal_2009, signal_2008, signal_1269}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1255 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1833, signal_1832, signal_1182}), .a ({signal_1831, signal_1830, signal_1181}), .clk ( clk ), .r ({Fresh[986], Fresh[985], Fresh[984]}), .c ({signal_2011, signal_2010, signal_1270}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1256 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1837, signal_1836, signal_1184}), .a ({signal_1835, signal_1834, signal_1183}), .clk ( clk ), .r ({Fresh[989], Fresh[988], Fresh[987]}), .c ({signal_2013, signal_2012, signal_1271}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1257 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1841, signal_1840, signal_1186}), .a ({signal_1839, signal_1838, signal_1185}), .clk ( clk ), .r ({Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_2015, signal_2014, signal_1272}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1258 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1845, signal_1844, signal_1188}), .a ({signal_1843, signal_1842, signal_1187}), .clk ( clk ), .r ({Fresh[995], Fresh[994], Fresh[993]}), .c ({signal_2017, signal_2016, signal_1273}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1259 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1849, signal_1848, signal_1190}), .a ({signal_1847, signal_1846, signal_1189}), .clk ( clk ), .r ({Fresh[998], Fresh[997], Fresh[996]}), .c ({signal_2019, signal_2018, signal_1274}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1260 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1853, signal_1852, signal_1192}), .a ({signal_1851, signal_1850, signal_1191}), .clk ( clk ), .r ({Fresh[1001], Fresh[1000], Fresh[999]}), .c ({signal_2021, signal_2020, signal_1275}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1261 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1857, signal_1856, signal_1194}), .a ({signal_1855, signal_1854, signal_1193}), .clk ( clk ), .r ({Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({signal_2023, signal_2022, signal_1276}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1262 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1861, signal_1860, signal_1196}), .a ({signal_1859, signal_1858, signal_1195}), .clk ( clk ), .r ({Fresh[1007], Fresh[1006], Fresh[1005]}), .c ({signal_2025, signal_2024, signal_1277}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1263 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1865, signal_1864, signal_1198}), .a ({signal_1863, signal_1862, signal_1197}), .clk ( clk ), .r ({Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({signal_2027, signal_2026, signal_1278}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1264 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1869, signal_1868, signal_1200}), .a ({signal_1867, signal_1866, signal_1199}), .clk ( clk ), .r ({Fresh[1013], Fresh[1012], Fresh[1011]}), .c ({signal_2029, signal_2028, signal_1279}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1265 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1873, signal_1872, signal_1202}), .a ({signal_1871, signal_1870, signal_1201}), .clk ( clk ), .r ({Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({signal_2031, signal_2030, signal_1280}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1266 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1877, signal_1876, signal_1204}), .a ({signal_1875, signal_1874, signal_1203}), .clk ( clk ), .r ({Fresh[1019], Fresh[1018], Fresh[1017]}), .c ({signal_2033, signal_2032, signal_1281}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1267 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1881, signal_1880, signal_1206}), .a ({signal_1879, signal_1878, signal_1205}), .clk ( clk ), .r ({Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_2035, signal_2034, signal_1282}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1268 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1885, signal_1884, signal_1208}), .a ({signal_1883, signal_1882, signal_1207}), .clk ( clk ), .r ({Fresh[1025], Fresh[1024], Fresh[1023]}), .c ({signal_2037, signal_2036, signal_1283}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1269 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1889, signal_1888, signal_1210}), .a ({signal_1887, signal_1886, signal_1209}), .clk ( clk ), .r ({Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({signal_2039, signal_2038, signal_1284}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1270 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1893, signal_1892, signal_1212}), .a ({signal_1891, signal_1890, signal_1211}), .clk ( clk ), .r ({Fresh[1031], Fresh[1030], Fresh[1029]}), .c ({signal_2041, signal_2040, signal_1285}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1271 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1897, signal_1896, signal_1214}), .a ({signal_1895, signal_1894, signal_1213}), .clk ( clk ), .r ({Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({signal_2043, signal_2042, signal_1286}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1272 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1901, signal_1900, signal_1216}), .a ({signal_1899, signal_1898, signal_1215}), .clk ( clk ), .r ({Fresh[1037], Fresh[1036], Fresh[1035]}), .c ({signal_2045, signal_2044, signal_1287}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1273 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1905, signal_1904, signal_1218}), .a ({signal_1903, signal_1902, signal_1217}), .clk ( clk ), .r ({Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({signal_2047, signal_2046, signal_1288}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1274 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1909, signal_1908, signal_1220}), .a ({signal_1907, signal_1906, signal_1219}), .clk ( clk ), .r ({Fresh[1043], Fresh[1042], Fresh[1041]}), .c ({signal_2049, signal_2048, signal_1289}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1275 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1913, signal_1912, signal_1222}), .a ({signal_1911, signal_1910, signal_1221}), .clk ( clk ), .r ({Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({signal_2051, signal_2050, signal_1290}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1276 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1917, signal_1916, signal_1224}), .a ({signal_1915, signal_1914, signal_1223}), .clk ( clk ), .r ({Fresh[1049], Fresh[1048], Fresh[1047]}), .c ({signal_2053, signal_2052, signal_1291}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1277 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1921, signal_1920, signal_1226}), .a ({signal_1919, signal_1918, signal_1225}), .clk ( clk ), .r ({Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_2055, signal_2054, signal_1292}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1278 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1925, signal_1924, signal_1228}), .a ({signal_1923, signal_1922, signal_1227}), .clk ( clk ), .r ({Fresh[1055], Fresh[1054], Fresh[1053]}), .c ({signal_2057, signal_2056, signal_1293}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1279 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1927, signal_1926, signal_1229}), .a ({signal_3647, signal_3645, signal_3643}), .clk ( clk ), .r ({Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({signal_2059, signal_2058, signal_1294}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1280 ( .s ({signal_3641, signal_3633, signal_3625}), .b ({signal_1931, signal_1930, signal_1231}), .a ({signal_1929, signal_1928, signal_1230}), .clk ( clk ), .r ({Fresh[1061], Fresh[1060], Fresh[1059]}), .c ({signal_2061, signal_2060, signal_1295}) ) ;
    buf_clk cell_1568 ( .C ( clk ), .D ( signal_3656 ), .Q ( signal_3657 ) ) ;
    buf_clk cell_1578 ( .C ( clk ), .D ( signal_3666 ), .Q ( signal_3667 ) ) ;
    buf_clk cell_1588 ( .C ( clk ), .D ( signal_3676 ), .Q ( signal_3677 ) ) ;
    buf_clk cell_1598 ( .C ( clk ), .D ( signal_3686 ), .Q ( signal_3687 ) ) ;
    buf_clk cell_1610 ( .C ( clk ), .D ( signal_3698 ), .Q ( signal_3699 ) ) ;
    buf_clk cell_1622 ( .C ( clk ), .D ( signal_3710 ), .Q ( signal_3711 ) ) ;
    buf_clk cell_1634 ( .C ( clk ), .D ( signal_3722 ), .Q ( signal_3723 ) ) ;
    buf_clk cell_1648 ( .C ( clk ), .D ( signal_3736 ), .Q ( signal_3737 ) ) ;
    buf_clk cell_1662 ( .C ( clk ), .D ( signal_3750 ), .Q ( signal_3751 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_1599 ( .C ( clk ), .D ( signal_3687 ), .Q ( signal_3688 ) ) ;
    buf_clk cell_1611 ( .C ( clk ), .D ( signal_3699 ), .Q ( signal_3700 ) ) ;
    buf_clk cell_1623 ( .C ( clk ), .D ( signal_3711 ), .Q ( signal_3712 ) ) ;
    buf_clk cell_1635 ( .C ( clk ), .D ( signal_3723 ), .Q ( signal_3724 ) ) ;
    buf_clk cell_1649 ( .C ( clk ), .D ( signal_3737 ), .Q ( signal_3738 ) ) ;
    buf_clk cell_1663 ( .C ( clk ), .D ( signal_3751 ), .Q ( signal_3752 ) ) ;

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1281 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1937, signal_1936, signal_1233}), .a ({signal_1935, signal_1934, signal_1232}), .clk ( clk ), .r ({Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({signal_2065, signal_2064, signal_1296}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1282 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1941, signal_1940, signal_1235}), .a ({signal_1939, signal_1938, signal_1234}), .clk ( clk ), .r ({Fresh[1067], Fresh[1066], Fresh[1065]}), .c ({signal_2067, signal_2066, signal_1297}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1283 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1945, signal_1944, signal_1237}), .a ({signal_1943, signal_1942, signal_1236}), .clk ( clk ), .r ({Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({signal_2069, signal_2068, signal_1298}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1284 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1949, signal_1948, signal_1239}), .a ({signal_1947, signal_1946, signal_1238}), .clk ( clk ), .r ({Fresh[1073], Fresh[1072], Fresh[1071]}), .c ({signal_2071, signal_2070, signal_1299}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1285 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1953, signal_1952, signal_1241}), .a ({signal_1951, signal_1950, signal_1240}), .clk ( clk ), .r ({Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({signal_2073, signal_2072, signal_1300}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1286 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1957, signal_1956, signal_1243}), .a ({signal_1955, signal_1954, signal_1242}), .clk ( clk ), .r ({Fresh[1079], Fresh[1078], Fresh[1077]}), .c ({signal_2075, signal_2074, signal_1301}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1287 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1961, signal_1960, signal_1245}), .a ({signal_1959, signal_1958, signal_1244}), .clk ( clk ), .r ({Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_2077, signal_2076, signal_1302}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1288 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1965, signal_1964, signal_1247}), .a ({signal_1963, signal_1962, signal_1246}), .clk ( clk ), .r ({Fresh[1085], Fresh[1084], Fresh[1083]}), .c ({signal_2079, signal_2078, signal_1303}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1289 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1969, signal_1968, signal_1249}), .a ({signal_1967, signal_1966, signal_1248}), .clk ( clk ), .r ({Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({signal_2081, signal_2080, signal_1304}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1290 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1973, signal_1972, signal_1251}), .a ({signal_1971, signal_1970, signal_1250}), .clk ( clk ), .r ({Fresh[1091], Fresh[1090], Fresh[1089]}), .c ({signal_2083, signal_2082, signal_1305}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1291 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1977, signal_1976, signal_1253}), .a ({signal_1975, signal_1974, signal_1252}), .clk ( clk ), .r ({Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({signal_2085, signal_2084, signal_1306}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1292 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1981, signal_1980, signal_1255}), .a ({signal_1979, signal_1978, signal_1254}), .clk ( clk ), .r ({Fresh[1097], Fresh[1096], Fresh[1095]}), .c ({signal_2087, signal_2086, signal_1307}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1293 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1985, signal_1984, signal_1257}), .a ({signal_1983, signal_1982, signal_1256}), .clk ( clk ), .r ({Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({signal_2089, signal_2088, signal_1308}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1294 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1989, signal_1988, signal_1259}), .a ({signal_1987, signal_1986, signal_1258}), .clk ( clk ), .r ({Fresh[1103], Fresh[1102], Fresh[1101]}), .c ({signal_2091, signal_2090, signal_1309}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1295 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1993, signal_1992, signal_1261}), .a ({signal_1991, signal_1990, signal_1260}), .clk ( clk ), .r ({Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({signal_2093, signal_2092, signal_1310}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1296 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_1997, signal_1996, signal_1263}), .a ({signal_1995, signal_1994, signal_1262}), .clk ( clk ), .r ({Fresh[1109], Fresh[1108], Fresh[1107]}), .c ({signal_2095, signal_2094, signal_1311}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1297 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2001, signal_2000, signal_1265}), .a ({signal_1999, signal_1998, signal_1264}), .clk ( clk ), .r ({Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_2097, signal_2096, signal_1312}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1298 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2005, signal_2004, signal_1267}), .a ({signal_2003, signal_2002, signal_1266}), .clk ( clk ), .r ({Fresh[1115], Fresh[1114], Fresh[1113]}), .c ({signal_2099, signal_2098, signal_1313}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1299 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2009, signal_2008, signal_1269}), .a ({signal_2007, signal_2006, signal_1268}), .clk ( clk ), .r ({Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({signal_2101, signal_2100, signal_1314}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1300 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2013, signal_2012, signal_1271}), .a ({signal_2011, signal_2010, signal_1270}), .clk ( clk ), .r ({Fresh[1121], Fresh[1120], Fresh[1119]}), .c ({signal_2103, signal_2102, signal_1315}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1301 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2017, signal_2016, signal_1273}), .a ({signal_2015, signal_2014, signal_1272}), .clk ( clk ), .r ({Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({signal_2105, signal_2104, signal_1316}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1302 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2021, signal_2020, signal_1275}), .a ({signal_2019, signal_2018, signal_1274}), .clk ( clk ), .r ({Fresh[1127], Fresh[1126], Fresh[1125]}), .c ({signal_2107, signal_2106, signal_1317}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1303 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2025, signal_2024, signal_1277}), .a ({signal_2023, signal_2022, signal_1276}), .clk ( clk ), .r ({Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({signal_2109, signal_2108, signal_1318}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1304 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2029, signal_2028, signal_1279}), .a ({signal_2027, signal_2026, signal_1278}), .clk ( clk ), .r ({Fresh[1133], Fresh[1132], Fresh[1131]}), .c ({signal_2111, signal_2110, signal_1319}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1305 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2033, signal_2032, signal_1281}), .a ({signal_2031, signal_2030, signal_1280}), .clk ( clk ), .r ({Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({signal_2113, signal_2112, signal_1320}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1306 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2037, signal_2036, signal_1283}), .a ({signal_2035, signal_2034, signal_1282}), .clk ( clk ), .r ({Fresh[1139], Fresh[1138], Fresh[1137]}), .c ({signal_2115, signal_2114, signal_1321}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1307 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2041, signal_2040, signal_1285}), .a ({signal_2039, signal_2038, signal_1284}), .clk ( clk ), .r ({Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_2117, signal_2116, signal_1322}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1308 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2045, signal_2044, signal_1287}), .a ({signal_2043, signal_2042, signal_1286}), .clk ( clk ), .r ({Fresh[1145], Fresh[1144], Fresh[1143]}), .c ({signal_2119, signal_2118, signal_1323}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1309 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2049, signal_2048, signal_1289}), .a ({signal_2047, signal_2046, signal_1288}), .clk ( clk ), .r ({Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({signal_2121, signal_2120, signal_1324}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1310 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2053, signal_2052, signal_1291}), .a ({signal_2051, signal_2050, signal_1290}), .clk ( clk ), .r ({Fresh[1151], Fresh[1150], Fresh[1149]}), .c ({signal_2123, signal_2122, signal_1325}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1311 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2057, signal_2056, signal_1293}), .a ({signal_2055, signal_2054, signal_1292}), .clk ( clk ), .r ({Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({signal_2125, signal_2124, signal_1326}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1312 ( .s ({signal_3677, signal_3667, signal_3657}), .b ({signal_2061, signal_2060, signal_1295}), .a ({signal_2059, signal_2058, signal_1294}), .clk ( clk ), .r ({Fresh[1157], Fresh[1156], Fresh[1155]}), .c ({signal_2127, signal_2126, signal_1327}) ) ;
    buf_clk cell_1600 ( .C ( clk ), .D ( signal_3688 ), .Q ( signal_3689 ) ) ;
    buf_clk cell_1612 ( .C ( clk ), .D ( signal_3700 ), .Q ( signal_3701 ) ) ;
    buf_clk cell_1624 ( .C ( clk ), .D ( signal_3712 ), .Q ( signal_3713 ) ) ;
    buf_clk cell_1636 ( .C ( clk ), .D ( signal_3724 ), .Q ( signal_3725 ) ) ;
    buf_clk cell_1650 ( .C ( clk ), .D ( signal_3738 ), .Q ( signal_3739 ) ) ;
    buf_clk cell_1664 ( .C ( clk ), .D ( signal_3752 ), .Q ( signal_3753 ) ) ;

    /* cells in depth 13 */
    buf_clk cell_1637 ( .C ( clk ), .D ( signal_3725 ), .Q ( signal_3726 ) ) ;
    buf_clk cell_1651 ( .C ( clk ), .D ( signal_3739 ), .Q ( signal_3740 ) ) ;
    buf_clk cell_1665 ( .C ( clk ), .D ( signal_3753 ), .Q ( signal_3754 ) ) ;

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1313 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2067, signal_2066, signal_1297}), .a ({signal_2065, signal_2064, signal_1296}), .clk ( clk ), .r ({Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({signal_2131, signal_2130, signal_1328}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1314 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2071, signal_2070, signal_1299}), .a ({signal_2069, signal_2068, signal_1298}), .clk ( clk ), .r ({Fresh[1163], Fresh[1162], Fresh[1161]}), .c ({signal_2133, signal_2132, signal_1329}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1315 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2075, signal_2074, signal_1301}), .a ({signal_2073, signal_2072, signal_1300}), .clk ( clk ), .r ({Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({signal_2135, signal_2134, signal_1330}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1316 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2079, signal_2078, signal_1303}), .a ({signal_2077, signal_2076, signal_1302}), .clk ( clk ), .r ({Fresh[1169], Fresh[1168], Fresh[1167]}), .c ({signal_2137, signal_2136, signal_1331}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1317 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2083, signal_2082, signal_1305}), .a ({signal_2081, signal_2080, signal_1304}), .clk ( clk ), .r ({Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_2139, signal_2138, signal_1332}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1318 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2087, signal_2086, signal_1307}), .a ({signal_2085, signal_2084, signal_1306}), .clk ( clk ), .r ({Fresh[1175], Fresh[1174], Fresh[1173]}), .c ({signal_2141, signal_2140, signal_1333}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1319 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2091, signal_2090, signal_1309}), .a ({signal_2089, signal_2088, signal_1308}), .clk ( clk ), .r ({Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({signal_2143, signal_2142, signal_1334}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1320 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2095, signal_2094, signal_1311}), .a ({signal_2093, signal_2092, signal_1310}), .clk ( clk ), .r ({Fresh[1181], Fresh[1180], Fresh[1179]}), .c ({signal_2145, signal_2144, signal_1335}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1321 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2099, signal_2098, signal_1313}), .a ({signal_2097, signal_2096, signal_1312}), .clk ( clk ), .r ({Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({signal_2147, signal_2146, signal_1336}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1322 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2103, signal_2102, signal_1315}), .a ({signal_2101, signal_2100, signal_1314}), .clk ( clk ), .r ({Fresh[1187], Fresh[1186], Fresh[1185]}), .c ({signal_2149, signal_2148, signal_1337}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1323 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2107, signal_2106, signal_1317}), .a ({signal_2105, signal_2104, signal_1316}), .clk ( clk ), .r ({Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({signal_2151, signal_2150, signal_1338}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1324 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2111, signal_2110, signal_1319}), .a ({signal_2109, signal_2108, signal_1318}), .clk ( clk ), .r ({Fresh[1193], Fresh[1192], Fresh[1191]}), .c ({signal_2153, signal_2152, signal_1339}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1325 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2115, signal_2114, signal_1321}), .a ({signal_2113, signal_2112, signal_1320}), .clk ( clk ), .r ({Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({signal_2155, signal_2154, signal_1340}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1326 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2119, signal_2118, signal_1323}), .a ({signal_2117, signal_2116, signal_1322}), .clk ( clk ), .r ({Fresh[1199], Fresh[1198], Fresh[1197]}), .c ({signal_2157, signal_2156, signal_1341}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1327 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2123, signal_2122, signal_1325}), .a ({signal_2121, signal_2120, signal_1324}), .clk ( clk ), .r ({Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_2159, signal_2158, signal_1342}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1328 ( .s ({signal_3713, signal_3701, signal_3689}), .b ({signal_2127, signal_2126, signal_1327}), .a ({signal_2125, signal_2124, signal_1326}), .clk ( clk ), .r ({Fresh[1205], Fresh[1204], Fresh[1203]}), .c ({signal_2161, signal_2160, signal_1343}) ) ;
    buf_clk cell_1638 ( .C ( clk ), .D ( signal_3726 ), .Q ( signal_3727 ) ) ;
    buf_clk cell_1652 ( .C ( clk ), .D ( signal_3740 ), .Q ( signal_3741 ) ) ;
    buf_clk cell_1666 ( .C ( clk ), .D ( signal_3754 ), .Q ( signal_3755 ) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1329 ( .s ({signal_3755, signal_3741, signal_3727}), .b ({signal_2133, signal_2132, signal_1329}), .a ({signal_2131, signal_2130, signal_1328}), .clk ( clk ), .r ({Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({signal_2165, signal_2164, signal_30}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1330 ( .s ({signal_3755, signal_3741, signal_3727}), .b ({signal_2137, signal_2136, signal_1331}), .a ({signal_2135, signal_2134, signal_1330}), .clk ( clk ), .r ({Fresh[1211], Fresh[1210], Fresh[1209]}), .c ({signal_2167, signal_2166, signal_29}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1331 ( .s ({signal_3755, signal_3741, signal_3727}), .b ({signal_2141, signal_2140, signal_1333}), .a ({signal_2139, signal_2138, signal_1332}), .clk ( clk ), .r ({Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({signal_2169, signal_2168, signal_28}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1332 ( .s ({signal_3755, signal_3741, signal_3727}), .b ({signal_2145, signal_2144, signal_1335}), .a ({signal_2143, signal_2142, signal_1334}), .clk ( clk ), .r ({Fresh[1217], Fresh[1216], Fresh[1215]}), .c ({signal_2171, signal_2170, signal_27}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1333 ( .s ({signal_3755, signal_3741, signal_3727}), .b ({signal_2149, signal_2148, signal_1337}), .a ({signal_2147, signal_2146, signal_1336}), .clk ( clk ), .r ({Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({signal_2173, signal_2172, signal_26}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1334 ( .s ({signal_3755, signal_3741, signal_3727}), .b ({signal_2153, signal_2152, signal_1339}), .a ({signal_2151, signal_2150, signal_1338}), .clk ( clk ), .r ({Fresh[1223], Fresh[1222], Fresh[1221]}), .c ({signal_2175, signal_2174, signal_25}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1335 ( .s ({signal_3755, signal_3741, signal_3727}), .b ({signal_2157, signal_2156, signal_1341}), .a ({signal_2155, signal_2154, signal_1340}), .clk ( clk ), .r ({Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({signal_2177, signal_2176, signal_24}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) cell_1336 ( .s ({signal_3755, signal_3741, signal_3727}), .b ({signal_2161, signal_2160, signal_1343}), .a ({signal_2159, signal_2158, signal_1342}), .clk ( clk ), .r ({Fresh[1229], Fresh[1228], Fresh[1227]}), .c ({signal_2179, signal_2178, signal_23}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_2179, signal_2178, signal_23}), .Q ({SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_2177, signal_2176, signal_24}), .Q ({SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_2175, signal_2174, signal_25}), .Q ({SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_2173, signal_2172, signal_26}), .Q ({SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_4 ( .clk ( clk ), .D ({signal_2171, signal_2170, signal_27}), .Q ({SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_5 ( .clk ( clk ), .D ({signal_2169, signal_2168, signal_28}), .Q ({SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_6 ( .clk ( clk ), .D ({signal_2167, signal_2166, signal_29}), .Q ({SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_7 ( .clk ( clk ), .D ({signal_2165, signal_2164, signal_30}), .Q ({SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
