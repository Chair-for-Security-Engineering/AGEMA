/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 16 time(s)  */

module sbox_HPC2_BDDsylvan_ClockGating_d2 (X_s0, clk, X_s1, X_s2, Fresh, rst, Y_s0, Y_s1, Y_s2, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input rst ;
    input [1229:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output Synch ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_2636 ;

    /* cells in depth 0 */
    ClockGatingController #(17) cell_546 ( .clk (clk), .rst (rst), .GatedClk (signal_2636), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_136 ( .s ({X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_556, signal_555, signal_151}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_137 ( .s ({X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({signal_558, signal_557, signal_152}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_138 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_562, signal_561, signal_153}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_139 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({signal_564, signal_563, signal_154}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_140 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_568, signal_567, signal_155}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_141 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({signal_570, signal_569, signal_156}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_142 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_556, signal_555, signal_151}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_572, signal_571, signal_157}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_143 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_558, signal_557, signal_152}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({signal_574, signal_573, signal_158}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_144 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_556, signal_555, signal_151}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_576, signal_575, signal_159}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_145 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_556, signal_555, signal_151}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({signal_578, signal_577, signal_160}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_146 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_558, signal_557, signal_152}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_580, signal_579, signal_161}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_147 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_558, signal_557, signal_152}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({signal_582, signal_581, signal_162}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_148 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_584, signal_583, signal_163}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_149 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({signal_586, signal_585, signal_164}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_150 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_564, signal_563, signal_154}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_588, signal_587, signal_165}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_151 ( .s ({X_s2[1], X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({signal_590, signal_589, signal_166}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_152 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_558, signal_557, signal_152}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_592, signal_591, signal_167}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_153 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_562, signal_561, signal_153}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({signal_594, signal_593, signal_168}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_154 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_562, signal_561, signal_153}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_596, signal_595, signal_169}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_155 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_564, signal_563, signal_154}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({signal_598, signal_597, signal_170}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_156 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_564, signal_563, signal_154}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_600, signal_599, signal_171}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_157 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_564, signal_563, signal_154}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({signal_602, signal_601, signal_172}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_158 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_562, signal_561, signal_153}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_604, signal_603, signal_173}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_159 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_562, signal_561, signal_153}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({signal_606, signal_605, signal_174}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_160 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_608, signal_607, signal_175}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_161 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_558, signal_557, signal_152}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({signal_610, signal_609, signal_176}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_162 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_564, signal_563, signal_154}), .a ({signal_562, signal_561, signal_153}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_612, signal_611, signal_177}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_163 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_558, signal_557, signal_152}), .a ({signal_564, signal_563, signal_154}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({signal_614, signal_613, signal_178}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_164 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_562, signal_561, signal_153}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_616, signal_615, signal_179}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_165 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_564, signal_563, signal_154}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({signal_618, signal_617, signal_180}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_166 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_570, signal_569, signal_156}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_620, signal_619, signal_181}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_167 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_574, signal_573, signal_158}), .a ({signal_572, signal_571, signal_157}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({signal_622, signal_621, signal_182}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_168 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_576, signal_575, signal_159}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_624, signal_623, signal_183}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_169 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_578, signal_577, signal_160}), .a ({signal_562, signal_561, signal_153}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({signal_626, signal_625, signal_184}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_170 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_628, signal_627, signal_185}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_171 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_582, signal_581, signal_162}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({signal_630, signal_629, signal_186}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_172 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_558, signal_557, signal_152}), .a ({signal_584, signal_583, signal_163}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_632, signal_631, signal_187}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_173 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({signal_634, signal_633, signal_188}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_174 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_572, signal_571, signal_157}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_636, signal_635, signal_189}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_175 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_576, signal_575, signal_159}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({signal_638, signal_637, signal_190}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_176 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_582, signal_581, signal_162}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_640, signal_639, signal_191}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_177 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_161}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({signal_642, signal_641, signal_192}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_178 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_558, signal_557, signal_152}), .a ({signal_574, signal_573, signal_158}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_644, signal_643, signal_193}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_179 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_556, signal_555, signal_151}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({signal_646, signal_645, signal_194}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_180 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_648, signal_647, signal_195}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_181 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_586, signal_585, signal_164}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({signal_650, signal_649, signal_196}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_182 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_586, signal_585, signal_164}), .a ({signal_570, signal_569, signal_156}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_652, signal_651, signal_197}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_183 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_558, signal_557, signal_152}), .a ({signal_590, signal_589, signal_166}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({signal_654, signal_653, signal_198}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_184 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_586, signal_585, signal_164}), .a ({signal_564, signal_563, signal_154}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_656, signal_655, signal_199}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_185 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_562, signal_561, signal_153}), .a ({signal_572, signal_571, signal_157}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({signal_658, signal_657, signal_200}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_186 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_572, signal_571, signal_157}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_660, signal_659, signal_201}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_187 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_574, signal_573, signal_158}), .a ({signal_570, signal_569, signal_156}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({signal_662, signal_661, signal_202}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_188 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_574, signal_573, signal_158}), .a ({signal_576, signal_575, signal_159}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_664, signal_663, signal_203}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_189 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_584, signal_583, signal_163}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({signal_666, signal_665, signal_204}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_190 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_578, signal_577, signal_160}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_668, signal_667, signal_205}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_191 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_564, signal_563, signal_154}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({signal_670, signal_669, signal_206}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_192 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_574, signal_573, signal_158}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_672, signal_671, signal_207}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_193 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_576, signal_575, signal_159}), .a ({signal_574, signal_573, signal_158}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({signal_674, signal_673, signal_208}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_194 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({signal_564, signal_563, signal_154}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_676, signal_675, signal_209}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_195 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_584, signal_583, signal_163}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({signal_678, signal_677, signal_210}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_196 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_584, signal_583, signal_163}), .a ({signal_578, signal_577, signal_160}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_680, signal_679, signal_211}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_197 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_570, signal_569, signal_156}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({signal_682, signal_681, signal_212}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_198 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_578, signal_577, signal_160}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_684, signal_683, signal_213}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_199 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({signal_576, signal_575, signal_159}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({signal_686, signal_685, signal_214}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_200 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_578, signal_577, signal_160}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_688, signal_687, signal_215}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_201 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_558, signal_557, signal_152}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({signal_690, signal_689, signal_216}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_202 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_556, signal_555, signal_151}), .a ({signal_570, signal_569, signal_156}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_692, signal_691, signal_217}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_203 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_586, signal_585, signal_164}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({signal_694, signal_693, signal_218}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_204 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_574, signal_573, signal_158}), .a ({signal_582, signal_581, signal_162}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({signal_696, signal_695, signal_219}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_205 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_562, signal_561, signal_153}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({signal_698, signal_697, signal_220}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_206 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_161}), .a ({signal_590, signal_589, signal_166}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_700, signal_699, signal_221}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_207 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({signal_702, signal_701, signal_222}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_208 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_161}), .a ({signal_574, signal_573, signal_158}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({signal_704, signal_703, signal_223}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_209 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_558, signal_557, signal_152}), .a ({signal_572, signal_571, signal_157}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({signal_706, signal_705, signal_224}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_210 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_564, signal_563, signal_154}), .a ({signal_570, signal_569, signal_156}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({signal_708, signal_707, signal_225}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_211 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_574, signal_573, signal_158}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({signal_710, signal_709, signal_226}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_212 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_572, signal_571, signal_157}), .a ({signal_590, signal_589, signal_166}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({signal_712, signal_711, signal_227}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_213 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_586, signal_585, signal_164}), .a ({signal_584, signal_583, signal_163}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({signal_714, signal_713, signal_228}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_214 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_574, signal_573, signal_158}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({signal_716, signal_715, signal_229}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_215 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_576, signal_575, signal_159}), .a ({signal_584, signal_583, signal_163}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({signal_718, signal_717, signal_230}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_216 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_161}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_720, signal_719, signal_231}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_217 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_161}), .a ({signal_576, signal_575, signal_159}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({signal_722, signal_721, signal_232}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_218 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_574, signal_573, signal_158}), .a ({signal_564, signal_563, signal_154}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({signal_724, signal_723, signal_233}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_219 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_584, signal_583, signal_163}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({signal_726, signal_725, signal_234}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_220 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({signal_728, signal_727, signal_235}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_221 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_574, signal_573, signal_158}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({signal_730, signal_729, signal_236}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_222 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_586, signal_585, signal_164}), .a ({signal_562, signal_561, signal_153}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({signal_732, signal_731, signal_237}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_223 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_586, signal_585, signal_164}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({signal_734, signal_733, signal_238}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_224 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_562, signal_561, signal_153}), .a ({signal_582, signal_581, signal_162}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({signal_736, signal_735, signal_239}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_225 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({signal_738, signal_737, signal_240}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_226 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_578, signal_577, signal_160}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_740, signal_739, signal_241}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_227 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_582, signal_581, signal_162}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({signal_742, signal_741, signal_242}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_228 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({signal_744, signal_743, signal_243}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_229 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({signal_582, signal_581, signal_162}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({signal_746, signal_745, signal_244}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_230 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_564, signal_563, signal_154}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({signal_748, signal_747, signal_245}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_231 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_572, signal_571, signal_157}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({signal_750, signal_749, signal_246}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_232 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_562, signal_561, signal_153}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({signal_752, signal_751, signal_247}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_233 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_584, signal_583, signal_163}), .a ({signal_590, signal_589, signal_166}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({signal_754, signal_753, signal_248}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_234 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({signal_570, signal_569, signal_156}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({signal_756, signal_755, signal_249}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_235 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_161}), .a ({signal_564, signal_563, signal_154}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({signal_758, signal_757, signal_250}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_236 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_576, signal_575, signal_159}), .a ({signal_578, signal_577, signal_160}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_760, signal_759, signal_251}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_237 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_586, signal_585, signal_164}), .a ({signal_576, signal_575, signal_159}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({signal_762, signal_761, signal_252}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_238 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_161}), .a ({signal_584, signal_583, signal_163}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({signal_764, signal_763, signal_253}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_239 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_582, signal_581, signal_162}), .a ({signal_578, signal_577, signal_160}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({signal_766, signal_765, signal_254}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_240 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_586, signal_585, signal_164}), .a ({signal_572, signal_571, signal_157}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({signal_768, signal_767, signal_255}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_241 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_578, signal_577, signal_160}), .a ({signal_574, signal_573, signal_158}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({signal_770, signal_769, signal_256}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_242 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_558, signal_557, signal_152}), .a ({signal_576, signal_575, signal_159}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({signal_772, signal_771, signal_257}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_243 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_590, signal_589, signal_166}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({signal_774, signal_773, signal_258}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_244 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_564, signal_563, signal_154}), .a ({signal_578, signal_577, signal_160}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({signal_776, signal_775, signal_259}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_245 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_161}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({signal_778, signal_777, signal_260}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_246 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_556, signal_555, signal_151}), .a ({signal_582, signal_581, signal_162}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_780, signal_779, signal_261}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_247 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_582, signal_581, signal_162}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({signal_782, signal_781, signal_262}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_248 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_578, signal_577, signal_160}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({signal_784, signal_783, signal_263}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_249 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_582, signal_581, signal_162}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({signal_786, signal_785, signal_264}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_250 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_578, signal_577, signal_160}), .a ({signal_572, signal_571, signal_157}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({signal_788, signal_787, signal_265}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_251 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_576, signal_575, signal_159}), .a ({signal_562, signal_561, signal_153}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({signal_790, signal_789, signal_266}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_252 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({signal_792, signal_791, signal_267}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_253 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_582, signal_581, signal_162}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({signal_794, signal_793, signal_268}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_254 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_584, signal_583, signal_163}), .a ({signal_570, signal_569, signal_156}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({signal_796, signal_795, signal_269}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_255 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_161}), .a ({signal_582, signal_581, signal_162}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({signal_798, signal_797, signal_270}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_256 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_564, signal_563, signal_154}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_800, signal_799, signal_271}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_257 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_564, signal_563, signal_154}), .a ({signal_574, signal_573, signal_158}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({signal_802, signal_801, signal_272}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_258 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_584, signal_583, signal_163}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({signal_804, signal_803, signal_273}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_259 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_572, signal_571, signal_157}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({signal_806, signal_805, signal_274}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_260 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_578, signal_577, signal_160}), .a ({signal_570, signal_569, signal_156}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({signal_808, signal_807, signal_275}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_261 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_562, signal_561, signal_153}), .a ({signal_574, signal_573, signal_158}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({signal_810, signal_809, signal_276}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_262 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_582, signal_581, signal_162}), .a ({signal_564, signal_563, signal_154}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({signal_812, signal_811, signal_277}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_263 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({signal_814, signal_813, signal_278}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_264 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_578, signal_577, signal_160}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({signal_816, signal_815, signal_279}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_265 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({signal_818, signal_817, signal_280}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_266 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_820, signal_819, signal_281}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_267 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_576, signal_575, signal_159}), .a ({signal_590, signal_589, signal_166}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({signal_822, signal_821, signal_282}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_268 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_572, signal_571, signal_157}), .a ({signal_562, signal_561, signal_153}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({signal_824, signal_823, signal_283}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_269 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_574, signal_573, signal_158}), .a ({signal_578, signal_577, signal_160}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({signal_826, signal_825, signal_284}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_270 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({signal_828, signal_827, signal_285}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_271 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_586, signal_585, signal_164}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({signal_830, signal_829, signal_286}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_272 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_576, signal_575, signal_159}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({signal_832, signal_831, signal_287}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_273 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({signal_584, signal_583, signal_163}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({signal_834, signal_833, signal_288}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_274 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({signal_836, signal_835, signal_289}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_275 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_576, signal_575, signal_159}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({signal_838, signal_837, signal_290}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_276 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_590, signal_589, signal_166}), .a ({signal_578, signal_577, signal_160}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_840, signal_839, signal_291}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_277 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_584, signal_583, signal_163}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({signal_842, signal_841, signal_292}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_278 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_572, signal_571, signal_157}), .a ({signal_582, signal_581, signal_162}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({signal_844, signal_843, signal_293}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_279 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_578, signal_577, signal_160}), .a ({signal_556, signal_555, signal_151}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({signal_846, signal_845, signal_294}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_280 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_584, signal_583, signal_163}), .a ({signal_572, signal_571, signal_157}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({signal_848, signal_847, signal_295}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_281 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_582, signal_581, signal_162}), .a ({signal_590, signal_589, signal_166}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({signal_850, signal_849, signal_296}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_282 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_572, signal_571, signal_157}), .a ({signal_578, signal_577, signal_160}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({signal_852, signal_851, signal_297}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_283 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_562, signal_561, signal_153}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({signal_854, signal_853, signal_298}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_284 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_574, signal_573, signal_158}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({signal_856, signal_855, signal_299}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_285 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_556, signal_555, signal_151}), .a ({signal_590, signal_589, signal_166}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({signal_858, signal_857, signal_300}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_286 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b0}), .a ({signal_580, signal_579, signal_161}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_860, signal_859, signal_301}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_287 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_576, signal_575, signal_159}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({signal_862, signal_861, signal_302}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_288 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_584, signal_583, signal_163}), .a ({signal_562, signal_561, signal_153}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({signal_864, signal_863, signal_303}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_289 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_584, signal_583, signal_163}), .a ({signal_574, signal_573, signal_158}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({signal_866, signal_865, signal_304}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_290 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_572, signal_571, signal_157}), .a ({signal_574, signal_573, signal_158}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({signal_868, signal_867, signal_305}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_291 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_572, signal_571, signal_157}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({signal_870, signal_869, signal_306}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_292 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_161}), .a ({signal_578, signal_577, signal_160}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({signal_872, signal_871, signal_307}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_293 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_578, signal_577, signal_160}), .a ({signal_582, signal_581, signal_162}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({signal_874, signal_873, signal_308}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_294 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_558, signal_557, signal_152}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({signal_876, signal_875, signal_309}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_295 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_590, signal_589, signal_166}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({signal_878, signal_877, signal_310}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_296 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_558, signal_557, signal_152}), .a ({signal_618, signal_617, signal_180}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_882, signal_881, signal_311}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_297 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_584, signal_583, signal_163}), .a ({signal_564, signal_563, signal_154}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({signal_884, signal_883, signal_312}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_298 ( .s ({X_s2[2], X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_586, signal_585, signal_164}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({signal_886, signal_885, signal_313}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_299 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_622, signal_621, signal_182}), .a ({signal_620, signal_619, signal_181}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({signal_888, signal_887, signal_314}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_300 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_626, signal_625, signal_184}), .a ({signal_624, signal_623, signal_183}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({signal_890, signal_889, signal_315}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_301 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_630, signal_629, signal_186}), .a ({signal_628, signal_627, signal_185}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({signal_892, signal_891, signal_316}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_302 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_634, signal_633, signal_188}), .a ({signal_632, signal_631, signal_187}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({signal_894, signal_893, signal_317}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_303 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_638, signal_637, signal_190}), .a ({signal_636, signal_635, signal_189}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({signal_896, signal_895, signal_318}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_304 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_636, signal_635, signal_189}), .a ({signal_640, signal_639, signal_191}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({signal_898, signal_897, signal_319}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_305 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_642, signal_641, signal_192}), .a ({signal_588, signal_587, signal_165}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({signal_900, signal_899, signal_320}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_306 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_646, signal_645, signal_194}), .a ({signal_644, signal_643, signal_193}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_902, signal_901, signal_321}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_307 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_650, signal_649, signal_196}), .a ({signal_648, signal_647, signal_195}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({signal_904, signal_903, signal_322}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_308 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_592, signal_591, signal_167}), .a ({signal_652, signal_651, signal_197}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({signal_906, signal_905, signal_323}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_309 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_656, signal_655, signal_199}), .a ({signal_654, signal_653, signal_198}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({signal_908, signal_907, signal_324}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_310 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_658, signal_657, signal_200}), .a ({signal_632, signal_631, signal_187}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({signal_910, signal_909, signal_325}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_311 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_662, signal_661, signal_202}), .a ({signal_660, signal_659, signal_201}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({signal_912, signal_911, signal_326}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_312 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_666, signal_665, signal_204}), .a ({signal_664, signal_663, signal_203}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({signal_914, signal_913, signal_327}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_313 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_670, signal_669, signal_206}), .a ({signal_668, signal_667, signal_205}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({signal_916, signal_915, signal_328}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_314 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_674, signal_673, signal_208}), .a ({signal_672, signal_671, signal_207}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({signal_918, signal_917, signal_329}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_315 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_678, signal_677, signal_210}), .a ({signal_676, signal_675, signal_209}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({signal_920, signal_919, signal_330}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_316 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_682, signal_681, signal_212}), .a ({signal_680, signal_679, signal_211}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_922, signal_921, signal_331}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_317 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_644, signal_643, signal_193}), .a ({signal_684, signal_683, signal_213}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({signal_924, signal_923, signal_332}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_318 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_688, signal_687, signal_215}), .a ({signal_686, signal_685, signal_214}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({signal_926, signal_925, signal_333}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_319 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_692, signal_691, signal_217}), .a ({signal_690, signal_689, signal_216}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({signal_928, signal_927, signal_334}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_320 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_696, signal_695, signal_219}), .a ({signal_694, signal_693, signal_218}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({signal_930, signal_929, signal_335}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_321 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_698, signal_697, signal_220}), .a ({signal_594, signal_593, signal_168}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({signal_932, signal_931, signal_336}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_322 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_702, signal_701, signal_222}), .a ({signal_700, signal_699, signal_221}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({signal_934, signal_933, signal_337}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_323 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_706, signal_705, signal_224}), .a ({signal_704, signal_703, signal_223}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({signal_936, signal_935, signal_338}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_324 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_710, signal_709, signal_226}), .a ({signal_708, signal_707, signal_225}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({signal_938, signal_937, signal_339}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_325 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_712, signal_711, signal_227}), .a ({signal_680, signal_679, signal_211}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({signal_940, signal_939, signal_340}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_326 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_632, signal_631, signal_187}), .a ({signal_628, signal_627, signal_185}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_942, signal_941, signal_341}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_327 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_716, signal_715, signal_229}), .a ({signal_714, signal_713, signal_228}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({signal_944, signal_943, signal_342}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_328 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_718, signal_717, signal_230}), .a ({1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({signal_946, signal_945, signal_343}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_329 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_596, signal_595, signal_169}), .a ({signal_708, signal_707, signal_225}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({signal_948, signal_947, signal_344}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_330 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_718, signal_717, signal_230}), .a ({signal_598, signal_597, signal_170}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({signal_950, signal_949, signal_345}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_331 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_626, signal_625, signal_184}), .a ({signal_600, signal_599, signal_171}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({signal_952, signal_951, signal_346}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_332 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_588, signal_587, signal_165}), .a ({signal_720, signal_719, signal_231}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({signal_954, signal_953, signal_347}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_333 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_724, signal_723, signal_233}), .a ({signal_722, signal_721, signal_232}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({signal_956, signal_955, signal_348}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_334 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_598, signal_597, signal_170}), .a ({signal_696, signal_695, signal_219}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({signal_958, signal_957, signal_349}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_335 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_718, signal_717, signal_230}), .a ({signal_726, signal_725, signal_234}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({signal_960, signal_959, signal_350}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_336 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_730, signal_729, signal_236}), .a ({signal_728, signal_727, signal_235}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_962, signal_961, signal_351}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_337 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_602, signal_601, signal_172}), .a ({signal_732, signal_731, signal_237}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({signal_964, signal_963, signal_352}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_338 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_734, signal_733, signal_238}), .a ({signal_604, signal_603, signal_173}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({signal_966, signal_965, signal_353}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_339 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_738, signal_737, signal_240}), .a ({signal_736, signal_735, signal_239}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({signal_968, signal_967, signal_354}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_340 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_742, signal_741, signal_242}), .a ({signal_740, signal_739, signal_241}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({signal_970, signal_969, signal_355}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_341 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_746, signal_745, signal_244}), .a ({signal_744, signal_743, signal_243}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({signal_972, signal_971, signal_356}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_342 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_630, signal_629, signal_186}), .a ({signal_748, signal_747, signal_245}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({signal_974, signal_973, signal_357}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_343 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_752, signal_751, signal_247}), .a ({signal_750, signal_749, signal_246}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({signal_976, signal_975, signal_358}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_344 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_734, signal_733, signal_238}), .a ({signal_754, signal_753, signal_248}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({signal_978, signal_977, signal_359}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_345 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_756, signal_755, signal_249}), .a ({signal_732, signal_731, signal_237}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({signal_980, signal_979, signal_360}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_346 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_758, signal_757, signal_250}), .a ({signal_702, signal_701, signal_222}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_982, signal_981, signal_361}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_347 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_760, signal_759, signal_251}), .a ({signal_662, signal_661, signal_202}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({signal_984, signal_983, signal_362}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_348 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_764, signal_763, signal_253}), .a ({signal_762, signal_761, signal_252}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({signal_986, signal_985, signal_363}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_349 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_766, signal_765, signal_254}), .a ({signal_676, signal_675, signal_209}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({signal_988, signal_987, signal_364}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_350 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_768, signal_767, signal_255}), .a ({signal_734, signal_733, signal_238}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({signal_990, signal_989, signal_365}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_351 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_772, signal_771, signal_257}), .a ({signal_770, signal_769, signal_256}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({signal_992, signal_991, signal_366}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_352 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_776, signal_775, signal_259}), .a ({signal_774, signal_773, signal_258}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({signal_994, signal_993, signal_367}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_353 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_600, signal_599, signal_171}), .a ({signal_778, signal_777, signal_260}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({signal_996, signal_995, signal_368}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_354 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_768, signal_767, signal_255}), .a ({signal_670, signal_669, signal_206}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({signal_998, signal_997, signal_369}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_355 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_648, signal_647, signal_195}), .a ({signal_780, signal_779, signal_261}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({signal_1000, signal_999, signal_370}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_356 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_696, signal_695, signal_219}), .a ({signal_644, signal_643, signal_193}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_1002, signal_1001, signal_371}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_357 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_738, signal_737, signal_240}), .a ({1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({signal_1004, signal_1003, signal_372}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_358 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_718, signal_717, signal_230}), .a ({signal_782, signal_781, signal_262}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({signal_1006, signal_1005, signal_373}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_359 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_784, signal_783, signal_263}), .a ({signal_636, signal_635, signal_189}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({signal_1008, signal_1007, signal_374}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_360 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_742, signal_741, signal_242}), .a ({signal_786, signal_785, signal_264}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({signal_1010, signal_1009, signal_375}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_361 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_790, signal_789, signal_266}), .a ({signal_788, signal_787, signal_265}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({signal_1012, signal_1011, signal_376}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_362 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_690, signal_689, signal_216}), .a ({signal_792, signal_791, signal_267}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({signal_1014, signal_1013, signal_377}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_363 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_636, signal_635, signal_189}), .a ({signal_794, signal_793, signal_268}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({signal_1016, signal_1015, signal_378}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_364 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_716, signal_715, signal_229}), .a ({signal_606, signal_605, signal_174}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({signal_1018, signal_1017, signal_379}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_365 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_796, signal_795, signal_269}), .a ({signal_724, signal_723, signal_233}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({signal_1020, signal_1019, signal_380}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_366 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_596, signal_595, signal_169}), .a ({signal_696, signal_695, signal_219}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_1022, signal_1021, signal_381}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_367 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_630, signal_629, signal_186}), .a ({signal_798, signal_797, signal_270}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({signal_1024, signal_1023, signal_382}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_368 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_700, signal_699, signal_221}), .a ({signal_640, signal_639, signal_191}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({signal_1026, signal_1025, signal_383}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_369 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_756, signal_755, signal_249}), .a ({signal_800, signal_799, signal_271}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({signal_1028, signal_1027, signal_384}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_370 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_702, signal_701, signal_222}), .a ({signal_802, signal_801, signal_272}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({signal_1030, signal_1029, signal_385}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_371 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_806, signal_805, signal_274}), .a ({signal_804, signal_803, signal_273}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({signal_1032, signal_1031, signal_386}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_372 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_808, signal_807, signal_275}), .a ({signal_632, signal_631, signal_187}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({signal_1034, signal_1033, signal_387}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_373 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_810, signal_809, signal_276}), .a ({signal_708, signal_707, signal_225}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({signal_1036, signal_1035, signal_388}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_374 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_792, signal_791, signal_267}), .a ({signal_568, signal_567, signal_155}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({signal_1038, signal_1037, signal_389}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_375 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_814, signal_813, signal_278}), .a ({signal_812, signal_811, signal_277}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({signal_1040, signal_1039, signal_390}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_376 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_584, signal_583, signal_163}), .a ({signal_816, signal_815, signal_279}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_1042, signal_1041, signal_391}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_377 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_818, signal_817, signal_280}), .a ({signal_782, signal_781, signal_262}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({signal_1044, signal_1043, signal_392}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_378 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_622, signal_621, signal_182}), .a ({signal_660, signal_659, signal_201}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({signal_1046, signal_1045, signal_393}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_379 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_640, signal_639, signal_191}), .a ({signal_820, signal_819, signal_281}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({signal_1048, signal_1047, signal_394}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_380 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_658, signal_657, signal_200}), .a ({signal_756, signal_755, signal_249}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({signal_1050, signal_1049, signal_395}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_381 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_620, signal_619, signal_181}), .a ({signal_694, signal_693, signal_218}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({signal_1052, signal_1051, signal_396}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_382 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_628, signal_627, signal_185}), .a ({signal_780, signal_779, signal_261}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({signal_1054, signal_1053, signal_397}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_383 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_822, signal_821, signal_282}), .a ({signal_718, signal_717, signal_230}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({signal_1056, signal_1055, signal_398}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_384 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_796, signal_795, signal_269}), .a ({signal_564, signal_563, signal_154}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({signal_1058, signal_1057, signal_399}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_385 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_824, signal_823, signal_283}), .a ({signal_642, signal_641, signal_192}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({signal_1060, signal_1059, signal_400}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_386 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_828, signal_827, signal_285}), .a ({signal_826, signal_825, signal_284}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_1062, signal_1061, signal_401}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_387 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_812, signal_811, signal_277}), .a ({signal_830, signal_829, signal_286}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({signal_1064, signal_1063, signal_402}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_388 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_662, signal_661, signal_202}), .a ({signal_558, signal_557, signal_152}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({signal_1066, signal_1065, signal_403}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_389 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_834, signal_833, signal_288}), .a ({signal_832, signal_831, signal_287}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({signal_1068, signal_1067, signal_404}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_390 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_744, signal_743, signal_243}), .a ({signal_632, signal_631, signal_187}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({signal_1070, signal_1069, signal_405}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_391 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_634, signal_633, signal_188}), .a ({signal_836, signal_835, signal_289}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({signal_1072, signal_1071, signal_406}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_392 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_714, signal_713, signal_228}), .a ({signal_608, signal_607, signal_175}), .clk (clk), .r ({Fresh[770], Fresh[769], Fresh[768]}), .c ({signal_1074, signal_1073, signal_407}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_393 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_840, signal_839, signal_291}), .a ({signal_838, signal_837, signal_290}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771]}), .c ({signal_1076, signal_1075, signal_408}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_394 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_842, signal_841, signal_292}), .a ({signal_576, signal_575, signal_159}), .clk (clk), .r ({Fresh[776], Fresh[775], Fresh[774]}), .c ({signal_1078, signal_1077, signal_409}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_395 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_730, signal_729, signal_236}), .a ({signal_844, signal_843, signal_293}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777]}), .c ({signal_1080, signal_1079, signal_410}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_396 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_562, signal_561, signal_153}), .a ({signal_818, signal_817, signal_280}), .clk (clk), .r ({Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_1082, signal_1081, signal_411}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_397 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_846, signal_845, signal_294}), .a ({signal_780, signal_779, signal_261}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783]}), .c ({signal_1084, signal_1083, signal_412}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_398 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_850, signal_849, signal_296}), .a ({signal_848, signal_847, signal_295}), .clk (clk), .r ({Fresh[788], Fresh[787], Fresh[786]}), .c ({signal_1086, signal_1085, signal_413}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_399 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_830, signal_829, signal_286}), .a ({signal_604, signal_603, signal_173}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789]}), .c ({signal_1088, signal_1087, signal_414}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_400 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_852, signal_851, signal_297}), .a ({signal_656, signal_655, signal_199}), .clk (clk), .r ({Fresh[794], Fresh[793], Fresh[792]}), .c ({signal_1090, signal_1089, signal_415}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_401 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_832, signal_831, signal_287}), .a ({signal_854, signal_853, signal_298}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795]}), .c ({signal_1092, signal_1091, signal_416}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_402 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_846, signal_845, signal_294}), .a ({signal_646, signal_645, signal_194}), .clk (clk), .r ({Fresh[800], Fresh[799], Fresh[798]}), .c ({signal_1094, signal_1093, signal_417}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_403 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_858, signal_857, signal_300}), .a ({signal_856, signal_855, signal_299}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801]}), .c ({signal_1096, signal_1095, signal_418}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_404 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_732, signal_731, signal_237}), .a ({signal_768, signal_767, signal_255}), .clk (clk), .r ({Fresh[806], Fresh[805], Fresh[804]}), .c ({signal_1098, signal_1097, signal_419}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_405 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_650, signal_649, signal_196}), .a ({signal_594, signal_593, signal_168}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807]}), .c ({signal_1100, signal_1099, signal_420}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_406 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_860, signal_859, signal_301}), .a ({signal_780, signal_779, signal_261}), .clk (clk), .r ({Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_1102, signal_1101, signal_421}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_407 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_610, signal_609, signal_176}), .a ({signal_840, signal_839, signal_291}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813]}), .c ({signal_1104, signal_1103, signal_422}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_408 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_812, signal_811, signal_277}), .a ({signal_612, signal_611, signal_177}), .clk (clk), .r ({Fresh[818], Fresh[817], Fresh[816]}), .c ({signal_1106, signal_1105, signal_423}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_409 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_862, signal_861, signal_302}), .a ({signal_812, signal_811, signal_277}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819]}), .c ({signal_1108, signal_1107, signal_424}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_410 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({1'b0, 1'b0, 1'b1}), .a ({signal_702, signal_701, signal_222}), .clk (clk), .r ({Fresh[824], Fresh[823], Fresh[822]}), .c ({signal_1110, signal_1109, signal_425}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_411 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_864, signal_863, signal_303}), .a ({signal_782, signal_781, signal_262}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825]}), .c ({signal_1112, signal_1111, signal_426}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_412 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_866, signal_865, signal_304}), .a ({signal_760, signal_759, signal_251}), .clk (clk), .r ({Fresh[830], Fresh[829], Fresh[828]}), .c ({signal_1114, signal_1113, signal_427}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_413 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_570, signal_569, signal_156}), .a ({signal_818, signal_817, signal_280}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831]}), .c ({signal_1116, signal_1115, signal_428}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_414 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_868, signal_867, signal_305}), .a ({signal_810, signal_809, signal_276}), .clk (clk), .r ({Fresh[836], Fresh[835], Fresh[834]}), .c ({signal_1118, signal_1117, signal_429}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_415 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_854, signal_853, signal_298}), .a ({signal_708, signal_707, signal_225}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837]}), .c ({signal_1120, signal_1119, signal_430}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_416 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_870, signal_869, signal_306}), .a ({signal_584, signal_583, signal_163}), .clk (clk), .r ({Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_1122, signal_1121, signal_431}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_417 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_614, signal_613, signal_178}), .a ({signal_872, signal_871, signal_307}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843]}), .c ({signal_1124, signal_1123, signal_432}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_418 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_874, signal_873, signal_308}), .a ({signal_616, signal_615, signal_179}), .clk (clk), .r ({Fresh[848], Fresh[847], Fresh[846]}), .c ({signal_1126, signal_1125, signal_433}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_419 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_876, signal_875, signal_309}), .a ({signal_866, signal_865, signal_304}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849]}), .c ({signal_1128, signal_1127, signal_434}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_420 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_878, signal_877, signal_310}), .a ({signal_812, signal_811, signal_277}), .clk (clk), .r ({Fresh[854], Fresh[853], Fresh[852]}), .c ({signal_1130, signal_1129, signal_435}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_421 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_690, signal_689, signal_216}), .a ({signal_700, signal_699, signal_221}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855]}), .c ({signal_1132, signal_1131, signal_436}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_422 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_850, signal_849, signal_296}), .a ({signal_600, signal_599, signal_171}), .clk (clk), .r ({Fresh[860], Fresh[859], Fresh[858]}), .c ({signal_1134, signal_1133, signal_437}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_423 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_884, signal_883, signal_312}), .a ({signal_696, signal_695, signal_219}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861]}), .c ({signal_1136, signal_1135, signal_438}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_424 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_680, signal_679, signal_211}), .a ({signal_886, signal_885, signal_313}), .clk (clk), .r ({Fresh[866], Fresh[865], Fresh[864]}), .c ({signal_1138, signal_1137, signal_439}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_425 ( .s ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_784, signal_783, signal_263}), .a ({signal_678, signal_677, signal_210}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867]}), .c ({signal_1140, signal_1139, signal_440}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_426 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_890, signal_889, signal_315}), .a ({signal_888, signal_887, signal_314}), .clk (clk), .r ({Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_1144, signal_1143, signal_441}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_427 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_894, signal_893, signal_317}), .a ({signal_892, signal_891, signal_316}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873]}), .c ({signal_1146, signal_1145, signal_442}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_428 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_898, signal_897, signal_319}), .a ({signal_896, signal_895, signal_318}), .clk (clk), .r ({Fresh[878], Fresh[877], Fresh[876]}), .c ({signal_1148, signal_1147, signal_443}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_429 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_902, signal_901, signal_321}), .a ({signal_900, signal_899, signal_320}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879]}), .c ({signal_1150, signal_1149, signal_444}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_430 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_906, signal_905, signal_323}), .a ({signal_904, signal_903, signal_322}), .clk (clk), .r ({Fresh[884], Fresh[883], Fresh[882]}), .c ({signal_1152, signal_1151, signal_445}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_431 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_910, signal_909, signal_325}), .a ({signal_908, signal_907, signal_324}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885]}), .c ({signal_1154, signal_1153, signal_446}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_432 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_914, signal_913, signal_327}), .a ({signal_912, signal_911, signal_326}), .clk (clk), .r ({Fresh[890], Fresh[889], Fresh[888]}), .c ({signal_1156, signal_1155, signal_447}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_433 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_918, signal_917, signal_329}), .a ({signal_916, signal_915, signal_328}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891]}), .c ({signal_1158, signal_1157, signal_448}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_434 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_922, signal_921, signal_331}), .a ({signal_920, signal_919, signal_330}), .clk (clk), .r ({Fresh[896], Fresh[895], Fresh[894]}), .c ({signal_1160, signal_1159, signal_449}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_435 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_926, signal_925, signal_333}), .a ({signal_924, signal_923, signal_332}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897]}), .c ({signal_1162, signal_1161, signal_450}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_436 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_930, signal_929, signal_335}), .a ({signal_928, signal_927, signal_334}), .clk (clk), .r ({Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_1164, signal_1163, signal_451}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_437 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_934, signal_933, signal_337}), .a ({signal_932, signal_931, signal_336}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903]}), .c ({signal_1166, signal_1165, signal_452}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_438 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_938, signal_937, signal_339}), .a ({signal_936, signal_935, signal_338}), .clk (clk), .r ({Fresh[908], Fresh[907], Fresh[906]}), .c ({signal_1168, signal_1167, signal_453}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_439 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_942, signal_941, signal_341}), .a ({signal_940, signal_939, signal_340}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909]}), .c ({signal_1170, signal_1169, signal_454}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_440 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_946, signal_945, signal_343}), .a ({signal_944, signal_943, signal_342}), .clk (clk), .r ({Fresh[914], Fresh[913], Fresh[912]}), .c ({signal_1172, signal_1171, signal_455}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_441 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_950, signal_949, signal_345}), .a ({signal_948, signal_947, signal_344}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915]}), .c ({signal_1174, signal_1173, signal_456}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_442 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_954, signal_953, signal_347}), .a ({signal_952, signal_951, signal_346}), .clk (clk), .r ({Fresh[920], Fresh[919], Fresh[918]}), .c ({signal_1176, signal_1175, signal_457}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_443 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_958, signal_957, signal_349}), .a ({signal_956, signal_955, signal_348}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921]}), .c ({signal_1178, signal_1177, signal_458}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_444 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_962, signal_961, signal_351}), .a ({signal_960, signal_959, signal_350}), .clk (clk), .r ({Fresh[926], Fresh[925], Fresh[924]}), .c ({signal_1180, signal_1179, signal_459}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_445 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_966, signal_965, signal_353}), .a ({signal_964, signal_963, signal_352}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927]}), .c ({signal_1182, signal_1181, signal_460}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_446 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_970, signal_969, signal_355}), .a ({signal_968, signal_967, signal_354}), .clk (clk), .r ({Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_1184, signal_1183, signal_461}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_447 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_974, signal_973, signal_357}), .a ({signal_972, signal_971, signal_356}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933]}), .c ({signal_1186, signal_1185, signal_462}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_448 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_978, signal_977, signal_359}), .a ({signal_976, signal_975, signal_358}), .clk (clk), .r ({Fresh[938], Fresh[937], Fresh[936]}), .c ({signal_1188, signal_1187, signal_463}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_449 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_982, signal_981, signal_361}), .a ({signal_980, signal_979, signal_360}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939]}), .c ({signal_1190, signal_1189, signal_464}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_450 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_986, signal_985, signal_363}), .a ({signal_984, signal_983, signal_362}), .clk (clk), .r ({Fresh[944], Fresh[943], Fresh[942]}), .c ({signal_1192, signal_1191, signal_465}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_451 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_990, signal_989, signal_365}), .a ({signal_988, signal_987, signal_364}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945]}), .c ({signal_1194, signal_1193, signal_466}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_452 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_994, signal_993, signal_367}), .a ({signal_992, signal_991, signal_366}), .clk (clk), .r ({Fresh[950], Fresh[949], Fresh[948]}), .c ({signal_1196, signal_1195, signal_467}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_453 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_998, signal_997, signal_369}), .a ({signal_996, signal_995, signal_368}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951]}), .c ({signal_1198, signal_1197, signal_468}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_454 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1002, signal_1001, signal_371}), .a ({signal_1000, signal_999, signal_370}), .clk (clk), .r ({Fresh[956], Fresh[955], Fresh[954]}), .c ({signal_1200, signal_1199, signal_469}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_455 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1006, signal_1005, signal_373}), .a ({signal_1004, signal_1003, signal_372}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957]}), .c ({signal_1202, signal_1201, signal_470}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_456 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1010, signal_1009, signal_375}), .a ({signal_1008, signal_1007, signal_374}), .clk (clk), .r ({Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_1204, signal_1203, signal_471}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_457 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1014, signal_1013, signal_377}), .a ({signal_1012, signal_1011, signal_376}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963]}), .c ({signal_1206, signal_1205, signal_472}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_458 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1018, signal_1017, signal_379}), .a ({signal_1016, signal_1015, signal_378}), .clk (clk), .r ({Fresh[968], Fresh[967], Fresh[966]}), .c ({signal_1208, signal_1207, signal_473}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_459 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1022, signal_1021, signal_381}), .a ({signal_1020, signal_1019, signal_380}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969]}), .c ({signal_1210, signal_1209, signal_474}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_460 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1026, signal_1025, signal_383}), .a ({signal_1024, signal_1023, signal_382}), .clk (clk), .r ({Fresh[974], Fresh[973], Fresh[972]}), .c ({signal_1212, signal_1211, signal_475}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_461 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1030, signal_1029, signal_385}), .a ({signal_1028, signal_1027, signal_384}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975]}), .c ({signal_1214, signal_1213, signal_476}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_462 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1034, signal_1033, signal_387}), .a ({signal_1032, signal_1031, signal_386}), .clk (clk), .r ({Fresh[980], Fresh[979], Fresh[978]}), .c ({signal_1216, signal_1215, signal_477}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_463 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1038, signal_1037, signal_389}), .a ({signal_1036, signal_1035, signal_388}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981]}), .c ({signal_1218, signal_1217, signal_478}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_464 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1042, signal_1041, signal_391}), .a ({signal_1040, signal_1039, signal_390}), .clk (clk), .r ({Fresh[986], Fresh[985], Fresh[984]}), .c ({signal_1220, signal_1219, signal_479}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_465 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1046, signal_1045, signal_393}), .a ({signal_1044, signal_1043, signal_392}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987]}), .c ({signal_1222, signal_1221, signal_480}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_466 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1050, signal_1049, signal_395}), .a ({signal_1048, signal_1047, signal_394}), .clk (clk), .r ({Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_1224, signal_1223, signal_481}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_467 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1054, signal_1053, signal_397}), .a ({signal_1052, signal_1051, signal_396}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993]}), .c ({signal_1226, signal_1225, signal_482}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_468 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1058, signal_1057, signal_399}), .a ({signal_1056, signal_1055, signal_398}), .clk (clk), .r ({Fresh[998], Fresh[997], Fresh[996]}), .c ({signal_1228, signal_1227, signal_483}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_469 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1062, signal_1061, signal_401}), .a ({signal_1060, signal_1059, signal_400}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999]}), .c ({signal_1230, signal_1229, signal_484}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_470 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1066, signal_1065, signal_403}), .a ({signal_1064, signal_1063, signal_402}), .clk (clk), .r ({Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({signal_1232, signal_1231, signal_485}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_471 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1070, signal_1069, signal_405}), .a ({signal_1068, signal_1067, signal_404}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005]}), .c ({signal_1234, signal_1233, signal_486}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_472 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1074, signal_1073, signal_407}), .a ({signal_1072, signal_1071, signal_406}), .clk (clk), .r ({Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({signal_1236, signal_1235, signal_487}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_473 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1078, signal_1077, signal_409}), .a ({signal_1076, signal_1075, signal_408}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011]}), .c ({signal_1238, signal_1237, signal_488}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_474 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1082, signal_1081, signal_411}), .a ({signal_1080, signal_1079, signal_410}), .clk (clk), .r ({Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({signal_1240, signal_1239, signal_489}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_475 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1086, signal_1085, signal_413}), .a ({signal_1084, signal_1083, signal_412}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017]}), .c ({signal_1242, signal_1241, signal_490}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_476 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1090, signal_1089, signal_415}), .a ({signal_1088, signal_1087, signal_414}), .clk (clk), .r ({Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_1244, signal_1243, signal_491}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_477 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1094, signal_1093, signal_417}), .a ({signal_1092, signal_1091, signal_416}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023]}), .c ({signal_1246, signal_1245, signal_492}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_478 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1098, signal_1097, signal_419}), .a ({signal_1096, signal_1095, signal_418}), .clk (clk), .r ({Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({signal_1248, signal_1247, signal_493}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_479 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1102, signal_1101, signal_421}), .a ({signal_1100, signal_1099, signal_420}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029]}), .c ({signal_1250, signal_1249, signal_494}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_480 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1106, signal_1105, signal_423}), .a ({signal_1104, signal_1103, signal_422}), .clk (clk), .r ({Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({signal_1252, signal_1251, signal_495}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_481 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1110, signal_1109, signal_425}), .a ({signal_1108, signal_1107, signal_424}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035]}), .c ({signal_1254, signal_1253, signal_496}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_482 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1114, signal_1113, signal_427}), .a ({signal_1112, signal_1111, signal_426}), .clk (clk), .r ({Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({signal_1256, signal_1255, signal_497}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_483 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1118, signal_1117, signal_429}), .a ({signal_1116, signal_1115, signal_428}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041]}), .c ({signal_1258, signal_1257, signal_498}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_484 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1122, signal_1121, signal_431}), .a ({signal_1120, signal_1119, signal_430}), .clk (clk), .r ({Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({signal_1260, signal_1259, signal_499}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_485 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1126, signal_1125, signal_433}), .a ({signal_1124, signal_1123, signal_432}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047]}), .c ({signal_1262, signal_1261, signal_500}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_486 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1130, signal_1129, signal_435}), .a ({signal_1128, signal_1127, signal_434}), .clk (clk), .r ({Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_1264, signal_1263, signal_501}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_487 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1134, signal_1133, signal_437}), .a ({signal_1132, signal_1131, signal_436}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053]}), .c ({signal_1266, signal_1265, signal_502}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_488 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1136, signal_1135, signal_438}), .a ({signal_882, signal_881, signal_311}), .clk (clk), .r ({Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({signal_1268, signal_1267, signal_503}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_489 ( .s ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_1140, signal_1139, signal_440}), .a ({signal_1138, signal_1137, signal_439}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059]}), .c ({signal_1270, signal_1269, signal_504}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_490 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1146, signal_1145, signal_442}), .a ({signal_1144, signal_1143, signal_441}), .clk (clk), .r ({Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({signal_1274, signal_1273, signal_505}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_491 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1150, signal_1149, signal_444}), .a ({signal_1148, signal_1147, signal_443}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065]}), .c ({signal_1276, signal_1275, signal_506}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_492 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1154, signal_1153, signal_446}), .a ({signal_1152, signal_1151, signal_445}), .clk (clk), .r ({Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({signal_1278, signal_1277, signal_507}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_493 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1158, signal_1157, signal_448}), .a ({signal_1156, signal_1155, signal_447}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071]}), .c ({signal_1280, signal_1279, signal_508}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_494 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1162, signal_1161, signal_450}), .a ({signal_1160, signal_1159, signal_449}), .clk (clk), .r ({Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({signal_1282, signal_1281, signal_509}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_495 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1166, signal_1165, signal_452}), .a ({signal_1164, signal_1163, signal_451}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077]}), .c ({signal_1284, signal_1283, signal_510}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_496 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1170, signal_1169, signal_454}), .a ({signal_1168, signal_1167, signal_453}), .clk (clk), .r ({Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_1286, signal_1285, signal_511}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_497 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1174, signal_1173, signal_456}), .a ({signal_1172, signal_1171, signal_455}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083]}), .c ({signal_1288, signal_1287, signal_512}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_498 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1178, signal_1177, signal_458}), .a ({signal_1176, signal_1175, signal_457}), .clk (clk), .r ({Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({signal_1290, signal_1289, signal_513}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_499 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1182, signal_1181, signal_460}), .a ({signal_1180, signal_1179, signal_459}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089]}), .c ({signal_1292, signal_1291, signal_514}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_500 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1186, signal_1185, signal_462}), .a ({signal_1184, signal_1183, signal_461}), .clk (clk), .r ({Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({signal_1294, signal_1293, signal_515}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_501 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1190, signal_1189, signal_464}), .a ({signal_1188, signal_1187, signal_463}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095]}), .c ({signal_1296, signal_1295, signal_516}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_502 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1194, signal_1193, signal_466}), .a ({signal_1192, signal_1191, signal_465}), .clk (clk), .r ({Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({signal_1298, signal_1297, signal_517}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_503 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1198, signal_1197, signal_468}), .a ({signal_1196, signal_1195, signal_467}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101]}), .c ({signal_1300, signal_1299, signal_518}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_504 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1202, signal_1201, signal_470}), .a ({signal_1200, signal_1199, signal_469}), .clk (clk), .r ({Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({signal_1302, signal_1301, signal_519}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_505 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1206, signal_1205, signal_472}), .a ({signal_1204, signal_1203, signal_471}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107]}), .c ({signal_1304, signal_1303, signal_520}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_506 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1210, signal_1209, signal_474}), .a ({signal_1208, signal_1207, signal_473}), .clk (clk), .r ({Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_1306, signal_1305, signal_521}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_507 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1214, signal_1213, signal_476}), .a ({signal_1212, signal_1211, signal_475}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113]}), .c ({signal_1308, signal_1307, signal_522}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_508 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1218, signal_1217, signal_478}), .a ({signal_1216, signal_1215, signal_477}), .clk (clk), .r ({Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({signal_1310, signal_1309, signal_523}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_509 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1222, signal_1221, signal_480}), .a ({signal_1220, signal_1219, signal_479}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119]}), .c ({signal_1312, signal_1311, signal_524}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_510 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1226, signal_1225, signal_482}), .a ({signal_1224, signal_1223, signal_481}), .clk (clk), .r ({Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({signal_1314, signal_1313, signal_525}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_511 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1230, signal_1229, signal_484}), .a ({signal_1228, signal_1227, signal_483}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125]}), .c ({signal_1316, signal_1315, signal_526}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_512 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1234, signal_1233, signal_486}), .a ({signal_1232, signal_1231, signal_485}), .clk (clk), .r ({Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({signal_1318, signal_1317, signal_527}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_513 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1238, signal_1237, signal_488}), .a ({signal_1236, signal_1235, signal_487}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131]}), .c ({signal_1320, signal_1319, signal_528}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_514 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1242, signal_1241, signal_490}), .a ({signal_1240, signal_1239, signal_489}), .clk (clk), .r ({Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({signal_1322, signal_1321, signal_529}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_515 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1246, signal_1245, signal_492}), .a ({signal_1244, signal_1243, signal_491}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137]}), .c ({signal_1324, signal_1323, signal_530}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_516 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1250, signal_1249, signal_494}), .a ({signal_1248, signal_1247, signal_493}), .clk (clk), .r ({Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_1326, signal_1325, signal_531}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_517 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1254, signal_1253, signal_496}), .a ({signal_1252, signal_1251, signal_495}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143]}), .c ({signal_1328, signal_1327, signal_532}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_518 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1258, signal_1257, signal_498}), .a ({signal_1256, signal_1255, signal_497}), .clk (clk), .r ({Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({signal_1330, signal_1329, signal_533}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_519 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1262, signal_1261, signal_500}), .a ({signal_1260, signal_1259, signal_499}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149]}), .c ({signal_1332, signal_1331, signal_534}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_520 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1266, signal_1265, signal_502}), .a ({signal_1264, signal_1263, signal_501}), .clk (clk), .r ({Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({signal_1334, signal_1333, signal_535}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_521 ( .s ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_1270, signal_1269, signal_504}), .a ({signal_1268, signal_1267, signal_503}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155]}), .c ({signal_1336, signal_1335, signal_536}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_522 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1276, signal_1275, signal_506}), .a ({signal_1274, signal_1273, signal_505}), .clk (clk), .r ({Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({signal_1340, signal_1339, signal_537}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_523 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1280, signal_1279, signal_508}), .a ({signal_1278, signal_1277, signal_507}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161]}), .c ({signal_1342, signal_1341, signal_538}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_524 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1284, signal_1283, signal_510}), .a ({signal_1282, signal_1281, signal_509}), .clk (clk), .r ({Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({signal_1344, signal_1343, signal_539}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_525 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1288, signal_1287, signal_512}), .a ({signal_1286, signal_1285, signal_511}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167]}), .c ({signal_1346, signal_1345, signal_540}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_526 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1292, signal_1291, signal_514}), .a ({signal_1290, signal_1289, signal_513}), .clk (clk), .r ({Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_1348, signal_1347, signal_541}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_527 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1296, signal_1295, signal_516}), .a ({signal_1294, signal_1293, signal_515}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173]}), .c ({signal_1350, signal_1349, signal_542}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_528 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1300, signal_1299, signal_518}), .a ({signal_1298, signal_1297, signal_517}), .clk (clk), .r ({Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({signal_1352, signal_1351, signal_543}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_529 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1304, signal_1303, signal_520}), .a ({signal_1302, signal_1301, signal_519}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179]}), .c ({signal_1354, signal_1353, signal_544}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_530 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1308, signal_1307, signal_522}), .a ({signal_1306, signal_1305, signal_521}), .clk (clk), .r ({Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({signal_1356, signal_1355, signal_545}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_531 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1312, signal_1311, signal_524}), .a ({signal_1310, signal_1309, signal_523}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185]}), .c ({signal_1358, signal_1357, signal_546}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_532 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1316, signal_1315, signal_526}), .a ({signal_1314, signal_1313, signal_525}), .clk (clk), .r ({Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({signal_1360, signal_1359, signal_547}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_533 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1320, signal_1319, signal_528}), .a ({signal_1318, signal_1317, signal_527}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191]}), .c ({signal_1362, signal_1361, signal_548}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_534 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1324, signal_1323, signal_530}), .a ({signal_1322, signal_1321, signal_529}), .clk (clk), .r ({Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({signal_1364, signal_1363, signal_549}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_535 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1328, signal_1327, signal_532}), .a ({signal_1326, signal_1325, signal_531}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197]}), .c ({signal_1366, signal_1365, signal_550}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_536 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1332, signal_1331, signal_534}), .a ({signal_1330, signal_1329, signal_533}), .clk (clk), .r ({Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_1368, signal_1367, signal_551}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_537 ( .s ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_1336, signal_1335, signal_536}), .a ({signal_1334, signal_1333, signal_535}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203]}), .c ({signal_1370, signal_1369, signal_552}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_538 ( .s ({X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_1342, signal_1341, signal_538}), .a ({signal_1340, signal_1339, signal_537}), .clk (clk), .r ({Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({signal_1374, signal_1373, signal_150}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_539 ( .s ({X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_1346, signal_1345, signal_540}), .a ({signal_1344, signal_1343, signal_539}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209]}), .c ({signal_1376, signal_1375, signal_149}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_540 ( .s ({X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_1350, signal_1349, signal_542}), .a ({signal_1348, signal_1347, signal_541}), .clk (clk), .r ({Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({signal_1378, signal_1377, signal_148}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_541 ( .s ({X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_1354, signal_1353, signal_544}), .a ({signal_1352, signal_1351, signal_543}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215]}), .c ({signal_1380, signal_1379, signal_147}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_542 ( .s ({X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_1358, signal_1357, signal_546}), .a ({signal_1356, signal_1355, signal_545}), .clk (clk), .r ({Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({signal_1382, signal_1381, signal_146}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_543 ( .s ({X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_1362, signal_1361, signal_548}), .a ({signal_1360, signal_1359, signal_547}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221]}), .c ({signal_1384, signal_1383, signal_145}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_544 ( .s ({X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_1366, signal_1365, signal_550}), .a ({signal_1364, signal_1363, signal_549}), .clk (clk), .r ({Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({signal_1386, signal_1385, signal_144}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(0)) cell_545 ( .s ({X_s2[7], X_s1[7], X_s0[7]}), .b ({signal_1370, signal_1369, signal_552}), .a ({signal_1368, signal_1367, signal_551}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227]}), .c ({signal_1388, signal_1387, signal_143}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(0)) cell_0 ( .clk (signal_2636), .D ({signal_1388, signal_1387, signal_143}), .Q ({Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_1 ( .clk (signal_2636), .D ({signal_1386, signal_1385, signal_144}), .Q ({Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_2 ( .clk (signal_2636), .D ({signal_1384, signal_1383, signal_145}), .Q ({Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_3 ( .clk (signal_2636), .D ({signal_1382, signal_1381, signal_146}), .Q ({Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_4 ( .clk (signal_2636), .D ({signal_1380, signal_1379, signal_147}), .Q ({Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_5 ( .clk (signal_2636), .D ({signal_1378, signal_1377, signal_148}), .Q ({Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_6 ( .clk (signal_2636), .D ({signal_1376, signal_1375, signal_149}), .Q ({Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_7 ( .clk (signal_2636), .D ({signal_1374, signal_1373, signal_150}), .Q ({Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
