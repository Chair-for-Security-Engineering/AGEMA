/* modified netlist. Source: module sbox in file ../sbox_lookup/sbox.v */
/* 10 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 11 register stage(s) in total */

module sbox_HPC1_Pipeline_d3 (SI_s0, clk, SI_s1, SI_s2, SI_s3, Fresh, SO_s0, SO_s1, SO_s2, SO_s3);
    input [3:0] SI_s0 ;
    input clk ;
    input [3:0] SI_s1 ;
    input [3:0] SI_s2 ;
    input [3:0] SI_s3 ;
    input [129:0] Fresh ;
    output [3:0] SO_s0 ;
    output [3:0] SO_s1 ;
    output [3:0] SO_s2 ;
    output [3:0] SO_s3 ;
    wire N9 ;
    wire N12 ;
    wire N19 ;
    wire N27 ;
    wire n40 ;
    wire n41 ;
    wire n42 ;
    wire n43 ;
    wire n44 ;
    wire n45 ;
    wire n46 ;
    wire n47 ;
    wire n48 ;
    wire n49 ;
    wire n50 ;
    wire n51 ;
    wire n52 ;
    wire n53 ;
    wire n54 ;
    wire new_AGEMA_signal_37 ;
    wire new_AGEMA_signal_38 ;
    wire new_AGEMA_signal_39 ;
    wire new_AGEMA_signal_46 ;
    wire new_AGEMA_signal_47 ;
    wire new_AGEMA_signal_48 ;
    wire new_AGEMA_signal_52 ;
    wire new_AGEMA_signal_53 ;
    wire new_AGEMA_signal_54 ;
    wire new_AGEMA_signal_55 ;
    wire new_AGEMA_signal_56 ;
    wire new_AGEMA_signal_57 ;
    wire new_AGEMA_signal_58 ;
    wire new_AGEMA_signal_59 ;
    wire new_AGEMA_signal_60 ;
    wire new_AGEMA_signal_61 ;
    wire new_AGEMA_signal_62 ;
    wire new_AGEMA_signal_63 ;
    wire new_AGEMA_signal_64 ;
    wire new_AGEMA_signal_65 ;
    wire new_AGEMA_signal_66 ;
    wire new_AGEMA_signal_67 ;
    wire new_AGEMA_signal_68 ;
    wire new_AGEMA_signal_69 ;
    wire new_AGEMA_signal_70 ;
    wire new_AGEMA_signal_71 ;
    wire new_AGEMA_signal_72 ;
    wire new_AGEMA_signal_73 ;
    wire new_AGEMA_signal_74 ;
    wire new_AGEMA_signal_75 ;
    wire new_AGEMA_signal_76 ;
    wire new_AGEMA_signal_77 ;
    wire new_AGEMA_signal_78 ;
    wire new_AGEMA_signal_79 ;
    wire new_AGEMA_signal_80 ;
    wire new_AGEMA_signal_81 ;
    wire new_AGEMA_signal_82 ;
    wire new_AGEMA_signal_83 ;
    wire new_AGEMA_signal_84 ;
    wire new_AGEMA_signal_85 ;
    wire new_AGEMA_signal_86 ;
    wire new_AGEMA_signal_87 ;
    wire new_AGEMA_signal_88 ;
    wire new_AGEMA_signal_89 ;
    wire new_AGEMA_signal_90 ;
    wire new_AGEMA_signal_91 ;
    wire new_AGEMA_signal_92 ;
    wire new_AGEMA_signal_93 ;
    wire new_AGEMA_signal_94 ;
    wire new_AGEMA_signal_95 ;
    wire new_AGEMA_signal_96 ;
    wire new_AGEMA_signal_97 ;
    wire new_AGEMA_signal_98 ;
    wire new_AGEMA_signal_99 ;
    wire new_AGEMA_signal_100 ;
    wire new_AGEMA_signal_101 ;
    wire new_AGEMA_signal_102 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(1)) U50 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_39, new_AGEMA_signal_38, new_AGEMA_signal_37, n53}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U53 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_54, new_AGEMA_signal_53, new_AGEMA_signal_52, n52}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U59 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, n51}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_23 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( new_AGEMA_signal_245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_25 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( new_AGEMA_signal_247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_27 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( new_AGEMA_signal_249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_29 ( .C ( clk ), .D ( SI_s3[3] ), .Q ( new_AGEMA_signal_251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_31 ( .C ( clk ), .D ( n53 ), .Q ( new_AGEMA_signal_253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_33 ( .C ( clk ), .D ( new_AGEMA_signal_37 ), .Q ( new_AGEMA_signal_255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_35 ( .C ( clk ), .D ( new_AGEMA_signal_38 ), .Q ( new_AGEMA_signal_257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_37 ( .C ( clk ), .D ( new_AGEMA_signal_39 ), .Q ( new_AGEMA_signal_259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_39 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( new_AGEMA_signal_261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_41 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( new_AGEMA_signal_263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_43 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( new_AGEMA_signal_265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_45 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( new_AGEMA_signal_267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_47 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( new_AGEMA_signal_269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_49 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( new_AGEMA_signal_271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_51 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( new_AGEMA_signal_273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_53 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( new_AGEMA_signal_275 ) ) ;

    /* cells in depth 2 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U51 ( .ina ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .inb ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .outt ({new_AGEMA_signal_48, new_AGEMA_signal_47, new_AGEMA_signal_46, n40}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) U52 ( .a ({new_AGEMA_signal_48, new_AGEMA_signal_47, new_AGEMA_signal_46, n40}), .b ({new_AGEMA_signal_252, new_AGEMA_signal_250, new_AGEMA_signal_248, new_AGEMA_signal_246}), .c ({new_AGEMA_signal_66, new_AGEMA_signal_65, new_AGEMA_signal_64, N12}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U54 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_54, new_AGEMA_signal_53, new_AGEMA_signal_52, n52}), .clk ( clk ), .rnd ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .outt ({new_AGEMA_signal_69, new_AGEMA_signal_68, new_AGEMA_signal_67, n41}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(1)) U55 ( .a ({new_AGEMA_signal_260, new_AGEMA_signal_258, new_AGEMA_signal_256, new_AGEMA_signal_254}), .b ({new_AGEMA_signal_69, new_AGEMA_signal_68, new_AGEMA_signal_67, n41}), .c ({new_AGEMA_signal_87, new_AGEMA_signal_86, new_AGEMA_signal_85, n42}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U57 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .outt ({new_AGEMA_signal_57, new_AGEMA_signal_56, new_AGEMA_signal_55, n43}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U60 ( .ina ({new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, n51}), .inb ({new_AGEMA_signal_39, new_AGEMA_signal_38, new_AGEMA_signal_37, n53}), .clk ( clk ), .rnd ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .outt ({new_AGEMA_signal_75, new_AGEMA_signal_74, new_AGEMA_signal_73, n45}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U61 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .outt ({new_AGEMA_signal_63, new_AGEMA_signal_62, new_AGEMA_signal_61, n48}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U67 ( .ina ({new_AGEMA_signal_54, new_AGEMA_signal_53, new_AGEMA_signal_52, n52}), .inb ({new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, n51}), .clk ( clk ), .rnd ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .outt ({new_AGEMA_signal_84, new_AGEMA_signal_83, new_AGEMA_signal_82, n54}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) U68 ( .a ({new_AGEMA_signal_84, new_AGEMA_signal_83, new_AGEMA_signal_82, n54}), .b ({new_AGEMA_signal_260, new_AGEMA_signal_258, new_AGEMA_signal_256, new_AGEMA_signal_254}), .c ({new_AGEMA_signal_93, new_AGEMA_signal_92, new_AGEMA_signal_91, N9}) ) ;
    buf_clk new_AGEMA_reg_buffer_24 ( .C ( clk ), .D ( new_AGEMA_signal_245 ), .Q ( new_AGEMA_signal_246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_26 ( .C ( clk ), .D ( new_AGEMA_signal_247 ), .Q ( new_AGEMA_signal_248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_28 ( .C ( clk ), .D ( new_AGEMA_signal_249 ), .Q ( new_AGEMA_signal_250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_30 ( .C ( clk ), .D ( new_AGEMA_signal_251 ), .Q ( new_AGEMA_signal_252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_32 ( .C ( clk ), .D ( new_AGEMA_signal_253 ), .Q ( new_AGEMA_signal_254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_34 ( .C ( clk ), .D ( new_AGEMA_signal_255 ), .Q ( new_AGEMA_signal_256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_36 ( .C ( clk ), .D ( new_AGEMA_signal_257 ), .Q ( new_AGEMA_signal_258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_38 ( .C ( clk ), .D ( new_AGEMA_signal_259 ), .Q ( new_AGEMA_signal_260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_40 ( .C ( clk ), .D ( new_AGEMA_signal_261 ), .Q ( new_AGEMA_signal_262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_42 ( .C ( clk ), .D ( new_AGEMA_signal_263 ), .Q ( new_AGEMA_signal_264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_44 ( .C ( clk ), .D ( new_AGEMA_signal_265 ), .Q ( new_AGEMA_signal_266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_46 ( .C ( clk ), .D ( new_AGEMA_signal_267 ), .Q ( new_AGEMA_signal_268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_48 ( .C ( clk ), .D ( new_AGEMA_signal_269 ), .Q ( new_AGEMA_signal_270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_50 ( .C ( clk ), .D ( new_AGEMA_signal_271 ), .Q ( new_AGEMA_signal_272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_52 ( .C ( clk ), .D ( new_AGEMA_signal_273 ), .Q ( new_AGEMA_signal_274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_54 ( .C ( clk ), .D ( new_AGEMA_signal_275 ), .Q ( new_AGEMA_signal_276 ) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_55 ( .C ( clk ), .D ( n45 ), .Q ( new_AGEMA_signal_277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_57 ( .C ( clk ), .D ( new_AGEMA_signal_73 ), .Q ( new_AGEMA_signal_279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_59 ( .C ( clk ), .D ( new_AGEMA_signal_74 ), .Q ( new_AGEMA_signal_281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_61 ( .C ( clk ), .D ( new_AGEMA_signal_75 ), .Q ( new_AGEMA_signal_283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_63 ( .C ( clk ), .D ( new_AGEMA_signal_262 ), .Q ( new_AGEMA_signal_285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_67 ( .C ( clk ), .D ( new_AGEMA_signal_264 ), .Q ( new_AGEMA_signal_289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_71 ( .C ( clk ), .D ( new_AGEMA_signal_266 ), .Q ( new_AGEMA_signal_293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_75 ( .C ( clk ), .D ( new_AGEMA_signal_268 ), .Q ( new_AGEMA_signal_297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_103 ( .C ( clk ), .D ( N9 ), .Q ( new_AGEMA_signal_325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_111 ( .C ( clk ), .D ( new_AGEMA_signal_91 ), .Q ( new_AGEMA_signal_333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_119 ( .C ( clk ), .D ( new_AGEMA_signal_92 ), .Q ( new_AGEMA_signal_341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_127 ( .C ( clk ), .D ( new_AGEMA_signal_93 ), .Q ( new_AGEMA_signal_349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_135 ( .C ( clk ), .D ( N12 ), .Q ( new_AGEMA_signal_357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_143 ( .C ( clk ), .D ( new_AGEMA_signal_64 ), .Q ( new_AGEMA_signal_365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_151 ( .C ( clk ), .D ( new_AGEMA_signal_65 ), .Q ( new_AGEMA_signal_373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_159 ( .C ( clk ), .D ( new_AGEMA_signal_66 ), .Q ( new_AGEMA_signal_381 ) ) ;

    /* cells in depth 4 */
    mux2_HPC1 #(.security_order(3), .pipeline(1)) U56 ( .ins ({new_AGEMA_signal_268, new_AGEMA_signal_266, new_AGEMA_signal_264, new_AGEMA_signal_262}), .inb ({new_AGEMA_signal_87, new_AGEMA_signal_86, new_AGEMA_signal_85, n42}), .ina ({new_AGEMA_signal_276, new_AGEMA_signal_274, new_AGEMA_signal_272, new_AGEMA_signal_270}), .clk ( clk ), .rnd ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .outt ({new_AGEMA_signal_96, new_AGEMA_signal_95, new_AGEMA_signal_94, N19}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U58 ( .ina ({new_AGEMA_signal_57, new_AGEMA_signal_56, new_AGEMA_signal_55, n43}), .inb ({new_AGEMA_signal_276, new_AGEMA_signal_274, new_AGEMA_signal_272, new_AGEMA_signal_270}), .clk ( clk ), .rnd ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .outt ({new_AGEMA_signal_72, new_AGEMA_signal_71, new_AGEMA_signal_70, n47}) ) ;
    or_HPC1 #(.security_order(3), .pipeline(1)) U62 ( .ina ({new_AGEMA_signal_252, new_AGEMA_signal_250, new_AGEMA_signal_248, new_AGEMA_signal_246}), .inb ({new_AGEMA_signal_63, new_AGEMA_signal_62, new_AGEMA_signal_61, n48}), .clk ( clk ), .rnd ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .outt ({new_AGEMA_signal_78, new_AGEMA_signal_77, new_AGEMA_signal_76, n44}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U65 ( .ina ({new_AGEMA_signal_252, new_AGEMA_signal_250, new_AGEMA_signal_248, new_AGEMA_signal_246}), .inb ({new_AGEMA_signal_63, new_AGEMA_signal_62, new_AGEMA_signal_61, n48}), .clk ( clk ), .rnd ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .outt ({new_AGEMA_signal_81, new_AGEMA_signal_80, new_AGEMA_signal_79, n49}) ) ;
    buf_clk new_AGEMA_reg_buffer_56 ( .C ( clk ), .D ( new_AGEMA_signal_277 ), .Q ( new_AGEMA_signal_278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_58 ( .C ( clk ), .D ( new_AGEMA_signal_279 ), .Q ( new_AGEMA_signal_280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_60 ( .C ( clk ), .D ( new_AGEMA_signal_281 ), .Q ( new_AGEMA_signal_282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_62 ( .C ( clk ), .D ( new_AGEMA_signal_283 ), .Q ( new_AGEMA_signal_284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_64 ( .C ( clk ), .D ( new_AGEMA_signal_285 ), .Q ( new_AGEMA_signal_286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_68 ( .C ( clk ), .D ( new_AGEMA_signal_289 ), .Q ( new_AGEMA_signal_290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_72 ( .C ( clk ), .D ( new_AGEMA_signal_293 ), .Q ( new_AGEMA_signal_294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_76 ( .C ( clk ), .D ( new_AGEMA_signal_297 ), .Q ( new_AGEMA_signal_298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_104 ( .C ( clk ), .D ( new_AGEMA_signal_325 ), .Q ( new_AGEMA_signal_326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_112 ( .C ( clk ), .D ( new_AGEMA_signal_333 ), .Q ( new_AGEMA_signal_334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_120 ( .C ( clk ), .D ( new_AGEMA_signal_341 ), .Q ( new_AGEMA_signal_342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_128 ( .C ( clk ), .D ( new_AGEMA_signal_349 ), .Q ( new_AGEMA_signal_350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_136 ( .C ( clk ), .D ( new_AGEMA_signal_357 ), .Q ( new_AGEMA_signal_358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_144 ( .C ( clk ), .D ( new_AGEMA_signal_365 ), .Q ( new_AGEMA_signal_366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_152 ( .C ( clk ), .D ( new_AGEMA_signal_373 ), .Q ( new_AGEMA_signal_374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_160 ( .C ( clk ), .D ( new_AGEMA_signal_381 ), .Q ( new_AGEMA_signal_382 ) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_65 ( .C ( clk ), .D ( new_AGEMA_signal_286 ), .Q ( new_AGEMA_signal_287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_69 ( .C ( clk ), .D ( new_AGEMA_signal_290 ), .Q ( new_AGEMA_signal_291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_73 ( .C ( clk ), .D ( new_AGEMA_signal_294 ), .Q ( new_AGEMA_signal_295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_77 ( .C ( clk ), .D ( new_AGEMA_signal_298 ), .Q ( new_AGEMA_signal_299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_79 ( .C ( clk ), .D ( n47 ), .Q ( new_AGEMA_signal_301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_81 ( .C ( clk ), .D ( new_AGEMA_signal_70 ), .Q ( new_AGEMA_signal_303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_83 ( .C ( clk ), .D ( new_AGEMA_signal_71 ), .Q ( new_AGEMA_signal_305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_85 ( .C ( clk ), .D ( new_AGEMA_signal_72 ), .Q ( new_AGEMA_signal_307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_87 ( .C ( clk ), .D ( n49 ), .Q ( new_AGEMA_signal_309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_91 ( .C ( clk ), .D ( new_AGEMA_signal_79 ), .Q ( new_AGEMA_signal_313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_95 ( .C ( clk ), .D ( new_AGEMA_signal_80 ), .Q ( new_AGEMA_signal_317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_99 ( .C ( clk ), .D ( new_AGEMA_signal_81 ), .Q ( new_AGEMA_signal_321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_105 ( .C ( clk ), .D ( new_AGEMA_signal_326 ), .Q ( new_AGEMA_signal_327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_113 ( .C ( clk ), .D ( new_AGEMA_signal_334 ), .Q ( new_AGEMA_signal_335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_121 ( .C ( clk ), .D ( new_AGEMA_signal_342 ), .Q ( new_AGEMA_signal_343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_129 ( .C ( clk ), .D ( new_AGEMA_signal_350 ), .Q ( new_AGEMA_signal_351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_137 ( .C ( clk ), .D ( new_AGEMA_signal_358 ), .Q ( new_AGEMA_signal_359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_145 ( .C ( clk ), .D ( new_AGEMA_signal_366 ), .Q ( new_AGEMA_signal_367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_153 ( .C ( clk ), .D ( new_AGEMA_signal_374 ), .Q ( new_AGEMA_signal_375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_161 ( .C ( clk ), .D ( new_AGEMA_signal_382 ), .Q ( new_AGEMA_signal_383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_167 ( .C ( clk ), .D ( N19 ), .Q ( new_AGEMA_signal_389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_173 ( .C ( clk ), .D ( new_AGEMA_signal_94 ), .Q ( new_AGEMA_signal_395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_179 ( .C ( clk ), .D ( new_AGEMA_signal_95 ), .Q ( new_AGEMA_signal_401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_185 ( .C ( clk ), .D ( new_AGEMA_signal_96 ), .Q ( new_AGEMA_signal_407 ) ) ;

    /* cells in depth 6 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U63 ( .ina ({new_AGEMA_signal_284, new_AGEMA_signal_282, new_AGEMA_signal_280, new_AGEMA_signal_278}), .inb ({new_AGEMA_signal_78, new_AGEMA_signal_77, new_AGEMA_signal_76, n44}), .clk ( clk ), .rnd ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .outt ({new_AGEMA_signal_90, new_AGEMA_signal_89, new_AGEMA_signal_88, n46}) ) ;
    buf_clk new_AGEMA_reg_buffer_66 ( .C ( clk ), .D ( new_AGEMA_signal_287 ), .Q ( new_AGEMA_signal_288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_70 ( .C ( clk ), .D ( new_AGEMA_signal_291 ), .Q ( new_AGEMA_signal_292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_74 ( .C ( clk ), .D ( new_AGEMA_signal_295 ), .Q ( new_AGEMA_signal_296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_78 ( .C ( clk ), .D ( new_AGEMA_signal_299 ), .Q ( new_AGEMA_signal_300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_80 ( .C ( clk ), .D ( new_AGEMA_signal_301 ), .Q ( new_AGEMA_signal_302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_82 ( .C ( clk ), .D ( new_AGEMA_signal_303 ), .Q ( new_AGEMA_signal_304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_84 ( .C ( clk ), .D ( new_AGEMA_signal_305 ), .Q ( new_AGEMA_signal_306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_86 ( .C ( clk ), .D ( new_AGEMA_signal_307 ), .Q ( new_AGEMA_signal_308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_88 ( .C ( clk ), .D ( new_AGEMA_signal_309 ), .Q ( new_AGEMA_signal_310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_92 ( .C ( clk ), .D ( new_AGEMA_signal_313 ), .Q ( new_AGEMA_signal_314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_96 ( .C ( clk ), .D ( new_AGEMA_signal_317 ), .Q ( new_AGEMA_signal_318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_100 ( .C ( clk ), .D ( new_AGEMA_signal_321 ), .Q ( new_AGEMA_signal_322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_106 ( .C ( clk ), .D ( new_AGEMA_signal_327 ), .Q ( new_AGEMA_signal_328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_114 ( .C ( clk ), .D ( new_AGEMA_signal_335 ), .Q ( new_AGEMA_signal_336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_122 ( .C ( clk ), .D ( new_AGEMA_signal_343 ), .Q ( new_AGEMA_signal_344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_130 ( .C ( clk ), .D ( new_AGEMA_signal_351 ), .Q ( new_AGEMA_signal_352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_138 ( .C ( clk ), .D ( new_AGEMA_signal_359 ), .Q ( new_AGEMA_signal_360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_146 ( .C ( clk ), .D ( new_AGEMA_signal_367 ), .Q ( new_AGEMA_signal_368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_154 ( .C ( clk ), .D ( new_AGEMA_signal_375 ), .Q ( new_AGEMA_signal_376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_162 ( .C ( clk ), .D ( new_AGEMA_signal_383 ), .Q ( new_AGEMA_signal_384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_168 ( .C ( clk ), .D ( new_AGEMA_signal_389 ), .Q ( new_AGEMA_signal_390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_174 ( .C ( clk ), .D ( new_AGEMA_signal_395 ), .Q ( new_AGEMA_signal_396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_180 ( .C ( clk ), .D ( new_AGEMA_signal_401 ), .Q ( new_AGEMA_signal_402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_186 ( .C ( clk ), .D ( new_AGEMA_signal_407 ), .Q ( new_AGEMA_signal_408 ) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_89 ( .C ( clk ), .D ( new_AGEMA_signal_310 ), .Q ( new_AGEMA_signal_311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_93 ( .C ( clk ), .D ( new_AGEMA_signal_314 ), .Q ( new_AGEMA_signal_315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_97 ( .C ( clk ), .D ( new_AGEMA_signal_318 ), .Q ( new_AGEMA_signal_319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_101 ( .C ( clk ), .D ( new_AGEMA_signal_322 ), .Q ( new_AGEMA_signal_323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_107 ( .C ( clk ), .D ( new_AGEMA_signal_328 ), .Q ( new_AGEMA_signal_329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_115 ( .C ( clk ), .D ( new_AGEMA_signal_336 ), .Q ( new_AGEMA_signal_337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_123 ( .C ( clk ), .D ( new_AGEMA_signal_344 ), .Q ( new_AGEMA_signal_345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_131 ( .C ( clk ), .D ( new_AGEMA_signal_352 ), .Q ( new_AGEMA_signal_353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_139 ( .C ( clk ), .D ( new_AGEMA_signal_360 ), .Q ( new_AGEMA_signal_361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_147 ( .C ( clk ), .D ( new_AGEMA_signal_368 ), .Q ( new_AGEMA_signal_369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_155 ( .C ( clk ), .D ( new_AGEMA_signal_376 ), .Q ( new_AGEMA_signal_377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_163 ( .C ( clk ), .D ( new_AGEMA_signal_384 ), .Q ( new_AGEMA_signal_385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_169 ( .C ( clk ), .D ( new_AGEMA_signal_390 ), .Q ( new_AGEMA_signal_391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_175 ( .C ( clk ), .D ( new_AGEMA_signal_396 ), .Q ( new_AGEMA_signal_397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_181 ( .C ( clk ), .D ( new_AGEMA_signal_402 ), .Q ( new_AGEMA_signal_403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_187 ( .C ( clk ), .D ( new_AGEMA_signal_408 ), .Q ( new_AGEMA_signal_409 ) ) ;

    /* cells in depth 8 */
    mux2_HPC1 #(.security_order(3), .pipeline(1)) U64 ( .ins ({new_AGEMA_signal_300, new_AGEMA_signal_296, new_AGEMA_signal_292, new_AGEMA_signal_288}), .inb ({new_AGEMA_signal_308, new_AGEMA_signal_306, new_AGEMA_signal_304, new_AGEMA_signal_302}), .ina ({new_AGEMA_signal_90, new_AGEMA_signal_89, new_AGEMA_signal_88, n46}), .clk ( clk ), .rnd ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .outt ({new_AGEMA_signal_99, new_AGEMA_signal_98, new_AGEMA_signal_97, n50}) ) ;
    buf_clk new_AGEMA_reg_buffer_90 ( .C ( clk ), .D ( new_AGEMA_signal_311 ), .Q ( new_AGEMA_signal_312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_94 ( .C ( clk ), .D ( new_AGEMA_signal_315 ), .Q ( new_AGEMA_signal_316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_98 ( .C ( clk ), .D ( new_AGEMA_signal_319 ), .Q ( new_AGEMA_signal_320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_102 ( .C ( clk ), .D ( new_AGEMA_signal_323 ), .Q ( new_AGEMA_signal_324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_108 ( .C ( clk ), .D ( new_AGEMA_signal_329 ), .Q ( new_AGEMA_signal_330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_116 ( .C ( clk ), .D ( new_AGEMA_signal_337 ), .Q ( new_AGEMA_signal_338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_124 ( .C ( clk ), .D ( new_AGEMA_signal_345 ), .Q ( new_AGEMA_signal_346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_132 ( .C ( clk ), .D ( new_AGEMA_signal_353 ), .Q ( new_AGEMA_signal_354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_140 ( .C ( clk ), .D ( new_AGEMA_signal_361 ), .Q ( new_AGEMA_signal_362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_148 ( .C ( clk ), .D ( new_AGEMA_signal_369 ), .Q ( new_AGEMA_signal_370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_156 ( .C ( clk ), .D ( new_AGEMA_signal_377 ), .Q ( new_AGEMA_signal_378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_164 ( .C ( clk ), .D ( new_AGEMA_signal_385 ), .Q ( new_AGEMA_signal_386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_170 ( .C ( clk ), .D ( new_AGEMA_signal_391 ), .Q ( new_AGEMA_signal_392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_176 ( .C ( clk ), .D ( new_AGEMA_signal_397 ), .Q ( new_AGEMA_signal_398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_182 ( .C ( clk ), .D ( new_AGEMA_signal_403 ), .Q ( new_AGEMA_signal_404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_188 ( .C ( clk ), .D ( new_AGEMA_signal_409 ), .Q ( new_AGEMA_signal_410 ) ) ;

    /* cells in depth 9 */
    buf_clk new_AGEMA_reg_buffer_109 ( .C ( clk ), .D ( new_AGEMA_signal_330 ), .Q ( new_AGEMA_signal_331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_117 ( .C ( clk ), .D ( new_AGEMA_signal_338 ), .Q ( new_AGEMA_signal_339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_125 ( .C ( clk ), .D ( new_AGEMA_signal_346 ), .Q ( new_AGEMA_signal_347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_133 ( .C ( clk ), .D ( new_AGEMA_signal_354 ), .Q ( new_AGEMA_signal_355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_141 ( .C ( clk ), .D ( new_AGEMA_signal_362 ), .Q ( new_AGEMA_signal_363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_149 ( .C ( clk ), .D ( new_AGEMA_signal_370 ), .Q ( new_AGEMA_signal_371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_157 ( .C ( clk ), .D ( new_AGEMA_signal_378 ), .Q ( new_AGEMA_signal_379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_165 ( .C ( clk ), .D ( new_AGEMA_signal_386 ), .Q ( new_AGEMA_signal_387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_171 ( .C ( clk ), .D ( new_AGEMA_signal_392 ), .Q ( new_AGEMA_signal_393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_177 ( .C ( clk ), .D ( new_AGEMA_signal_398 ), .Q ( new_AGEMA_signal_399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_183 ( .C ( clk ), .D ( new_AGEMA_signal_404 ), .Q ( new_AGEMA_signal_405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_189 ( .C ( clk ), .D ( new_AGEMA_signal_410 ), .Q ( new_AGEMA_signal_411 ) ) ;

    /* cells in depth 10 */
    nand_HPC1 #(.security_order(3), .pipeline(1)) U66 ( .ina ({new_AGEMA_signal_99, new_AGEMA_signal_98, new_AGEMA_signal_97, n50}), .inb ({new_AGEMA_signal_324, new_AGEMA_signal_320, new_AGEMA_signal_316, new_AGEMA_signal_312}), .clk ( clk ), .rnd ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .outt ({new_AGEMA_signal_102, new_AGEMA_signal_101, new_AGEMA_signal_100, N27}) ) ;
    buf_clk new_AGEMA_reg_buffer_110 ( .C ( clk ), .D ( new_AGEMA_signal_331 ), .Q ( new_AGEMA_signal_332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_118 ( .C ( clk ), .D ( new_AGEMA_signal_339 ), .Q ( new_AGEMA_signal_340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_126 ( .C ( clk ), .D ( new_AGEMA_signal_347 ), .Q ( new_AGEMA_signal_348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_134 ( .C ( clk ), .D ( new_AGEMA_signal_355 ), .Q ( new_AGEMA_signal_356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_142 ( .C ( clk ), .D ( new_AGEMA_signal_363 ), .Q ( new_AGEMA_signal_364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_150 ( .C ( clk ), .D ( new_AGEMA_signal_371 ), .Q ( new_AGEMA_signal_372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_158 ( .C ( clk ), .D ( new_AGEMA_signal_379 ), .Q ( new_AGEMA_signal_380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_166 ( .C ( clk ), .D ( new_AGEMA_signal_387 ), .Q ( new_AGEMA_signal_388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_172 ( .C ( clk ), .D ( new_AGEMA_signal_393 ), .Q ( new_AGEMA_signal_394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_178 ( .C ( clk ), .D ( new_AGEMA_signal_399 ), .Q ( new_AGEMA_signal_400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_184 ( .C ( clk ), .D ( new_AGEMA_signal_405 ), .Q ( new_AGEMA_signal_406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_190 ( .C ( clk ), .D ( new_AGEMA_signal_411 ), .Q ( new_AGEMA_signal_412 ) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_356, new_AGEMA_signal_348, new_AGEMA_signal_340, new_AGEMA_signal_332}), .Q ({SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_388, new_AGEMA_signal_380, new_AGEMA_signal_372, new_AGEMA_signal_364}), .Q ({SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_412, new_AGEMA_signal_406, new_AGEMA_signal_400, new_AGEMA_signal_394}), .Q ({SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_102, new_AGEMA_signal_101, new_AGEMA_signal_100, N27}), .Q ({SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
