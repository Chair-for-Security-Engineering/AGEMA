/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module sbox_HPC2_AIG_ClockGating_d4 (X_s0, clk, X_s1, X_s2, X_s3, X_s4, Fresh, rst, Y_s0, Y_s1, Y_s2, Y_s3, Y_s4, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [7:0] X_s4 ;
    input rst ;
    input [339:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    output [7:0] Y_s4 ;
    output Synch ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_1208 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_136 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_286, signal_285, signal_284, signal_283, signal_151}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_137 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_294, signal_293, signal_292, signal_291, signal_152}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_138 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_302, signal_301, signal_300, signal_299, signal_153}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_139 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_306, signal_305, signal_304, signal_303, signal_154}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_140 ( .a ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_314, signal_313, signal_312, signal_311, signal_155}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_141 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .c ({signal_326, signal_325, signal_324, signal_323, signal_156}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_142 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_330, signal_329, signal_328, signal_327, signal_157}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_143 ( .a ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_334, signal_333, signal_332, signal_331, signal_158}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_144 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_342, signal_341, signal_340, signal_339, signal_159}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_145 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_346, signal_345, signal_344, signal_343, signal_160}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_146 ( .a ({signal_286, signal_285, signal_284, signal_283, signal_151}), .b ({signal_314, signal_313, signal_312, signal_311, signal_155}), .c ({signal_350, signal_349, signal_348, signal_347, signal_161}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_147 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_326, signal_325, signal_324, signal_323, signal_156}), .c ({signal_354, signal_353, signal_352, signal_351, signal_162}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_148 ( .a ({signal_302, signal_301, signal_300, signal_299, signal_153}), .b ({signal_306, signal_305, signal_304, signal_303, signal_154}), .c ({signal_358, signal_357, signal_356, signal_355, signal_163}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_149 ( .a ({signal_314, signal_313, signal_312, signal_311, signal_155}), .b ({signal_330, signal_329, signal_328, signal_327, signal_157}), .c ({signal_362, signal_361, signal_360, signal_359, signal_164}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_150 ( .a ({signal_314, signal_313, signal_312, signal_311, signal_155}), .b ({signal_334, signal_333, signal_332, signal_331, signal_158}), .c ({signal_366, signal_365, signal_364, signal_363, signal_165}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_151 ( .a ({signal_326, signal_325, signal_324, signal_323, signal_156}), .b ({signal_342, signal_341, signal_340, signal_339, signal_159}), .c ({signal_370, signal_369, signal_368, signal_367, signal_166}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_152 ( .a ({signal_326, signal_325, signal_324, signal_323, signal_156}), .b ({signal_346, signal_345, signal_344, signal_343, signal_160}), .c ({signal_374, signal_373, signal_372, signal_371, signal_167}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_153 ( .a ({signal_286, signal_285, signal_284, signal_283, signal_151}), .b ({signal_334, signal_333, signal_332, signal_331, signal_158}), .c ({signal_378, signal_377, signal_376, signal_375, signal_168}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_160 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_350, signal_349, signal_348, signal_347, signal_161}), .c ({signal_406, signal_405, signal_404, signal_403, signal_175}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_161 ( .a ({signal_326, signal_325, signal_324, signal_323, signal_156}), .b ({signal_350, signal_349, signal_348, signal_347, signal_161}), .c ({signal_410, signal_409, signal_408, signal_407, signal_176}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_162 ( .a ({signal_330, signal_329, signal_328, signal_327, signal_157}), .b ({signal_350, signal_349, signal_348, signal_347, signal_161}), .c ({signal_414, signal_413, signal_412, signal_411, signal_177}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_163 ( .a ({signal_354, signal_353, signal_352, signal_351, signal_162}), .b ({signal_366, signal_365, signal_364, signal_363, signal_165}), .c ({signal_418, signal_417, signal_416, signal_415, signal_178}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_164 ( .a ({signal_286, signal_285, signal_284, signal_283, signal_151}), .b ({signal_370, signal_369, signal_368, signal_367, signal_166}), .c ({signal_422, signal_421, signal_420, signal_419, signal_179}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_165 ( .a ({signal_294, signal_293, signal_292, signal_291, signal_152}), .b ({signal_374, signal_373, signal_372, signal_371, signal_167}), .c ({signal_426, signal_425, signal_424, signal_423, signal_180}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_166 ( .a ({signal_302, signal_301, signal_300, signal_299, signal_153}), .b ({signal_366, signal_365, signal_364, signal_363, signal_165}), .c ({signal_430, signal_429, signal_428, signal_427, signal_181}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_170 ( .a ({signal_294, signal_293, signal_292, signal_291, signal_152}), .b ({signal_410, signal_409, signal_408, signal_407, signal_176}), .c ({signal_446, signal_445, signal_444, signal_443, signal_185}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_171 ( .a ({signal_418, signal_417, signal_416, signal_415, signal_178}), .b ({signal_422, signal_421, signal_420, signal_419, signal_179}), .c ({signal_450, signal_449, signal_448, signal_447, signal_186}) ) ;
    ClockGatingController #(9) cell_268 ( .clk (clk), .rst (rst), .GatedClk (signal_1208), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_154 ( .a ({signal_350, signal_349, signal_348, signal_347, signal_161}), .b ({signal_358, signal_357, signal_356, signal_355, signal_163}), .clk (clk), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_382, signal_381, signal_380, signal_379, signal_169}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_155 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_370, signal_369, signal_368, signal_367, signal_166}), .clk (clk), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({signal_386, signal_385, signal_384, signal_383, signal_170}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_156 ( .a ({signal_302, signal_301, signal_300, signal_299, signal_153}), .b ({signal_366, signal_365, signal_364, signal_363, signal_165}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({signal_390, signal_389, signal_388, signal_387, signal_171}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_157 ( .a ({signal_354, signal_353, signal_352, signal_351, signal_162}), .b ({signal_374, signal_373, signal_372, signal_371, signal_167}), .clk (clk), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_394, signal_393, signal_392, signal_391, signal_172}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_158 ( .a ({signal_286, signal_285, signal_284, signal_283, signal_151}), .b ({signal_362, signal_361, signal_360, signal_359, signal_164}), .clk (clk), .r ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({signal_398, signal_397, signal_396, signal_395, signal_173}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_159 ( .a ({signal_306, signal_305, signal_304, signal_303, signal_154}), .b ({signal_378, signal_377, signal_376, signal_375, signal_168}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .c ({signal_402, signal_401, signal_400, signal_399, signal_174}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_167 ( .a ({signal_406, signal_405, signal_404, signal_403, signal_175}), .b ({signal_426, signal_425, signal_424, signal_423, signal_180}), .clk (clk), .r ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_434, signal_433, signal_432, signal_431, signal_182}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_168 ( .a ({signal_418, signal_417, signal_416, signal_415, signal_178}), .b ({signal_422, signal_421, signal_420, signal_419, signal_179}), .clk (clk), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .c ({signal_438, signal_437, signal_436, signal_435, signal_183}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_169 ( .a ({signal_294, signal_293, signal_292, signal_291, signal_152}), .b ({signal_410, signal_409, signal_408, signal_407, signal_176}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({signal_442, signal_441, signal_440, signal_439, signal_184}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_172 ( .a ({signal_414, signal_413, signal_412, signal_411, signal_177}), .b ({signal_382, signal_381, signal_380, signal_379, signal_169}), .c ({signal_454, signal_453, signal_452, signal_451, signal_187}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_173 ( .a ({signal_382, signal_381, signal_380, signal_379, signal_169}), .b ({signal_386, signal_385, signal_384, signal_383, signal_170}), .c ({signal_458, signal_457, signal_456, signal_455, signal_188}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_174 ( .a ({signal_430, signal_429, signal_428, signal_427, signal_181}), .b ({signal_390, signal_389, signal_388, signal_387, signal_171}), .c ({signal_462, signal_461, signal_460, signal_459, signal_189}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_175 ( .a ({signal_398, signal_397, signal_396, signal_395, signal_173}), .b ({signal_402, signal_401, signal_400, signal_399, signal_174}), .c ({signal_466, signal_465, signal_464, signal_463, signal_190}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_176 ( .a ({signal_390, signal_389, signal_388, signal_387, signal_171}), .b ({signal_438, signal_437, signal_436, signal_435, signal_183}), .c ({signal_470, signal_469, signal_468, signal_467, signal_191}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_177 ( .a ({signal_398, signal_397, signal_396, signal_395, signal_173}), .b ({signal_442, signal_441, signal_440, signal_439, signal_184}), .c ({signal_474, signal_473, signal_472, signal_471, signal_192}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_178 ( .a ({signal_434, signal_433, signal_432, signal_431, signal_182}), .b ({signal_454, signal_453, signal_452, signal_451, signal_187}), .c ({signal_478, signal_477, signal_476, signal_475, signal_193}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_179 ( .a ({signal_446, signal_445, signal_444, signal_443, signal_185}), .b ({signal_458, signal_457, signal_456, signal_455, signal_188}), .c ({signal_482, signal_481, signal_480, signal_479, signal_194}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_180 ( .a ({signal_394, signal_393, signal_392, signal_391, signal_172}), .b ({signal_462, signal_461, signal_460, signal_459, signal_189}), .c ({signal_486, signal_485, signal_484, signal_483, signal_195}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_181 ( .a ({signal_470, signal_469, signal_468, signal_467, signal_191}), .b ({signal_474, signal_473, signal_472, signal_471, signal_192}), .c ({signal_490, signal_489, signal_488, signal_487, signal_196}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_182 ( .a ({signal_466, signal_465, signal_464, signal_463, signal_190}), .b ({signal_478, signal_477, signal_476, signal_475, signal_193}), .c ({signal_494, signal_493, signal_492, signal_491, signal_197}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_183 ( .a ({signal_474, signal_473, signal_472, signal_471, signal_192}), .b ({signal_482, signal_481, signal_480, signal_479, signal_194}), .c ({signal_498, signal_497, signal_496, signal_495, signal_198}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_184 ( .a ({signal_466, signal_465, signal_464, signal_463, signal_190}), .b ({signal_486, signal_485, signal_484, signal_483, signal_195}), .c ({signal_502, signal_501, signal_500, signal_499, signal_199}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_187 ( .a ({signal_450, signal_449, signal_448, signal_447, signal_186}), .b ({signal_490, signal_489, signal_488, signal_487, signal_196}), .c ({signal_514, signal_513, signal_512, signal_511, signal_202}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_188 ( .a ({signal_494, signal_493, signal_492, signal_491, signal_197}), .b ({signal_498, signal_497, signal_496, signal_495, signal_198}), .c ({signal_518, signal_517, signal_516, signal_515, signal_203}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_190 ( .a ({signal_502, signal_501, signal_500, signal_499, signal_199}), .b ({signal_514, signal_513, signal_512, signal_511, signal_202}), .c ({signal_526, signal_525, signal_524, signal_523, signal_205}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_185 ( .a ({signal_494, signal_493, signal_492, signal_491, signal_197}), .b ({signal_502, signal_501, signal_500, signal_499, signal_199}), .clk (clk), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_506, signal_505, signal_504, signal_503, signal_200}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_186 ( .a ({signal_498, signal_497, signal_496, signal_495, signal_198}), .b ({signal_502, signal_501, signal_500, signal_499, signal_199}), .clk (clk), .r ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({signal_510, signal_509, signal_508, signal_507, signal_201}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_189 ( .a ({signal_494, signal_493, signal_492, signal_491, signal_197}), .b ({signal_514, signal_513, signal_512, signal_511, signal_202}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .c ({signal_522, signal_521, signal_520, signal_519, signal_204}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_191 ( .a ({signal_498, signal_497, signal_496, signal_495, signal_198}), .b ({signal_506, signal_505, signal_504, signal_503, signal_200}), .c ({signal_530, signal_529, signal_528, signal_527, signal_206}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_192 ( .a ({signal_514, signal_513, signal_512, signal_511, signal_202}), .b ({signal_506, signal_505, signal_504, signal_503, signal_200}), .c ({signal_534, signal_533, signal_532, signal_531, signal_207}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_193 ( .a ({signal_506, signal_505, signal_504, signal_503, signal_200}), .b ({signal_518, signal_517, signal_516, signal_515, signal_203}), .c ({signal_538, signal_537, signal_536, signal_535, signal_208}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_198 ( .a ({signal_506, signal_505, signal_504, signal_503, signal_200}), .b ({signal_526, signal_525, signal_524, signal_523, signal_205}), .c ({signal_558, signal_557, signal_556, signal_555, signal_213}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_194 ( .a ({signal_518, signal_517, signal_516, signal_515, signal_203}), .b ({signal_534, signal_533, signal_532, signal_531, signal_207}), .clk (clk), .r ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_542, signal_541, signal_540, signal_539, signal_209}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_195 ( .a ({signal_526, signal_525, signal_524, signal_523, signal_205}), .b ({signal_530, signal_529, signal_528, signal_527, signal_206}), .clk (clk), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .c ({signal_546, signal_545, signal_544, signal_543, signal_210}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_196 ( .a ({signal_518, signal_517, signal_516, signal_515, signal_203}), .b ({signal_522, signal_521, signal_520, signal_519, signal_204}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({signal_550, signal_549, signal_548, signal_547, signal_211}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_197 ( .a ({signal_510, signal_509, signal_508, signal_507, signal_201}), .b ({signal_526, signal_525, signal_524, signal_523, signal_205}), .clk (clk), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_554, signal_553, signal_552, signal_551, signal_212}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_199 ( .a ({signal_498, signal_497, signal_496, signal_495, signal_198}), .b ({signal_542, signal_541, signal_540, signal_539, signal_209}), .c ({signal_562, signal_561, signal_560, signal_559, signal_214}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_200 ( .a ({signal_538, signal_537, signal_536, signal_535, signal_208}), .b ({signal_550, signal_549, signal_548, signal_547, signal_211}), .c ({signal_566, signal_565, signal_564, signal_563, signal_215}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_201 ( .a ({signal_514, signal_513, signal_512, signal_511, signal_202}), .b ({signal_546, signal_545, signal_544, signal_543, signal_210}), .c ({signal_570, signal_569, signal_568, signal_567, signal_216}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_202 ( .a ({signal_554, signal_553, signal_552, signal_551, signal_212}), .b ({signal_558, signal_557, signal_556, signal_555, signal_213}), .c ({signal_574, signal_573, signal_572, signal_571, signal_217}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_211 ( .a ({signal_566, signal_565, signal_564, signal_563, signal_215}), .b ({signal_574, signal_573, signal_572, signal_571, signal_217}), .c ({signal_610, signal_609, signal_608, signal_607, signal_226}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_212 ( .a ({signal_562, signal_561, signal_560, signal_559, signal_214}), .b ({signal_570, signal_569, signal_568, signal_567, signal_216}), .c ({signal_614, signal_613, signal_612, signal_611, signal_227}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_213 ( .a ({signal_562, signal_561, signal_560, signal_559, signal_214}), .b ({signal_566, signal_565, signal_564, signal_563, signal_215}), .c ({signal_618, signal_617, signal_616, signal_615, signal_228}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_214 ( .a ({signal_570, signal_569, signal_568, signal_567, signal_216}), .b ({signal_574, signal_573, signal_572, signal_571, signal_217}), .c ({signal_622, signal_621, signal_620, signal_619, signal_229}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_223 ( .a ({signal_610, signal_609, signal_608, signal_607, signal_226}), .b ({signal_614, signal_613, signal_612, signal_611, signal_227}), .c ({signal_658, signal_657, signal_656, signal_655, signal_238}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_203 ( .a ({signal_406, signal_405, signal_404, signal_403, signal_175}), .b ({signal_574, signal_573, signal_572, signal_571, signal_217}), .clk (clk), .r ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .c ({signal_578, signal_577, signal_576, signal_575, signal_218}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_204 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_570, signal_569, signal_568, signal_567, signal_216}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .c ({signal_582, signal_581, signal_580, signal_579, signal_219}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_205 ( .a ({signal_354, signal_353, signal_352, signal_351, signal_162}), .b ({signal_566, signal_565, signal_564, signal_563, signal_215}), .clk (clk), .r ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_586, signal_585, signal_584, signal_583, signal_220}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_206 ( .a ({signal_418, signal_417, signal_416, signal_415, signal_178}), .b ({signal_562, signal_561, signal_560, signal_559, signal_214}), .clk (clk), .r ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .c ({signal_590, signal_589, signal_588, signal_587, signal_221}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_207 ( .a ({signal_426, signal_425, signal_424, signal_423, signal_180}), .b ({signal_574, signal_573, signal_572, signal_571, signal_217}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .c ({signal_594, signal_593, signal_592, signal_591, signal_222}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_208 ( .a ({signal_370, signal_369, signal_368, signal_367, signal_166}), .b ({signal_570, signal_569, signal_568, signal_567, signal_216}), .clk (clk), .r ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_598, signal_597, signal_596, signal_595, signal_223}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_209 ( .a ({signal_374, signal_373, signal_372, signal_371, signal_167}), .b ({signal_566, signal_565, signal_564, signal_563, signal_215}), .clk (clk), .r ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .c ({signal_602, signal_601, signal_600, signal_599, signal_224}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_210 ( .a ({signal_422, signal_421, signal_420, signal_419, signal_179}), .b ({signal_562, signal_561, signal_560, signal_559, signal_214}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .c ({signal_606, signal_605, signal_604, signal_603, signal_225}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_215 ( .a ({signal_350, signal_349, signal_348, signal_347, signal_161}), .b ({signal_622, signal_621, signal_620, signal_619, signal_229}), .clk (clk), .r ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_626, signal_625, signal_624, signal_623, signal_230}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_216 ( .a ({signal_366, signal_365, signal_364, signal_363, signal_165}), .b ({signal_618, signal_617, signal_616, signal_615, signal_228}), .clk (clk), .r ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .c ({signal_630, signal_629, signal_628, signal_627, signal_231}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_217 ( .a ({signal_362, signal_361, signal_360, signal_359, signal_164}), .b ({signal_614, signal_613, signal_612, signal_611, signal_227}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .c ({signal_634, signal_633, signal_632, signal_631, signal_232}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_218 ( .a ({signal_410, signal_409, signal_408, signal_407, signal_176}), .b ({signal_610, signal_609, signal_608, signal_607, signal_226}), .clk (clk), .r ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_638, signal_637, signal_636, signal_635, signal_233}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_219 ( .a ({signal_358, signal_357, signal_356, signal_355, signal_163}), .b ({signal_622, signal_621, signal_620, signal_619, signal_229}), .clk (clk), .r ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .c ({signal_642, signal_641, signal_640, signal_639, signal_234}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_220 ( .a ({signal_302, signal_301, signal_300, signal_299, signal_153}), .b ({signal_618, signal_617, signal_616, signal_615, signal_228}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .c ({signal_646, signal_645, signal_644, signal_643, signal_235}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_221 ( .a ({signal_286, signal_285, signal_284, signal_283, signal_151}), .b ({signal_614, signal_613, signal_612, signal_611, signal_227}), .clk (clk), .r ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_650, signal_649, signal_648, signal_647, signal_236}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_222 ( .a ({signal_294, signal_293, signal_292, signal_291, signal_152}), .b ({signal_610, signal_609, signal_608, signal_607, signal_226}), .clk (clk), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .c ({signal_654, signal_653, signal_652, signal_651, signal_237}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_224 ( .a ({signal_586, signal_585, signal_584, signal_583, signal_220}), .b ({signal_594, signal_593, signal_592, signal_591, signal_222}), .c ({signal_662, signal_661, signal_660, signal_659, signal_239}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_225 ( .a ({signal_590, signal_589, signal_588, signal_587, signal_221}), .b ({signal_602, signal_601, signal_600, signal_599, signal_224}), .c ({signal_666, signal_665, signal_664, signal_663, signal_240}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_226 ( .a ({signal_582, signal_581, signal_580, signal_579, signal_219}), .b ({signal_590, signal_589, signal_588, signal_587, signal_221}), .c ({signal_670, signal_669, signal_668, signal_667, signal_241}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_227 ( .a ({signal_378, signal_377, signal_376, signal_375, signal_168}), .b ({signal_658, signal_657, signal_656, signal_655, signal_238}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .c ({signal_674, signal_673, signal_672, signal_671, signal_242}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_228 ( .a ({signal_306, signal_305, signal_304, signal_303, signal_154}), .b ({signal_658, signal_657, signal_656, signal_655, signal_238}), .clk (clk), .r ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_678, signal_677, signal_676, signal_675, signal_243}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_229 ( .a ({signal_582, signal_581, signal_580, signal_579, signal_219}), .b ({signal_626, signal_625, signal_624, signal_623, signal_230}), .c ({signal_682, signal_681, signal_680, signal_679, signal_244}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_230 ( .a ({signal_578, signal_577, signal_576, signal_575, signal_218}), .b ({signal_642, signal_641, signal_640, signal_639, signal_234}), .c ({signal_686, signal_685, signal_684, signal_683, signal_245}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_231 ( .a ({signal_638, signal_637, signal_636, signal_635, signal_233}), .b ({signal_646, signal_645, signal_644, signal_643, signal_235}), .c ({signal_690, signal_689, signal_688, signal_687, signal_246}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_232 ( .a ({signal_630, signal_629, signal_628, signal_627, signal_231}), .b ({signal_650, signal_649, signal_648, signal_647, signal_236}), .c ({signal_694, signal_693, signal_692, signal_691, signal_247}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_233 ( .a ({signal_634, signal_633, signal_632, signal_631, signal_232}), .b ({signal_650, signal_649, signal_648, signal_647, signal_236}), .c ({signal_698, signal_697, signal_696, signal_695, signal_248}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_234 ( .a ({signal_642, signal_641, signal_640, signal_639, signal_234}), .b ({signal_662, signal_661, signal_660, signal_659, signal_239}), .c ({signal_702, signal_701, signal_700, signal_699, signal_249}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_235 ( .a ({signal_598, signal_597, signal_596, signal_595, signal_223}), .b ({signal_662, signal_661, signal_660, signal_659, signal_239}), .c ({signal_706, signal_705, signal_704, signal_703, signal_250}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_236 ( .a ({signal_646, signal_645, signal_644, signal_643, signal_235}), .b ({signal_666, signal_665, signal_664, signal_663, signal_240}), .c ({signal_710, signal_709, signal_708, signal_707, signal_251}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_237 ( .a ({signal_650, signal_649, signal_648, signal_647, signal_236}), .b ({signal_678, signal_677, signal_676, signal_675, signal_243}), .c ({signal_714, signal_713, signal_712, signal_711, signal_252}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_238 ( .a ({signal_678, signal_677, signal_676, signal_675, signal_243}), .b ({signal_694, signal_693, signal_692, signal_691, signal_247}), .c ({signal_718, signal_717, signal_716, signal_715, signal_253}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_239 ( .a ({signal_626, signal_625, signal_624, signal_623, signal_230}), .b ({signal_686, signal_685, signal_684, signal_683, signal_245}), .c ({signal_722, signal_721, signal_720, signal_719, signal_254}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_240 ( .a ({signal_634, signal_633, signal_632, signal_631, signal_232}), .b ({signal_674, signal_673, signal_672, signal_671, signal_242}), .c ({signal_726, signal_725, signal_724, signal_723, signal_255}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_241 ( .a ({signal_674, signal_673, signal_672, signal_671, signal_242}), .b ({signal_690, signal_689, signal_688, signal_687, signal_246}), .c ({signal_730, signal_729, signal_728, signal_727, signal_256}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_242 ( .a ({signal_606, signal_605, signal_604, signal_603, signal_225}), .b ({signal_682, signal_681, signal_680, signal_679, signal_244}), .c ({signal_734, signal_733, signal_732, signal_731, signal_257}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_243 ( .a ({signal_654, signal_653, signal_652, signal_651, signal_237}), .b ({signal_690, signal_689, signal_688, signal_687, signal_246}), .c ({signal_738, signal_737, signal_736, signal_735, signal_258}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_244 ( .a ({signal_670, signal_669, signal_668, signal_667, signal_241}), .b ({signal_686, signal_685, signal_684, signal_683, signal_245}), .c ({signal_742, signal_741, signal_740, signal_739, signal_259}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_245 ( .a ({signal_682, signal_681, signal_680, signal_679, signal_244}), .b ({signal_710, signal_709, signal_708, signal_707, signal_251}), .c ({signal_746, signal_745, signal_744, signal_743, signal_260}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_246 ( .a ({signal_586, signal_585, signal_584, signal_583, signal_220}), .b ({signal_714, signal_713, signal_712, signal_711, signal_252}), .c ({signal_750, signal_749, signal_748, signal_747, signal_261}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_247 ( .a ({signal_594, signal_593, signal_592, signal_591, signal_222}), .b ({signal_714, signal_713, signal_712, signal_711, signal_252}), .c ({signal_754, signal_753, signal_752, signal_751, signal_262}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_248 ( .a ({signal_662, signal_661, signal_660, signal_659, signal_239}), .b ({signal_714, signal_713, signal_712, signal_711, signal_252}), .c ({signal_758, signal_757, signal_756, signal_755, signal_263}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_249 ( .a ({signal_662, signal_661, signal_660, signal_659, signal_239}), .b ({signal_722, signal_721, signal_720, signal_719, signal_254}), .c ({signal_762, signal_761, signal_760, signal_759, signal_264}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_250 ( .a ({signal_702, signal_701, signal_700, signal_699, signal_249}), .b ({signal_726, signal_725, signal_724, signal_723, signal_255}), .c ({signal_766, signal_765, signal_764, signal_763, signal_265}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_251 ( .a ({signal_718, signal_717, signal_716, signal_715, signal_253}), .b ({signal_730, signal_729, signal_728, signal_727, signal_256}), .c ({signal_770, signal_769, signal_768, signal_767, signal_266}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_252 ( .a ({signal_722, signal_721, signal_720, signal_719, signal_254}), .b ({signal_726, signal_725, signal_724, signal_723, signal_255}), .c ({signal_774, signal_773, signal_772, signal_771, signal_267}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_253 ( .a ({signal_666, signal_665, signal_664, signal_663, signal_240}), .b ({signal_730, signal_729, signal_728, signal_727, signal_256}), .c ({signal_778, signal_777, signal_776, signal_775, signal_268}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_254 ( .a ({signal_698, signal_697, signal_696, signal_695, signal_248}), .b ({signal_734, signal_733, signal_732, signal_731, signal_257}), .c ({signal_782, signal_781, signal_780, signal_779, signal_269}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_255 ( .a ({signal_706, signal_705, signal_704, signal_703, signal_250}), .b ({signal_734, signal_733, signal_732, signal_731, signal_257}), .c ({signal_786, signal_785, signal_784, signal_783, signal_270}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_256 ( .a ({signal_718, signal_717, signal_716, signal_715, signal_253}), .b ({signal_746, signal_745, signal_744, signal_743, signal_260}), .c ({signal_790, signal_789, signal_788, signal_787, signal_271}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_257 ( .a ({signal_790, signal_789, signal_788, signal_787, signal_271}), .b ({signal_794, signal_793, signal_792, signal_791, signal_150}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_258 ( .a ({signal_718, signal_717, signal_716, signal_715, signal_253}), .b ({signal_766, signal_765, signal_764, signal_763, signal_265}), .c ({signal_798, signal_797, signal_796, signal_795, signal_143}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_259 ( .a ({signal_754, signal_753, signal_752, signal_751, signal_262}), .b ({signal_774, signal_773, signal_772, signal_771, signal_267}), .c ({signal_802, signal_801, signal_800, signal_799, signal_272}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_260 ( .a ({signal_738, signal_737, signal_736, signal_735, signal_258}), .b ({signal_782, signal_781, signal_780, signal_779, signal_269}), .c ({signal_806, signal_805, signal_804, signal_803, signal_273}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_261 ( .a ({signal_718, signal_717, signal_716, signal_715, signal_253}), .b ({signal_762, signal_761, signal_760, signal_759, signal_264}), .c ({signal_810, signal_809, signal_808, signal_807, signal_146}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_262 ( .a ({signal_742, signal_741, signal_740, signal_739, signal_259}), .b ({signal_758, signal_757, signal_756, signal_755, signal_263}), .c ({signal_814, signal_813, signal_812, signal_811, signal_147}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_263 ( .a ({signal_770, signal_769, signal_768, signal_767, signal_266}), .b ({signal_786, signal_785, signal_784, signal_783, signal_270}), .c ({signal_818, signal_817, signal_816, signal_815, signal_148}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_264 ( .a ({signal_750, signal_749, signal_748, signal_747, signal_261}), .b ({signal_778, signal_777, signal_776, signal_775, signal_268}), .c ({signal_822, signal_821, signal_820, signal_819, signal_274}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_265 ( .a ({signal_802, signal_801, signal_800, signal_799, signal_272}), .b ({signal_826, signal_825, signal_824, signal_823, signal_144}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_266 ( .a ({signal_806, signal_805, signal_804, signal_803, signal_273}), .b ({signal_830, signal_829, signal_828, signal_827, signal_145}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_267 ( .a ({signal_822, signal_821, signal_820, signal_819, signal_274}), .b ({signal_834, signal_833, signal_832, signal_831, signal_149}) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(0)) cell_0 ( .clk (signal_1208), .D ({signal_798, signal_797, signal_796, signal_795, signal_143}), .Q ({Y_s4[7], Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_1 ( .clk (signal_1208), .D ({signal_826, signal_825, signal_824, signal_823, signal_144}), .Q ({Y_s4[6], Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_2 ( .clk (signal_1208), .D ({signal_830, signal_829, signal_828, signal_827, signal_145}), .Q ({Y_s4[5], Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_3 ( .clk (signal_1208), .D ({signal_810, signal_809, signal_808, signal_807, signal_146}), .Q ({Y_s4[4], Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_4 ( .clk (signal_1208), .D ({signal_814, signal_813, signal_812, signal_811, signal_147}), .Q ({Y_s4[3], Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_5 ( .clk (signal_1208), .D ({signal_818, signal_817, signal_816, signal_815, signal_148}), .Q ({Y_s4[2], Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_6 ( .clk (signal_1208), .D ({signal_834, signal_833, signal_832, signal_831, signal_149}), .Q ({Y_s4[1], Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_7 ( .clk (signal_1208), .D ({signal_794, signal_793, signal_792, signal_791, signal_150}), .Q ({Y_s4[0], Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
