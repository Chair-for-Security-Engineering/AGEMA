/* modified netlist. Source: module sbox in file Designs/AESSbox//Canright/AGEMA/sbox.v */
/* 16 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 17 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d3 (X_s0, clk, X_s1, X_s2, X_s3, Fresh, Y_s0, Y_s1, Y_s2, Y_s3);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [527:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(1)) cell_176 ( .a ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_442, signal_441, signal_440, signal_192}) ) ;
    INV_X1 cell_177 ( .A ( 1'b1 ), .ZN ( signal_193 ) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_178 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_451, signal_450, signal_449, signal_194}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_179 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .c ({signal_460, signal_459, signal_458, signal_195}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_180 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_463, signal_462, signal_461, signal_196}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_181 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_466, signal_465, signal_464, signal_197}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_182 ( .a ({X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_472, signal_471, signal_470, signal_198}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_183 ( .a ({signal_463, signal_462, signal_461, signal_196}), .b ({signal_475, signal_474, signal_473, signal_199}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_186 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_463, signal_462, signal_461, signal_196}), .c ({signal_484, signal_483, signal_482, signal_202}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_187 ( .a ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_460, signal_459, signal_458, signal_195}), .c ({signal_490, signal_489, signal_488, signal_203}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_188 ( .a ({signal_460, signal_459, signal_458, signal_195}), .b ({signal_466, signal_465, signal_464, signal_197}), .c ({signal_493, signal_492, signal_491, signal_204}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_189 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_466, signal_465, signal_464, signal_197}), .c ({signal_499, signal_498, signal_497, signal_205}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_190 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_472, signal_471, signal_470, signal_198}), .c ({signal_502, signal_501, signal_500, signal_206}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_191 ( .a ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_466, signal_465, signal_464, signal_197}), .c ({signal_505, signal_504, signal_503, signal_207}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_192 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_472, signal_471, signal_470, signal_198}), .c ({signal_508, signal_507, signal_506, signal_208}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_193 ( .a ({signal_493, signal_492, signal_491, signal_204}), .b ({signal_511, signal_510, signal_509, signal_209}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_194 ( .a ({signal_505, signal_504, signal_503, signal_207}), .b ({signal_514, signal_513, signal_512, signal_210}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_201 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_505, signal_504, signal_503, signal_207}), .c ({signal_535, signal_534, signal_533, signal_217}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_202 ( .a ({signal_490, signal_489, signal_488, signal_203}), .b ({signal_499, signal_498, signal_497, signal_205}), .c ({signal_538, signal_537, signal_536, signal_218}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_203 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_499, signal_498, signal_497, signal_205}), .c ({signal_541, signal_540, signal_539, signal_219}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_204 ( .a ({X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_499, signal_498, signal_497, signal_205}), .c ({signal_544, signal_543, signal_542, signal_220}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_205 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_505, signal_504, signal_503, signal_207}), .c ({signal_547, signal_546, signal_545, signal_221}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_206 ( .a ({signal_463, signal_462, signal_461, signal_196}), .b ({signal_508, signal_507, signal_506, signal_208}), .c ({signal_550, signal_549, signal_548, signal_222}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_208 ( .a ({signal_535, signal_534, signal_533, signal_217}), .b ({signal_556, signal_555, signal_554, signal_224}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_209 ( .a ({signal_538, signal_537, signal_536, signal_218}), .b ({signal_559, signal_558, signal_557, signal_225}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_210 ( .a ({signal_547, signal_546, signal_545, signal_221}), .b ({signal_562, signal_561, signal_560, signal_226}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_211 ( .a ({signal_550, signal_549, signal_548, signal_222}), .b ({signal_565, signal_564, signal_563, signal_227}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_219 ( .a ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_544, signal_543, signal_542, signal_220}), .c ({signal_589, signal_588, signal_587, signal_235}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_220 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_547, signal_546, signal_545, signal_221}), .c ({signal_592, signal_591, signal_590, signal_236}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_222 ( .a ({signal_589, signal_588, signal_587, signal_235}), .b ({signal_598, signal_597, signal_596, signal_238}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_223 ( .a ({signal_592, signal_591, signal_590, signal_236}), .b ({signal_601, signal_600, signal_599, signal_239}) ) ;

    /* cells in depth 1 */
    buf_clk cell_909 ( .C ( clk ), .D ( signal_193 ), .Q ( signal_2249 ) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_184 ( .a ({signal_442, signal_441, signal_440, signal_192}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_478, signal_477, signal_476, signal_200}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_185 ( .a ({1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_451, signal_450, signal_449, signal_194}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_481, signal_480, signal_479, signal_201}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_195 ( .a ({signal_478, signal_477, signal_476, signal_200}), .b ({signal_517, signal_516, signal_515, signal_211}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_196 ( .a ({signal_481, signal_480, signal_479, signal_201}), .b ({signal_520, signal_519, signal_518, signal_212}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_197 ( .a ({1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_490, signal_489, signal_488, signal_203}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_523, signal_522, signal_521, signal_213}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_198 ( .a ({1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_502, signal_501, signal_500, signal_206}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_526, signal_525, signal_524, signal_214}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_199 ( .a ({1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_475, signal_474, signal_473, signal_199}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_529, signal_528, signal_527, signal_215}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_200 ( .a ({1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_484, signal_483, signal_482, signal_202}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_532, signal_531, signal_530, signal_216}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_207 ( .a ({signal_523, signal_522, signal_521, signal_213}), .b ({signal_553, signal_552, signal_551, signal_223}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_212 ( .a ({signal_526, signal_525, signal_524, signal_214}), .b ({signal_568, signal_567, signal_566, signal_228}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_213 ( .a ({signal_529, signal_528, signal_527, signal_215}), .b ({signal_571, signal_570, signal_569, signal_229}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_214 ( .a ({signal_532, signal_531, signal_530, signal_216}), .b ({signal_574, signal_573, signal_572, signal_230}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_215 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_514, signal_513, signal_512, signal_210}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_577, signal_576, signal_575, signal_231}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_216 ( .a ({1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_541, signal_540, signal_539, signal_219}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_580, signal_579, signal_578, signal_232}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_217 ( .a ({1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_544, signal_543, signal_542, signal_220}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_583, signal_582, signal_581, signal_233}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_218 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_511, signal_510, signal_509, signal_209}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_586, signal_585, signal_584, signal_234}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_221 ( .a ({signal_577, signal_576, signal_575, signal_231}), .b ({signal_595, signal_594, signal_593, signal_237}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_224 ( .a ({signal_580, signal_579, signal_578, signal_232}), .b ({signal_604, signal_603, signal_602, signal_240}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_225 ( .a ({signal_583, signal_582, signal_581, signal_233}), .b ({signal_607, signal_606, signal_605, signal_241}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_226 ( .a ({signal_586, signal_585, signal_584, signal_234}), .b ({signal_610, signal_609, signal_608, signal_242}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_228 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_559, signal_558, signal_557, signal_225}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_616, signal_615, signal_614, signal_244}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_229 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_562, signal_561, signal_560, signal_226}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_619, signal_618, signal_617, signal_245}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_230 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_556, signal_555, signal_554, signal_224}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_622, signal_621, signal_620, signal_246}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_231 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_565, signal_564, signal_563, signal_227}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_625, signal_624, signal_623, signal_247}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_232 ( .a ({signal_616, signal_615, signal_614, signal_244}), .b ({signal_628, signal_627, signal_626, signal_248}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_233 ( .a ({signal_619, signal_618, signal_617, signal_245}), .b ({signal_631, signal_630, signal_629, signal_249}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_234 ( .a ({signal_622, signal_621, signal_620, signal_246}), .b ({signal_634, signal_633, signal_632, signal_250}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_235 ( .a ({signal_625, signal_624, signal_623, signal_247}), .b ({signal_637, signal_636, signal_635, signal_251}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_238 ( .a ({1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_601, signal_600, signal_599, signal_239}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_646, signal_645, signal_644, signal_254}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_239 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_598, signal_597, signal_596, signal_238}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_649, signal_648, signal_647, signal_255}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_241 ( .a ({signal_646, signal_645, signal_644, signal_254}), .b ({signal_655, signal_654, signal_653, signal_257}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_242 ( .a ({signal_649, signal_648, signal_647, signal_255}), .b ({signal_658, signal_657, signal_656, signal_258}) ) ;
    buf_clk cell_910 ( .C ( clk ), .D ( signal_2249 ), .Q ( signal_2250 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_911 ( .C ( clk ), .D ( signal_2250 ), .Q ( signal_2251 ) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_227 ( .a ({signal_553, signal_552, signal_551, signal_223}), .b ({signal_517, signal_516, signal_515, signal_211}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_613, signal_612, signal_611, signal_243}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_236 ( .a ({signal_568, signal_567, signal_566, signal_228}), .b ({signal_595, signal_594, signal_593, signal_237}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_640, signal_639, signal_638, signal_252}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_237 ( .a ({signal_607, signal_606, signal_605, signal_241}), .b ({signal_610, signal_609, signal_608, signal_242}), .clk ( clk ), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_643, signal_642, signal_641, signal_253}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_240 ( .a ({signal_643, signal_642, signal_641, signal_253}), .b ({signal_652, signal_651, signal_650, signal_256}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_243 ( .a ({signal_571, signal_570, signal_569, signal_229}), .b ({signal_628, signal_627, signal_626, signal_248}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_661, signal_660, signal_659, signal_259}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_244 ( .a ({signal_604, signal_603, signal_602, signal_240}), .b ({signal_631, signal_630, signal_629, signal_249}), .clk ( clk ), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_664, signal_663, signal_662, signal_260}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_245 ( .a ({signal_520, signal_519, signal_518, signal_212}), .b ({signal_634, signal_633, signal_632, signal_250}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_667, signal_666, signal_665, signal_261}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_246 ( .a ({signal_574, signal_573, signal_572, signal_230}), .b ({signal_637, signal_636, signal_635, signal_251}), .clk ( clk ), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_670, signal_669, signal_668, signal_262}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_247 ( .a ({signal_655, signal_654, signal_653, signal_257}), .b ({signal_658, signal_657, signal_656, signal_258}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_673, signal_672, signal_671, signal_263}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_251 ( .a ({signal_613, signal_612, signal_611, signal_243}), .b ({signal_670, signal_669, signal_668, signal_262}), .c ({signal_685, signal_684, signal_683, signal_267}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_252 ( .a ({signal_640, signal_639, signal_638, signal_252}), .b ({signal_670, signal_669, signal_668, signal_262}), .c ({signal_688, signal_687, signal_686, signal_268}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_253 ( .a ({signal_667, signal_666, signal_665, signal_261}), .b ({signal_643, signal_642, signal_641, signal_253}), .c ({signal_691, signal_690, signal_689, signal_269}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_254 ( .a ({signal_661, signal_660, signal_659, signal_259}), .b ({signal_664, signal_663, signal_662, signal_260}), .c ({signal_694, signal_693, signal_692, signal_270}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_255 ( .a ({signal_664, signal_663, signal_662, signal_260}), .b ({signal_643, signal_642, signal_641, signal_253}), .c ({signal_697, signal_696, signal_695, signal_271}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_256 ( .a ({signal_661, signal_660, signal_659, signal_259}), .b ({signal_667, signal_666, signal_665, signal_261}), .c ({signal_700, signal_699, signal_698, signal_272}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_257 ( .a ({signal_673, signal_672, signal_671, signal_263}), .b ({signal_703, signal_702, signal_701, signal_273}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_258 ( .a ({signal_688, signal_687, signal_686, signal_268}), .b ({signal_706, signal_705, signal_704, signal_274}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_259 ( .a ({signal_691, signal_690, signal_689, signal_269}), .b ({signal_709, signal_708, signal_707, signal_275}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_260 ( .a ({signal_697, signal_696, signal_695, signal_271}), .b ({signal_712, signal_711, signal_710, signal_276}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_261 ( .a ({signal_700, signal_699, signal_698, signal_272}), .b ({signal_715, signal_714, signal_713, signal_277}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_264 ( .a ({signal_640, signal_639, signal_638, signal_252}), .b ({signal_673, signal_672, signal_671, signal_263}), .c ({signal_724, signal_723, signal_722, signal_280}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_265 ( .a ({signal_613, signal_612, signal_611, signal_243}), .b ({signal_673, signal_672, signal_671, signal_263}), .c ({signal_727, signal_726, signal_725, signal_281}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_266 ( .a ({signal_697, signal_696, signal_695, signal_271}), .b ({signal_700, signal_699, signal_698, signal_272}), .c ({signal_730, signal_729, signal_728, signal_282}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_267 ( .a ({signal_724, signal_723, signal_722, signal_280}), .b ({signal_733, signal_732, signal_731, signal_283}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_268 ( .a ({signal_727, signal_726, signal_725, signal_281}), .b ({signal_736, signal_735, signal_734, signal_284}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_273 ( .a ({signal_688, signal_687, signal_686, signal_268}), .b ({signal_727, signal_726, signal_725, signal_281}), .c ({signal_751, signal_750, signal_749, signal_289}) ) ;
    buf_clk cell_912 ( .C ( clk ), .D ( signal_2251 ), .Q ( signal_2252 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_477 ( .C ( clk ), .D ( signal_262 ), .Q ( signal_1817 ) ) ;
    buf_clk cell_483 ( .C ( clk ), .D ( signal_668 ), .Q ( signal_1823 ) ) ;
    buf_clk cell_489 ( .C ( clk ), .D ( signal_669 ), .Q ( signal_1829 ) ) ;
    buf_clk cell_495 ( .C ( clk ), .D ( signal_670 ), .Q ( signal_1835 ) ) ;
    buf_clk cell_501 ( .C ( clk ), .D ( signal_243 ), .Q ( signal_1841 ) ) ;
    buf_clk cell_507 ( .C ( clk ), .D ( signal_611 ), .Q ( signal_1847 ) ) ;
    buf_clk cell_513 ( .C ( clk ), .D ( signal_612 ), .Q ( signal_1853 ) ) ;
    buf_clk cell_519 ( .C ( clk ), .D ( signal_613 ), .Q ( signal_1859 ) ) ;
    buf_clk cell_525 ( .C ( clk ), .D ( signal_252 ), .Q ( signal_1865 ) ) ;
    buf_clk cell_531 ( .C ( clk ), .D ( signal_638 ), .Q ( signal_1871 ) ) ;
    buf_clk cell_537 ( .C ( clk ), .D ( signal_639 ), .Q ( signal_1877 ) ) ;
    buf_clk cell_543 ( .C ( clk ), .D ( signal_640 ), .Q ( signal_1883 ) ) ;
    buf_clk cell_549 ( .C ( clk ), .D ( signal_263 ), .Q ( signal_1889 ) ) ;
    buf_clk cell_555 ( .C ( clk ), .D ( signal_671 ), .Q ( signal_1895 ) ) ;
    buf_clk cell_561 ( .C ( clk ), .D ( signal_672 ), .Q ( signal_1901 ) ) ;
    buf_clk cell_567 ( .C ( clk ), .D ( signal_673 ), .Q ( signal_1907 ) ) ;
    buf_clk cell_573 ( .C ( clk ), .D ( signal_259 ), .Q ( signal_1913 ) ) ;
    buf_clk cell_579 ( .C ( clk ), .D ( signal_659 ), .Q ( signal_1919 ) ) ;
    buf_clk cell_585 ( .C ( clk ), .D ( signal_660 ), .Q ( signal_1925 ) ) ;
    buf_clk cell_591 ( .C ( clk ), .D ( signal_661 ), .Q ( signal_1931 ) ) ;
    buf_clk cell_597 ( .C ( clk ), .D ( signal_260 ), .Q ( signal_1937 ) ) ;
    buf_clk cell_603 ( .C ( clk ), .D ( signal_662 ), .Q ( signal_1943 ) ) ;
    buf_clk cell_609 ( .C ( clk ), .D ( signal_663 ), .Q ( signal_1949 ) ) ;
    buf_clk cell_615 ( .C ( clk ), .D ( signal_664 ), .Q ( signal_1955 ) ) ;
    buf_clk cell_621 ( .C ( clk ), .D ( signal_261 ), .Q ( signal_1961 ) ) ;
    buf_clk cell_627 ( .C ( clk ), .D ( signal_665 ), .Q ( signal_1967 ) ) ;
    buf_clk cell_633 ( .C ( clk ), .D ( signal_666 ), .Q ( signal_1973 ) ) ;
    buf_clk cell_639 ( .C ( clk ), .D ( signal_667 ), .Q ( signal_1979 ) ) ;
    buf_clk cell_645 ( .C ( clk ), .D ( signal_253 ), .Q ( signal_1985 ) ) ;
    buf_clk cell_651 ( .C ( clk ), .D ( signal_641 ), .Q ( signal_1991 ) ) ;
    buf_clk cell_657 ( .C ( clk ), .D ( signal_642 ), .Q ( signal_1997 ) ) ;
    buf_clk cell_663 ( .C ( clk ), .D ( signal_643 ), .Q ( signal_2003 ) ) ;
    buf_clk cell_669 ( .C ( clk ), .D ( signal_267 ), .Q ( signal_2009 ) ) ;
    buf_clk cell_675 ( .C ( clk ), .D ( signal_683 ), .Q ( signal_2015 ) ) ;
    buf_clk cell_681 ( .C ( clk ), .D ( signal_684 ), .Q ( signal_2021 ) ) ;
    buf_clk cell_687 ( .C ( clk ), .D ( signal_685 ), .Q ( signal_2027 ) ) ;
    buf_clk cell_693 ( .C ( clk ), .D ( signal_280 ), .Q ( signal_2033 ) ) ;
    buf_clk cell_699 ( .C ( clk ), .D ( signal_722 ), .Q ( signal_2039 ) ) ;
    buf_clk cell_705 ( .C ( clk ), .D ( signal_723 ), .Q ( signal_2045 ) ) ;
    buf_clk cell_711 ( .C ( clk ), .D ( signal_724 ), .Q ( signal_2051 ) ) ;
    buf_clk cell_717 ( .C ( clk ), .D ( signal_268 ), .Q ( signal_2057 ) ) ;
    buf_clk cell_723 ( .C ( clk ), .D ( signal_686 ), .Q ( signal_2063 ) ) ;
    buf_clk cell_729 ( .C ( clk ), .D ( signal_687 ), .Q ( signal_2069 ) ) ;
    buf_clk cell_735 ( .C ( clk ), .D ( signal_688 ), .Q ( signal_2075 ) ) ;
    buf_clk cell_741 ( .C ( clk ), .D ( signal_281 ), .Q ( signal_2081 ) ) ;
    buf_clk cell_747 ( .C ( clk ), .D ( signal_725 ), .Q ( signal_2087 ) ) ;
    buf_clk cell_753 ( .C ( clk ), .D ( signal_726 ), .Q ( signal_2093 ) ) ;
    buf_clk cell_759 ( .C ( clk ), .D ( signal_727 ), .Q ( signal_2099 ) ) ;
    buf_clk cell_765 ( .C ( clk ), .D ( signal_270 ), .Q ( signal_2105 ) ) ;
    buf_clk cell_771 ( .C ( clk ), .D ( signal_692 ), .Q ( signal_2111 ) ) ;
    buf_clk cell_777 ( .C ( clk ), .D ( signal_693 ), .Q ( signal_2117 ) ) ;
    buf_clk cell_783 ( .C ( clk ), .D ( signal_694 ), .Q ( signal_2123 ) ) ;
    buf_clk cell_789 ( .C ( clk ), .D ( signal_269 ), .Q ( signal_2129 ) ) ;
    buf_clk cell_795 ( .C ( clk ), .D ( signal_689 ), .Q ( signal_2135 ) ) ;
    buf_clk cell_801 ( .C ( clk ), .D ( signal_690 ), .Q ( signal_2141 ) ) ;
    buf_clk cell_807 ( .C ( clk ), .D ( signal_691 ), .Q ( signal_2147 ) ) ;
    buf_clk cell_813 ( .C ( clk ), .D ( signal_272 ), .Q ( signal_2153 ) ) ;
    buf_clk cell_819 ( .C ( clk ), .D ( signal_698 ), .Q ( signal_2159 ) ) ;
    buf_clk cell_825 ( .C ( clk ), .D ( signal_699 ), .Q ( signal_2165 ) ) ;
    buf_clk cell_831 ( .C ( clk ), .D ( signal_700 ), .Q ( signal_2171 ) ) ;
    buf_clk cell_837 ( .C ( clk ), .D ( signal_271 ), .Q ( signal_2177 ) ) ;
    buf_clk cell_843 ( .C ( clk ), .D ( signal_695 ), .Q ( signal_2183 ) ) ;
    buf_clk cell_849 ( .C ( clk ), .D ( signal_696 ), .Q ( signal_2189 ) ) ;
    buf_clk cell_855 ( .C ( clk ), .D ( signal_697 ), .Q ( signal_2195 ) ) ;
    buf_clk cell_861 ( .C ( clk ), .D ( signal_289 ), .Q ( signal_2201 ) ) ;
    buf_clk cell_867 ( .C ( clk ), .D ( signal_749 ), .Q ( signal_2207 ) ) ;
    buf_clk cell_873 ( .C ( clk ), .D ( signal_750 ), .Q ( signal_2213 ) ) ;
    buf_clk cell_879 ( .C ( clk ), .D ( signal_751 ), .Q ( signal_2219 ) ) ;
    buf_clk cell_885 ( .C ( clk ), .D ( signal_282 ), .Q ( signal_2225 ) ) ;
    buf_clk cell_891 ( .C ( clk ), .D ( signal_728 ), .Q ( signal_2231 ) ) ;
    buf_clk cell_897 ( .C ( clk ), .D ( signal_729 ), .Q ( signal_2237 ) ) ;
    buf_clk cell_903 ( .C ( clk ), .D ( signal_730 ), .Q ( signal_2243 ) ) ;
    buf_clk cell_913 ( .C ( clk ), .D ( signal_2252 ), .Q ( signal_2253 ) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_248 ( .a ({signal_661, signal_660, signal_659, signal_259}), .b ({signal_670, signal_669, signal_668, signal_262}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_676, signal_675, signal_674, signal_264}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_249 ( .a ({signal_613, signal_612, signal_611, signal_243}), .b ({signal_664, signal_663, signal_662, signal_260}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_679, signal_678, signal_677, signal_265}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_250 ( .a ({signal_640, signal_639, signal_638, signal_252}), .b ({signal_667, signal_666, signal_665, signal_261}), .clk ( clk ), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_682, signal_681, signal_680, signal_266}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_262 ( .a ({signal_685, signal_684, signal_683, signal_267}), .b ({signal_694, signal_693, signal_692, signal_270}), .clk ( clk ), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_718, signal_717, signal_716, signal_278}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_263 ( .a ({signal_688, signal_687, signal_686, signal_268}), .b ({signal_700, signal_699, signal_698, signal_272}), .clk ( clk ), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_721, signal_720, signal_719, signal_279}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_269 ( .a ({signal_706, signal_705, signal_704, signal_274}), .b ({signal_715, signal_714, signal_713, signal_277}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_739, signal_738, signal_737, signal_285}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_270 ( .a ({signal_652, signal_651, signal_650, signal_256}), .b ({signal_703, signal_702, signal_701, signal_273}), .clk ( clk ), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_742, signal_741, signal_740, signal_286}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_271 ( .a ({signal_691, signal_690, signal_689, signal_269}), .b ({signal_724, signal_723, signal_722, signal_280}), .clk ( clk ), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_745, signal_744, signal_743, signal_287}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_272 ( .a ({signal_697, signal_696, signal_695, signal_271}), .b ({signal_727, signal_726, signal_725, signal_281}), .clk ( clk ), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_748, signal_747, signal_746, signal_288}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_274 ( .a ({signal_712, signal_711, signal_710, signal_276}), .b ({signal_736, signal_735, signal_734, signal_284}), .clk ( clk ), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_754, signal_753, signal_752, signal_290}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_275 ( .a ({signal_709, signal_708, signal_707, signal_275}), .b ({signal_733, signal_732, signal_731, signal_283}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({signal_757, signal_756, signal_755, signal_291}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_276 ( .a ({signal_730, signal_729, signal_728, signal_282}), .b ({signal_751, signal_750, signal_749, signal_289}), .clk ( clk ), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_760, signal_759, signal_758, signal_292}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_277 ( .a ({signal_679, signal_678, signal_677, signal_265}), .b ({signal_739, signal_738, signal_737, signal_285}), .c ({signal_763, signal_762, signal_761, signal_293}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_278 ( .a ({signal_718, signal_717, signal_716, signal_278}), .b ({signal_748, signal_747, signal_746, signal_288}), .c ({signal_766, signal_765, signal_764, signal_294}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_279 ( .a ({signal_742, signal_741, signal_740, signal_286}), .b ({signal_745, signal_744, signal_743, signal_287}), .c ({signal_769, signal_768, signal_767, signal_295}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_280 ( .a ({signal_676, signal_675, signal_674, signal_264}), .b ({signal_754, signal_753, signal_752, signal_290}), .c ({signal_772, signal_771, signal_770, signal_296}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_281 ( .a ({signal_682, signal_681, signal_680, signal_266}), .b ({signal_757, signal_756, signal_755, signal_291}), .c ({signal_775, signal_774, signal_773, signal_297}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_282 ( .a ({signal_718, signal_717, signal_716, signal_278}), .b ({signal_760, signal_759, signal_758, signal_292}), .c ({signal_778, signal_777, signal_776, signal_298}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_283 ( .a ({signal_763, signal_762, signal_761, signal_293}), .b ({signal_766, signal_765, signal_764, signal_294}), .c ({signal_781, signal_780, signal_779, signal_299}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_284 ( .a ({signal_748, signal_747, signal_746, signal_288}), .b ({signal_760, signal_759, signal_758, signal_292}), .c ({signal_784, signal_783, signal_782, signal_300}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_285 ( .a ({signal_721, signal_720, signal_719, signal_279}), .b ({signal_769, signal_768, signal_767, signal_295}), .c ({signal_787, signal_786, signal_785, signal_301}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_286 ( .a ({signal_781, signal_780, signal_779, signal_299}), .b ({signal_790, signal_789, signal_788, signal_302}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_287 ( .a ({signal_772, signal_771, signal_770, signal_296}), .b ({signal_778, signal_777, signal_776, signal_298}), .c ({signal_793, signal_792, signal_791, signal_303}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_288 ( .a ({signal_775, signal_774, signal_773, signal_297}), .b ({signal_784, signal_783, signal_782, signal_300}), .c ({signal_796, signal_795, signal_794, signal_304}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_289 ( .a ({signal_748, signal_747, signal_746, signal_288}), .b ({signal_787, signal_786, signal_785, signal_301}), .c ({signal_799, signal_798, signal_797, signal_305}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_290 ( .a ({signal_793, signal_792, signal_791, signal_303}), .b ({signal_802, signal_801, signal_800, signal_306}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_291 ( .a ({signal_796, signal_795, signal_794, signal_304}), .b ({signal_805, signal_804, signal_803, signal_307}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_292 ( .a ({signal_799, signal_798, signal_797, signal_305}), .b ({signal_808, signal_807, signal_806, signal_308}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_294 ( .a ({signal_781, signal_780, signal_779, signal_299}), .b ({signal_793, signal_792, signal_791, signal_303}), .c ({signal_814, signal_813, signal_812, signal_310}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_295 ( .a ({signal_796, signal_795, signal_794, signal_304}), .b ({signal_799, signal_798, signal_797, signal_305}), .c ({signal_817, signal_816, signal_815, signal_311}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_296 ( .a ({signal_814, signal_813, signal_812, signal_310}), .b ({signal_820, signal_819, signal_818, signal_312}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_297 ( .a ({signal_817, signal_816, signal_815, signal_311}), .b ({signal_823, signal_822, signal_821, signal_313}) ) ;
    buf_clk cell_478 ( .C ( clk ), .D ( signal_1817 ), .Q ( signal_1818 ) ) ;
    buf_clk cell_484 ( .C ( clk ), .D ( signal_1823 ), .Q ( signal_1824 ) ) ;
    buf_clk cell_490 ( .C ( clk ), .D ( signal_1829 ), .Q ( signal_1830 ) ) ;
    buf_clk cell_496 ( .C ( clk ), .D ( signal_1835 ), .Q ( signal_1836 ) ) ;
    buf_clk cell_502 ( .C ( clk ), .D ( signal_1841 ), .Q ( signal_1842 ) ) ;
    buf_clk cell_508 ( .C ( clk ), .D ( signal_1847 ), .Q ( signal_1848 ) ) ;
    buf_clk cell_514 ( .C ( clk ), .D ( signal_1853 ), .Q ( signal_1854 ) ) ;
    buf_clk cell_520 ( .C ( clk ), .D ( signal_1859 ), .Q ( signal_1860 ) ) ;
    buf_clk cell_526 ( .C ( clk ), .D ( signal_1865 ), .Q ( signal_1866 ) ) ;
    buf_clk cell_532 ( .C ( clk ), .D ( signal_1871 ), .Q ( signal_1872 ) ) ;
    buf_clk cell_538 ( .C ( clk ), .D ( signal_1877 ), .Q ( signal_1878 ) ) ;
    buf_clk cell_544 ( .C ( clk ), .D ( signal_1883 ), .Q ( signal_1884 ) ) ;
    buf_clk cell_550 ( .C ( clk ), .D ( signal_1889 ), .Q ( signal_1890 ) ) ;
    buf_clk cell_556 ( .C ( clk ), .D ( signal_1895 ), .Q ( signal_1896 ) ) ;
    buf_clk cell_562 ( .C ( clk ), .D ( signal_1901 ), .Q ( signal_1902 ) ) ;
    buf_clk cell_568 ( .C ( clk ), .D ( signal_1907 ), .Q ( signal_1908 ) ) ;
    buf_clk cell_574 ( .C ( clk ), .D ( signal_1913 ), .Q ( signal_1914 ) ) ;
    buf_clk cell_580 ( .C ( clk ), .D ( signal_1919 ), .Q ( signal_1920 ) ) ;
    buf_clk cell_586 ( .C ( clk ), .D ( signal_1925 ), .Q ( signal_1926 ) ) ;
    buf_clk cell_592 ( .C ( clk ), .D ( signal_1931 ), .Q ( signal_1932 ) ) ;
    buf_clk cell_598 ( .C ( clk ), .D ( signal_1937 ), .Q ( signal_1938 ) ) ;
    buf_clk cell_604 ( .C ( clk ), .D ( signal_1943 ), .Q ( signal_1944 ) ) ;
    buf_clk cell_610 ( .C ( clk ), .D ( signal_1949 ), .Q ( signal_1950 ) ) ;
    buf_clk cell_616 ( .C ( clk ), .D ( signal_1955 ), .Q ( signal_1956 ) ) ;
    buf_clk cell_622 ( .C ( clk ), .D ( signal_1961 ), .Q ( signal_1962 ) ) ;
    buf_clk cell_628 ( .C ( clk ), .D ( signal_1967 ), .Q ( signal_1968 ) ) ;
    buf_clk cell_634 ( .C ( clk ), .D ( signal_1973 ), .Q ( signal_1974 ) ) ;
    buf_clk cell_640 ( .C ( clk ), .D ( signal_1979 ), .Q ( signal_1980 ) ) ;
    buf_clk cell_646 ( .C ( clk ), .D ( signal_1985 ), .Q ( signal_1986 ) ) ;
    buf_clk cell_652 ( .C ( clk ), .D ( signal_1991 ), .Q ( signal_1992 ) ) ;
    buf_clk cell_658 ( .C ( clk ), .D ( signal_1997 ), .Q ( signal_1998 ) ) ;
    buf_clk cell_664 ( .C ( clk ), .D ( signal_2003 ), .Q ( signal_2004 ) ) ;
    buf_clk cell_670 ( .C ( clk ), .D ( signal_2009 ), .Q ( signal_2010 ) ) ;
    buf_clk cell_676 ( .C ( clk ), .D ( signal_2015 ), .Q ( signal_2016 ) ) ;
    buf_clk cell_682 ( .C ( clk ), .D ( signal_2021 ), .Q ( signal_2022 ) ) ;
    buf_clk cell_688 ( .C ( clk ), .D ( signal_2027 ), .Q ( signal_2028 ) ) ;
    buf_clk cell_694 ( .C ( clk ), .D ( signal_2033 ), .Q ( signal_2034 ) ) ;
    buf_clk cell_700 ( .C ( clk ), .D ( signal_2039 ), .Q ( signal_2040 ) ) ;
    buf_clk cell_706 ( .C ( clk ), .D ( signal_2045 ), .Q ( signal_2046 ) ) ;
    buf_clk cell_712 ( .C ( clk ), .D ( signal_2051 ), .Q ( signal_2052 ) ) ;
    buf_clk cell_718 ( .C ( clk ), .D ( signal_2057 ), .Q ( signal_2058 ) ) ;
    buf_clk cell_724 ( .C ( clk ), .D ( signal_2063 ), .Q ( signal_2064 ) ) ;
    buf_clk cell_730 ( .C ( clk ), .D ( signal_2069 ), .Q ( signal_2070 ) ) ;
    buf_clk cell_736 ( .C ( clk ), .D ( signal_2075 ), .Q ( signal_2076 ) ) ;
    buf_clk cell_742 ( .C ( clk ), .D ( signal_2081 ), .Q ( signal_2082 ) ) ;
    buf_clk cell_748 ( .C ( clk ), .D ( signal_2087 ), .Q ( signal_2088 ) ) ;
    buf_clk cell_754 ( .C ( clk ), .D ( signal_2093 ), .Q ( signal_2094 ) ) ;
    buf_clk cell_760 ( .C ( clk ), .D ( signal_2099 ), .Q ( signal_2100 ) ) ;
    buf_clk cell_766 ( .C ( clk ), .D ( signal_2105 ), .Q ( signal_2106 ) ) ;
    buf_clk cell_772 ( .C ( clk ), .D ( signal_2111 ), .Q ( signal_2112 ) ) ;
    buf_clk cell_778 ( .C ( clk ), .D ( signal_2117 ), .Q ( signal_2118 ) ) ;
    buf_clk cell_784 ( .C ( clk ), .D ( signal_2123 ), .Q ( signal_2124 ) ) ;
    buf_clk cell_790 ( .C ( clk ), .D ( signal_2129 ), .Q ( signal_2130 ) ) ;
    buf_clk cell_796 ( .C ( clk ), .D ( signal_2135 ), .Q ( signal_2136 ) ) ;
    buf_clk cell_802 ( .C ( clk ), .D ( signal_2141 ), .Q ( signal_2142 ) ) ;
    buf_clk cell_808 ( .C ( clk ), .D ( signal_2147 ), .Q ( signal_2148 ) ) ;
    buf_clk cell_814 ( .C ( clk ), .D ( signal_2153 ), .Q ( signal_2154 ) ) ;
    buf_clk cell_820 ( .C ( clk ), .D ( signal_2159 ), .Q ( signal_2160 ) ) ;
    buf_clk cell_826 ( .C ( clk ), .D ( signal_2165 ), .Q ( signal_2166 ) ) ;
    buf_clk cell_832 ( .C ( clk ), .D ( signal_2171 ), .Q ( signal_2172 ) ) ;
    buf_clk cell_838 ( .C ( clk ), .D ( signal_2177 ), .Q ( signal_2178 ) ) ;
    buf_clk cell_844 ( .C ( clk ), .D ( signal_2183 ), .Q ( signal_2184 ) ) ;
    buf_clk cell_850 ( .C ( clk ), .D ( signal_2189 ), .Q ( signal_2190 ) ) ;
    buf_clk cell_856 ( .C ( clk ), .D ( signal_2195 ), .Q ( signal_2196 ) ) ;
    buf_clk cell_862 ( .C ( clk ), .D ( signal_2201 ), .Q ( signal_2202 ) ) ;
    buf_clk cell_868 ( .C ( clk ), .D ( signal_2207 ), .Q ( signal_2208 ) ) ;
    buf_clk cell_874 ( .C ( clk ), .D ( signal_2213 ), .Q ( signal_2214 ) ) ;
    buf_clk cell_880 ( .C ( clk ), .D ( signal_2219 ), .Q ( signal_2220 ) ) ;
    buf_clk cell_886 ( .C ( clk ), .D ( signal_2225 ), .Q ( signal_2226 ) ) ;
    buf_clk cell_892 ( .C ( clk ), .D ( signal_2231 ), .Q ( signal_2232 ) ) ;
    buf_clk cell_898 ( .C ( clk ), .D ( signal_2237 ), .Q ( signal_2238 ) ) ;
    buf_clk cell_904 ( .C ( clk ), .D ( signal_2243 ), .Q ( signal_2244 ) ) ;
    buf_clk cell_914 ( .C ( clk ), .D ( signal_2253 ), .Q ( signal_2254 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_429 ( .C ( clk ), .D ( signal_308 ), .Q ( signal_1769 ) ) ;
    buf_clk cell_431 ( .C ( clk ), .D ( signal_806 ), .Q ( signal_1771 ) ) ;
    buf_clk cell_433 ( .C ( clk ), .D ( signal_807 ), .Q ( signal_1773 ) ) ;
    buf_clk cell_435 ( .C ( clk ), .D ( signal_808 ), .Q ( signal_1775 ) ) ;
    buf_clk cell_437 ( .C ( clk ), .D ( signal_302 ), .Q ( signal_1777 ) ) ;
    buf_clk cell_439 ( .C ( clk ), .D ( signal_788 ), .Q ( signal_1779 ) ) ;
    buf_clk cell_441 ( .C ( clk ), .D ( signal_789 ), .Q ( signal_1781 ) ) ;
    buf_clk cell_443 ( .C ( clk ), .D ( signal_790 ), .Q ( signal_1783 ) ) ;
    buf_clk cell_445 ( .C ( clk ), .D ( signal_307 ), .Q ( signal_1785 ) ) ;
    buf_clk cell_447 ( .C ( clk ), .D ( signal_803 ), .Q ( signal_1787 ) ) ;
    buf_clk cell_449 ( .C ( clk ), .D ( signal_804 ), .Q ( signal_1789 ) ) ;
    buf_clk cell_451 ( .C ( clk ), .D ( signal_805 ), .Q ( signal_1791 ) ) ;
    buf_clk cell_453 ( .C ( clk ), .D ( signal_306 ), .Q ( signal_1793 ) ) ;
    buf_clk cell_455 ( .C ( clk ), .D ( signal_800 ), .Q ( signal_1795 ) ) ;
    buf_clk cell_457 ( .C ( clk ), .D ( signal_801 ), .Q ( signal_1797 ) ) ;
    buf_clk cell_459 ( .C ( clk ), .D ( signal_802 ), .Q ( signal_1799 ) ) ;
    buf_clk cell_461 ( .C ( clk ), .D ( signal_311 ), .Q ( signal_1801 ) ) ;
    buf_clk cell_463 ( .C ( clk ), .D ( signal_815 ), .Q ( signal_1803 ) ) ;
    buf_clk cell_465 ( .C ( clk ), .D ( signal_816 ), .Q ( signal_1805 ) ) ;
    buf_clk cell_467 ( .C ( clk ), .D ( signal_817 ), .Q ( signal_1807 ) ) ;
    buf_clk cell_469 ( .C ( clk ), .D ( signal_310 ), .Q ( signal_1809 ) ) ;
    buf_clk cell_471 ( .C ( clk ), .D ( signal_812 ), .Q ( signal_1811 ) ) ;
    buf_clk cell_473 ( .C ( clk ), .D ( signal_813 ), .Q ( signal_1813 ) ) ;
    buf_clk cell_475 ( .C ( clk ), .D ( signal_814 ), .Q ( signal_1815 ) ) ;
    buf_clk cell_479 ( .C ( clk ), .D ( signal_1818 ), .Q ( signal_1819 ) ) ;
    buf_clk cell_485 ( .C ( clk ), .D ( signal_1824 ), .Q ( signal_1825 ) ) ;
    buf_clk cell_491 ( .C ( clk ), .D ( signal_1830 ), .Q ( signal_1831 ) ) ;
    buf_clk cell_497 ( .C ( clk ), .D ( signal_1836 ), .Q ( signal_1837 ) ) ;
    buf_clk cell_503 ( .C ( clk ), .D ( signal_1842 ), .Q ( signal_1843 ) ) ;
    buf_clk cell_509 ( .C ( clk ), .D ( signal_1848 ), .Q ( signal_1849 ) ) ;
    buf_clk cell_515 ( .C ( clk ), .D ( signal_1854 ), .Q ( signal_1855 ) ) ;
    buf_clk cell_521 ( .C ( clk ), .D ( signal_1860 ), .Q ( signal_1861 ) ) ;
    buf_clk cell_527 ( .C ( clk ), .D ( signal_1866 ), .Q ( signal_1867 ) ) ;
    buf_clk cell_533 ( .C ( clk ), .D ( signal_1872 ), .Q ( signal_1873 ) ) ;
    buf_clk cell_539 ( .C ( clk ), .D ( signal_1878 ), .Q ( signal_1879 ) ) ;
    buf_clk cell_545 ( .C ( clk ), .D ( signal_1884 ), .Q ( signal_1885 ) ) ;
    buf_clk cell_551 ( .C ( clk ), .D ( signal_1890 ), .Q ( signal_1891 ) ) ;
    buf_clk cell_557 ( .C ( clk ), .D ( signal_1896 ), .Q ( signal_1897 ) ) ;
    buf_clk cell_563 ( .C ( clk ), .D ( signal_1902 ), .Q ( signal_1903 ) ) ;
    buf_clk cell_569 ( .C ( clk ), .D ( signal_1908 ), .Q ( signal_1909 ) ) ;
    buf_clk cell_575 ( .C ( clk ), .D ( signal_1914 ), .Q ( signal_1915 ) ) ;
    buf_clk cell_581 ( .C ( clk ), .D ( signal_1920 ), .Q ( signal_1921 ) ) ;
    buf_clk cell_587 ( .C ( clk ), .D ( signal_1926 ), .Q ( signal_1927 ) ) ;
    buf_clk cell_593 ( .C ( clk ), .D ( signal_1932 ), .Q ( signal_1933 ) ) ;
    buf_clk cell_599 ( .C ( clk ), .D ( signal_1938 ), .Q ( signal_1939 ) ) ;
    buf_clk cell_605 ( .C ( clk ), .D ( signal_1944 ), .Q ( signal_1945 ) ) ;
    buf_clk cell_611 ( .C ( clk ), .D ( signal_1950 ), .Q ( signal_1951 ) ) ;
    buf_clk cell_617 ( .C ( clk ), .D ( signal_1956 ), .Q ( signal_1957 ) ) ;
    buf_clk cell_623 ( .C ( clk ), .D ( signal_1962 ), .Q ( signal_1963 ) ) ;
    buf_clk cell_629 ( .C ( clk ), .D ( signal_1968 ), .Q ( signal_1969 ) ) ;
    buf_clk cell_635 ( .C ( clk ), .D ( signal_1974 ), .Q ( signal_1975 ) ) ;
    buf_clk cell_641 ( .C ( clk ), .D ( signal_1980 ), .Q ( signal_1981 ) ) ;
    buf_clk cell_647 ( .C ( clk ), .D ( signal_1986 ), .Q ( signal_1987 ) ) ;
    buf_clk cell_653 ( .C ( clk ), .D ( signal_1992 ), .Q ( signal_1993 ) ) ;
    buf_clk cell_659 ( .C ( clk ), .D ( signal_1998 ), .Q ( signal_1999 ) ) ;
    buf_clk cell_665 ( .C ( clk ), .D ( signal_2004 ), .Q ( signal_2005 ) ) ;
    buf_clk cell_671 ( .C ( clk ), .D ( signal_2010 ), .Q ( signal_2011 ) ) ;
    buf_clk cell_677 ( .C ( clk ), .D ( signal_2016 ), .Q ( signal_2017 ) ) ;
    buf_clk cell_683 ( .C ( clk ), .D ( signal_2022 ), .Q ( signal_2023 ) ) ;
    buf_clk cell_689 ( .C ( clk ), .D ( signal_2028 ), .Q ( signal_2029 ) ) ;
    buf_clk cell_695 ( .C ( clk ), .D ( signal_2034 ), .Q ( signal_2035 ) ) ;
    buf_clk cell_701 ( .C ( clk ), .D ( signal_2040 ), .Q ( signal_2041 ) ) ;
    buf_clk cell_707 ( .C ( clk ), .D ( signal_2046 ), .Q ( signal_2047 ) ) ;
    buf_clk cell_713 ( .C ( clk ), .D ( signal_2052 ), .Q ( signal_2053 ) ) ;
    buf_clk cell_719 ( .C ( clk ), .D ( signal_2058 ), .Q ( signal_2059 ) ) ;
    buf_clk cell_725 ( .C ( clk ), .D ( signal_2064 ), .Q ( signal_2065 ) ) ;
    buf_clk cell_731 ( .C ( clk ), .D ( signal_2070 ), .Q ( signal_2071 ) ) ;
    buf_clk cell_737 ( .C ( clk ), .D ( signal_2076 ), .Q ( signal_2077 ) ) ;
    buf_clk cell_743 ( .C ( clk ), .D ( signal_2082 ), .Q ( signal_2083 ) ) ;
    buf_clk cell_749 ( .C ( clk ), .D ( signal_2088 ), .Q ( signal_2089 ) ) ;
    buf_clk cell_755 ( .C ( clk ), .D ( signal_2094 ), .Q ( signal_2095 ) ) ;
    buf_clk cell_761 ( .C ( clk ), .D ( signal_2100 ), .Q ( signal_2101 ) ) ;
    buf_clk cell_767 ( .C ( clk ), .D ( signal_2106 ), .Q ( signal_2107 ) ) ;
    buf_clk cell_773 ( .C ( clk ), .D ( signal_2112 ), .Q ( signal_2113 ) ) ;
    buf_clk cell_779 ( .C ( clk ), .D ( signal_2118 ), .Q ( signal_2119 ) ) ;
    buf_clk cell_785 ( .C ( clk ), .D ( signal_2124 ), .Q ( signal_2125 ) ) ;
    buf_clk cell_791 ( .C ( clk ), .D ( signal_2130 ), .Q ( signal_2131 ) ) ;
    buf_clk cell_797 ( .C ( clk ), .D ( signal_2136 ), .Q ( signal_2137 ) ) ;
    buf_clk cell_803 ( .C ( clk ), .D ( signal_2142 ), .Q ( signal_2143 ) ) ;
    buf_clk cell_809 ( .C ( clk ), .D ( signal_2148 ), .Q ( signal_2149 ) ) ;
    buf_clk cell_815 ( .C ( clk ), .D ( signal_2154 ), .Q ( signal_2155 ) ) ;
    buf_clk cell_821 ( .C ( clk ), .D ( signal_2160 ), .Q ( signal_2161 ) ) ;
    buf_clk cell_827 ( .C ( clk ), .D ( signal_2166 ), .Q ( signal_2167 ) ) ;
    buf_clk cell_833 ( .C ( clk ), .D ( signal_2172 ), .Q ( signal_2173 ) ) ;
    buf_clk cell_839 ( .C ( clk ), .D ( signal_2178 ), .Q ( signal_2179 ) ) ;
    buf_clk cell_845 ( .C ( clk ), .D ( signal_2184 ), .Q ( signal_2185 ) ) ;
    buf_clk cell_851 ( .C ( clk ), .D ( signal_2190 ), .Q ( signal_2191 ) ) ;
    buf_clk cell_857 ( .C ( clk ), .D ( signal_2196 ), .Q ( signal_2197 ) ) ;
    buf_clk cell_863 ( .C ( clk ), .D ( signal_2202 ), .Q ( signal_2203 ) ) ;
    buf_clk cell_869 ( .C ( clk ), .D ( signal_2208 ), .Q ( signal_2209 ) ) ;
    buf_clk cell_875 ( .C ( clk ), .D ( signal_2214 ), .Q ( signal_2215 ) ) ;
    buf_clk cell_881 ( .C ( clk ), .D ( signal_2220 ), .Q ( signal_2221 ) ) ;
    buf_clk cell_887 ( .C ( clk ), .D ( signal_2226 ), .Q ( signal_2227 ) ) ;
    buf_clk cell_893 ( .C ( clk ), .D ( signal_2232 ), .Q ( signal_2233 ) ) ;
    buf_clk cell_899 ( .C ( clk ), .D ( signal_2238 ), .Q ( signal_2239 ) ) ;
    buf_clk cell_905 ( .C ( clk ), .D ( signal_2244 ), .Q ( signal_2245 ) ) ;
    buf_clk cell_915 ( .C ( clk ), .D ( signal_2254 ), .Q ( signal_2255 ) ) ;

    /* cells in depth 8 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_293 ( .a ({signal_793, signal_792, signal_791, signal_303}), .b ({signal_796, signal_795, signal_794, signal_304}), .clk ( clk ), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({signal_811, signal_810, signal_809, signal_309}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_298 ( .a ({signal_790, signal_789, signal_788, signal_302}), .b ({signal_808, signal_807, signal_806, signal_308}), .clk ( clk ), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({signal_826, signal_825, signal_824, signal_314}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_299 ( .a ({signal_814, signal_813, signal_812, signal_310}), .b ({signal_817, signal_816, signal_815, signal_311}), .clk ( clk ), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({signal_829, signal_828, signal_827, signal_315}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_300 ( .a ({signal_820, signal_819, signal_818, signal_312}), .b ({signal_823, signal_822, signal_821, signal_313}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({signal_832, signal_831, signal_830, signal_316}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_301 ( .a ({signal_811, signal_810, signal_809, signal_309}), .b ({signal_829, signal_828, signal_827, signal_315}), .c ({signal_835, signal_834, signal_833, signal_317}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_302 ( .a ({signal_835, signal_834, signal_833, signal_317}), .b ({signal_838, signal_837, signal_836, signal_318}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_303 ( .a ({signal_826, signal_825, signal_824, signal_314}), .b ({signal_832, signal_831, signal_830, signal_316}), .c ({signal_841, signal_840, signal_839, signal_319}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_304 ( .a ({signal_841, signal_840, signal_839, signal_319}), .b ({signal_844, signal_843, signal_842, signal_320}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_307 ( .a ({signal_835, signal_834, signal_833, signal_317}), .b ({signal_841, signal_840, signal_839, signal_319}), .c ({signal_853, signal_852, signal_851, signal_323}) ) ;
    buf_clk cell_430 ( .C ( clk ), .D ( signal_1769 ), .Q ( signal_1770 ) ) ;
    buf_clk cell_432 ( .C ( clk ), .D ( signal_1771 ), .Q ( signal_1772 ) ) ;
    buf_clk cell_434 ( .C ( clk ), .D ( signal_1773 ), .Q ( signal_1774 ) ) ;
    buf_clk cell_436 ( .C ( clk ), .D ( signal_1775 ), .Q ( signal_1776 ) ) ;
    buf_clk cell_438 ( .C ( clk ), .D ( signal_1777 ), .Q ( signal_1778 ) ) ;
    buf_clk cell_440 ( .C ( clk ), .D ( signal_1779 ), .Q ( signal_1780 ) ) ;
    buf_clk cell_442 ( .C ( clk ), .D ( signal_1781 ), .Q ( signal_1782 ) ) ;
    buf_clk cell_444 ( .C ( clk ), .D ( signal_1783 ), .Q ( signal_1784 ) ) ;
    buf_clk cell_446 ( .C ( clk ), .D ( signal_1785 ), .Q ( signal_1786 ) ) ;
    buf_clk cell_448 ( .C ( clk ), .D ( signal_1787 ), .Q ( signal_1788 ) ) ;
    buf_clk cell_450 ( .C ( clk ), .D ( signal_1789 ), .Q ( signal_1790 ) ) ;
    buf_clk cell_452 ( .C ( clk ), .D ( signal_1791 ), .Q ( signal_1792 ) ) ;
    buf_clk cell_454 ( .C ( clk ), .D ( signal_1793 ), .Q ( signal_1794 ) ) ;
    buf_clk cell_456 ( .C ( clk ), .D ( signal_1795 ), .Q ( signal_1796 ) ) ;
    buf_clk cell_458 ( .C ( clk ), .D ( signal_1797 ), .Q ( signal_1798 ) ) ;
    buf_clk cell_460 ( .C ( clk ), .D ( signal_1799 ), .Q ( signal_1800 ) ) ;
    buf_clk cell_462 ( .C ( clk ), .D ( signal_1801 ), .Q ( signal_1802 ) ) ;
    buf_clk cell_464 ( .C ( clk ), .D ( signal_1803 ), .Q ( signal_1804 ) ) ;
    buf_clk cell_466 ( .C ( clk ), .D ( signal_1805 ), .Q ( signal_1806 ) ) ;
    buf_clk cell_468 ( .C ( clk ), .D ( signal_1807 ), .Q ( signal_1808 ) ) ;
    buf_clk cell_470 ( .C ( clk ), .D ( signal_1809 ), .Q ( signal_1810 ) ) ;
    buf_clk cell_472 ( .C ( clk ), .D ( signal_1811 ), .Q ( signal_1812 ) ) ;
    buf_clk cell_474 ( .C ( clk ), .D ( signal_1813 ), .Q ( signal_1814 ) ) ;
    buf_clk cell_476 ( .C ( clk ), .D ( signal_1815 ), .Q ( signal_1816 ) ) ;
    buf_clk cell_480 ( .C ( clk ), .D ( signal_1819 ), .Q ( signal_1820 ) ) ;
    buf_clk cell_486 ( .C ( clk ), .D ( signal_1825 ), .Q ( signal_1826 ) ) ;
    buf_clk cell_492 ( .C ( clk ), .D ( signal_1831 ), .Q ( signal_1832 ) ) ;
    buf_clk cell_498 ( .C ( clk ), .D ( signal_1837 ), .Q ( signal_1838 ) ) ;
    buf_clk cell_504 ( .C ( clk ), .D ( signal_1843 ), .Q ( signal_1844 ) ) ;
    buf_clk cell_510 ( .C ( clk ), .D ( signal_1849 ), .Q ( signal_1850 ) ) ;
    buf_clk cell_516 ( .C ( clk ), .D ( signal_1855 ), .Q ( signal_1856 ) ) ;
    buf_clk cell_522 ( .C ( clk ), .D ( signal_1861 ), .Q ( signal_1862 ) ) ;
    buf_clk cell_528 ( .C ( clk ), .D ( signal_1867 ), .Q ( signal_1868 ) ) ;
    buf_clk cell_534 ( .C ( clk ), .D ( signal_1873 ), .Q ( signal_1874 ) ) ;
    buf_clk cell_540 ( .C ( clk ), .D ( signal_1879 ), .Q ( signal_1880 ) ) ;
    buf_clk cell_546 ( .C ( clk ), .D ( signal_1885 ), .Q ( signal_1886 ) ) ;
    buf_clk cell_552 ( .C ( clk ), .D ( signal_1891 ), .Q ( signal_1892 ) ) ;
    buf_clk cell_558 ( .C ( clk ), .D ( signal_1897 ), .Q ( signal_1898 ) ) ;
    buf_clk cell_564 ( .C ( clk ), .D ( signal_1903 ), .Q ( signal_1904 ) ) ;
    buf_clk cell_570 ( .C ( clk ), .D ( signal_1909 ), .Q ( signal_1910 ) ) ;
    buf_clk cell_576 ( .C ( clk ), .D ( signal_1915 ), .Q ( signal_1916 ) ) ;
    buf_clk cell_582 ( .C ( clk ), .D ( signal_1921 ), .Q ( signal_1922 ) ) ;
    buf_clk cell_588 ( .C ( clk ), .D ( signal_1927 ), .Q ( signal_1928 ) ) ;
    buf_clk cell_594 ( .C ( clk ), .D ( signal_1933 ), .Q ( signal_1934 ) ) ;
    buf_clk cell_600 ( .C ( clk ), .D ( signal_1939 ), .Q ( signal_1940 ) ) ;
    buf_clk cell_606 ( .C ( clk ), .D ( signal_1945 ), .Q ( signal_1946 ) ) ;
    buf_clk cell_612 ( .C ( clk ), .D ( signal_1951 ), .Q ( signal_1952 ) ) ;
    buf_clk cell_618 ( .C ( clk ), .D ( signal_1957 ), .Q ( signal_1958 ) ) ;
    buf_clk cell_624 ( .C ( clk ), .D ( signal_1963 ), .Q ( signal_1964 ) ) ;
    buf_clk cell_630 ( .C ( clk ), .D ( signal_1969 ), .Q ( signal_1970 ) ) ;
    buf_clk cell_636 ( .C ( clk ), .D ( signal_1975 ), .Q ( signal_1976 ) ) ;
    buf_clk cell_642 ( .C ( clk ), .D ( signal_1981 ), .Q ( signal_1982 ) ) ;
    buf_clk cell_648 ( .C ( clk ), .D ( signal_1987 ), .Q ( signal_1988 ) ) ;
    buf_clk cell_654 ( .C ( clk ), .D ( signal_1993 ), .Q ( signal_1994 ) ) ;
    buf_clk cell_660 ( .C ( clk ), .D ( signal_1999 ), .Q ( signal_2000 ) ) ;
    buf_clk cell_666 ( .C ( clk ), .D ( signal_2005 ), .Q ( signal_2006 ) ) ;
    buf_clk cell_672 ( .C ( clk ), .D ( signal_2011 ), .Q ( signal_2012 ) ) ;
    buf_clk cell_678 ( .C ( clk ), .D ( signal_2017 ), .Q ( signal_2018 ) ) ;
    buf_clk cell_684 ( .C ( clk ), .D ( signal_2023 ), .Q ( signal_2024 ) ) ;
    buf_clk cell_690 ( .C ( clk ), .D ( signal_2029 ), .Q ( signal_2030 ) ) ;
    buf_clk cell_696 ( .C ( clk ), .D ( signal_2035 ), .Q ( signal_2036 ) ) ;
    buf_clk cell_702 ( .C ( clk ), .D ( signal_2041 ), .Q ( signal_2042 ) ) ;
    buf_clk cell_708 ( .C ( clk ), .D ( signal_2047 ), .Q ( signal_2048 ) ) ;
    buf_clk cell_714 ( .C ( clk ), .D ( signal_2053 ), .Q ( signal_2054 ) ) ;
    buf_clk cell_720 ( .C ( clk ), .D ( signal_2059 ), .Q ( signal_2060 ) ) ;
    buf_clk cell_726 ( .C ( clk ), .D ( signal_2065 ), .Q ( signal_2066 ) ) ;
    buf_clk cell_732 ( .C ( clk ), .D ( signal_2071 ), .Q ( signal_2072 ) ) ;
    buf_clk cell_738 ( .C ( clk ), .D ( signal_2077 ), .Q ( signal_2078 ) ) ;
    buf_clk cell_744 ( .C ( clk ), .D ( signal_2083 ), .Q ( signal_2084 ) ) ;
    buf_clk cell_750 ( .C ( clk ), .D ( signal_2089 ), .Q ( signal_2090 ) ) ;
    buf_clk cell_756 ( .C ( clk ), .D ( signal_2095 ), .Q ( signal_2096 ) ) ;
    buf_clk cell_762 ( .C ( clk ), .D ( signal_2101 ), .Q ( signal_2102 ) ) ;
    buf_clk cell_768 ( .C ( clk ), .D ( signal_2107 ), .Q ( signal_2108 ) ) ;
    buf_clk cell_774 ( .C ( clk ), .D ( signal_2113 ), .Q ( signal_2114 ) ) ;
    buf_clk cell_780 ( .C ( clk ), .D ( signal_2119 ), .Q ( signal_2120 ) ) ;
    buf_clk cell_786 ( .C ( clk ), .D ( signal_2125 ), .Q ( signal_2126 ) ) ;
    buf_clk cell_792 ( .C ( clk ), .D ( signal_2131 ), .Q ( signal_2132 ) ) ;
    buf_clk cell_798 ( .C ( clk ), .D ( signal_2137 ), .Q ( signal_2138 ) ) ;
    buf_clk cell_804 ( .C ( clk ), .D ( signal_2143 ), .Q ( signal_2144 ) ) ;
    buf_clk cell_810 ( .C ( clk ), .D ( signal_2149 ), .Q ( signal_2150 ) ) ;
    buf_clk cell_816 ( .C ( clk ), .D ( signal_2155 ), .Q ( signal_2156 ) ) ;
    buf_clk cell_822 ( .C ( clk ), .D ( signal_2161 ), .Q ( signal_2162 ) ) ;
    buf_clk cell_828 ( .C ( clk ), .D ( signal_2167 ), .Q ( signal_2168 ) ) ;
    buf_clk cell_834 ( .C ( clk ), .D ( signal_2173 ), .Q ( signal_2174 ) ) ;
    buf_clk cell_840 ( .C ( clk ), .D ( signal_2179 ), .Q ( signal_2180 ) ) ;
    buf_clk cell_846 ( .C ( clk ), .D ( signal_2185 ), .Q ( signal_2186 ) ) ;
    buf_clk cell_852 ( .C ( clk ), .D ( signal_2191 ), .Q ( signal_2192 ) ) ;
    buf_clk cell_858 ( .C ( clk ), .D ( signal_2197 ), .Q ( signal_2198 ) ) ;
    buf_clk cell_864 ( .C ( clk ), .D ( signal_2203 ), .Q ( signal_2204 ) ) ;
    buf_clk cell_870 ( .C ( clk ), .D ( signal_2209 ), .Q ( signal_2210 ) ) ;
    buf_clk cell_876 ( .C ( clk ), .D ( signal_2215 ), .Q ( signal_2216 ) ) ;
    buf_clk cell_882 ( .C ( clk ), .D ( signal_2221 ), .Q ( signal_2222 ) ) ;
    buf_clk cell_888 ( .C ( clk ), .D ( signal_2227 ), .Q ( signal_2228 ) ) ;
    buf_clk cell_894 ( .C ( clk ), .D ( signal_2233 ), .Q ( signal_2234 ) ) ;
    buf_clk cell_900 ( .C ( clk ), .D ( signal_2239 ), .Q ( signal_2240 ) ) ;
    buf_clk cell_906 ( .C ( clk ), .D ( signal_2245 ), .Q ( signal_2246 ) ) ;
    buf_clk cell_916 ( .C ( clk ), .D ( signal_2255 ), .Q ( signal_2256 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_481 ( .C ( clk ), .D ( signal_1820 ), .Q ( signal_1821 ) ) ;
    buf_clk cell_487 ( .C ( clk ), .D ( signal_1826 ), .Q ( signal_1827 ) ) ;
    buf_clk cell_493 ( .C ( clk ), .D ( signal_1832 ), .Q ( signal_1833 ) ) ;
    buf_clk cell_499 ( .C ( clk ), .D ( signal_1838 ), .Q ( signal_1839 ) ) ;
    buf_clk cell_505 ( .C ( clk ), .D ( signal_1844 ), .Q ( signal_1845 ) ) ;
    buf_clk cell_511 ( .C ( clk ), .D ( signal_1850 ), .Q ( signal_1851 ) ) ;
    buf_clk cell_517 ( .C ( clk ), .D ( signal_1856 ), .Q ( signal_1857 ) ) ;
    buf_clk cell_523 ( .C ( clk ), .D ( signal_1862 ), .Q ( signal_1863 ) ) ;
    buf_clk cell_529 ( .C ( clk ), .D ( signal_1868 ), .Q ( signal_1869 ) ) ;
    buf_clk cell_535 ( .C ( clk ), .D ( signal_1874 ), .Q ( signal_1875 ) ) ;
    buf_clk cell_541 ( .C ( clk ), .D ( signal_1880 ), .Q ( signal_1881 ) ) ;
    buf_clk cell_547 ( .C ( clk ), .D ( signal_1886 ), .Q ( signal_1887 ) ) ;
    buf_clk cell_553 ( .C ( clk ), .D ( signal_1892 ), .Q ( signal_1893 ) ) ;
    buf_clk cell_559 ( .C ( clk ), .D ( signal_1898 ), .Q ( signal_1899 ) ) ;
    buf_clk cell_565 ( .C ( clk ), .D ( signal_1904 ), .Q ( signal_1905 ) ) ;
    buf_clk cell_571 ( .C ( clk ), .D ( signal_1910 ), .Q ( signal_1911 ) ) ;
    buf_clk cell_577 ( .C ( clk ), .D ( signal_1916 ), .Q ( signal_1917 ) ) ;
    buf_clk cell_583 ( .C ( clk ), .D ( signal_1922 ), .Q ( signal_1923 ) ) ;
    buf_clk cell_589 ( .C ( clk ), .D ( signal_1928 ), .Q ( signal_1929 ) ) ;
    buf_clk cell_595 ( .C ( clk ), .D ( signal_1934 ), .Q ( signal_1935 ) ) ;
    buf_clk cell_601 ( .C ( clk ), .D ( signal_1940 ), .Q ( signal_1941 ) ) ;
    buf_clk cell_607 ( .C ( clk ), .D ( signal_1946 ), .Q ( signal_1947 ) ) ;
    buf_clk cell_613 ( .C ( clk ), .D ( signal_1952 ), .Q ( signal_1953 ) ) ;
    buf_clk cell_619 ( .C ( clk ), .D ( signal_1958 ), .Q ( signal_1959 ) ) ;
    buf_clk cell_625 ( .C ( clk ), .D ( signal_1964 ), .Q ( signal_1965 ) ) ;
    buf_clk cell_631 ( .C ( clk ), .D ( signal_1970 ), .Q ( signal_1971 ) ) ;
    buf_clk cell_637 ( .C ( clk ), .D ( signal_1976 ), .Q ( signal_1977 ) ) ;
    buf_clk cell_643 ( .C ( clk ), .D ( signal_1982 ), .Q ( signal_1983 ) ) ;
    buf_clk cell_649 ( .C ( clk ), .D ( signal_1988 ), .Q ( signal_1989 ) ) ;
    buf_clk cell_655 ( .C ( clk ), .D ( signal_1994 ), .Q ( signal_1995 ) ) ;
    buf_clk cell_661 ( .C ( clk ), .D ( signal_2000 ), .Q ( signal_2001 ) ) ;
    buf_clk cell_667 ( .C ( clk ), .D ( signal_2006 ), .Q ( signal_2007 ) ) ;
    buf_clk cell_673 ( .C ( clk ), .D ( signal_2012 ), .Q ( signal_2013 ) ) ;
    buf_clk cell_679 ( .C ( clk ), .D ( signal_2018 ), .Q ( signal_2019 ) ) ;
    buf_clk cell_685 ( .C ( clk ), .D ( signal_2024 ), .Q ( signal_2025 ) ) ;
    buf_clk cell_691 ( .C ( clk ), .D ( signal_2030 ), .Q ( signal_2031 ) ) ;
    buf_clk cell_697 ( .C ( clk ), .D ( signal_2036 ), .Q ( signal_2037 ) ) ;
    buf_clk cell_703 ( .C ( clk ), .D ( signal_2042 ), .Q ( signal_2043 ) ) ;
    buf_clk cell_709 ( .C ( clk ), .D ( signal_2048 ), .Q ( signal_2049 ) ) ;
    buf_clk cell_715 ( .C ( clk ), .D ( signal_2054 ), .Q ( signal_2055 ) ) ;
    buf_clk cell_721 ( .C ( clk ), .D ( signal_2060 ), .Q ( signal_2061 ) ) ;
    buf_clk cell_727 ( .C ( clk ), .D ( signal_2066 ), .Q ( signal_2067 ) ) ;
    buf_clk cell_733 ( .C ( clk ), .D ( signal_2072 ), .Q ( signal_2073 ) ) ;
    buf_clk cell_739 ( .C ( clk ), .D ( signal_2078 ), .Q ( signal_2079 ) ) ;
    buf_clk cell_745 ( .C ( clk ), .D ( signal_2084 ), .Q ( signal_2085 ) ) ;
    buf_clk cell_751 ( .C ( clk ), .D ( signal_2090 ), .Q ( signal_2091 ) ) ;
    buf_clk cell_757 ( .C ( clk ), .D ( signal_2096 ), .Q ( signal_2097 ) ) ;
    buf_clk cell_763 ( .C ( clk ), .D ( signal_2102 ), .Q ( signal_2103 ) ) ;
    buf_clk cell_769 ( .C ( clk ), .D ( signal_2108 ), .Q ( signal_2109 ) ) ;
    buf_clk cell_775 ( .C ( clk ), .D ( signal_2114 ), .Q ( signal_2115 ) ) ;
    buf_clk cell_781 ( .C ( clk ), .D ( signal_2120 ), .Q ( signal_2121 ) ) ;
    buf_clk cell_787 ( .C ( clk ), .D ( signal_2126 ), .Q ( signal_2127 ) ) ;
    buf_clk cell_793 ( .C ( clk ), .D ( signal_2132 ), .Q ( signal_2133 ) ) ;
    buf_clk cell_799 ( .C ( clk ), .D ( signal_2138 ), .Q ( signal_2139 ) ) ;
    buf_clk cell_805 ( .C ( clk ), .D ( signal_2144 ), .Q ( signal_2145 ) ) ;
    buf_clk cell_811 ( .C ( clk ), .D ( signal_2150 ), .Q ( signal_2151 ) ) ;
    buf_clk cell_817 ( .C ( clk ), .D ( signal_2156 ), .Q ( signal_2157 ) ) ;
    buf_clk cell_823 ( .C ( clk ), .D ( signal_2162 ), .Q ( signal_2163 ) ) ;
    buf_clk cell_829 ( .C ( clk ), .D ( signal_2168 ), .Q ( signal_2169 ) ) ;
    buf_clk cell_835 ( .C ( clk ), .D ( signal_2174 ), .Q ( signal_2175 ) ) ;
    buf_clk cell_841 ( .C ( clk ), .D ( signal_2180 ), .Q ( signal_2181 ) ) ;
    buf_clk cell_847 ( .C ( clk ), .D ( signal_2186 ), .Q ( signal_2187 ) ) ;
    buf_clk cell_853 ( .C ( clk ), .D ( signal_2192 ), .Q ( signal_2193 ) ) ;
    buf_clk cell_859 ( .C ( clk ), .D ( signal_2198 ), .Q ( signal_2199 ) ) ;
    buf_clk cell_865 ( .C ( clk ), .D ( signal_2204 ), .Q ( signal_2205 ) ) ;
    buf_clk cell_871 ( .C ( clk ), .D ( signal_2210 ), .Q ( signal_2211 ) ) ;
    buf_clk cell_877 ( .C ( clk ), .D ( signal_2216 ), .Q ( signal_2217 ) ) ;
    buf_clk cell_883 ( .C ( clk ), .D ( signal_2222 ), .Q ( signal_2223 ) ) ;
    buf_clk cell_889 ( .C ( clk ), .D ( signal_2228 ), .Q ( signal_2229 ) ) ;
    buf_clk cell_895 ( .C ( clk ), .D ( signal_2234 ), .Q ( signal_2235 ) ) ;
    buf_clk cell_901 ( .C ( clk ), .D ( signal_2240 ), .Q ( signal_2241 ) ) ;
    buf_clk cell_907 ( .C ( clk ), .D ( signal_2246 ), .Q ( signal_2247 ) ) ;
    buf_clk cell_917 ( .C ( clk ), .D ( signal_2256 ), .Q ( signal_2257 ) ) ;

    /* cells in depth 10 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_305 ( .a ({signal_1776, signal_1774, signal_1772, signal_1770}), .b ({signal_838, signal_837, signal_836, signal_318}), .clk ( clk ), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_847, signal_846, signal_845, signal_321}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_306 ( .a ({signal_1784, signal_1782, signal_1780, signal_1778}), .b ({signal_838, signal_837, signal_836, signal_318}), .clk ( clk ), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({signal_850, signal_849, signal_848, signal_322}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_308 ( .a ({signal_1792, signal_1790, signal_1788, signal_1786}), .b ({signal_844, signal_843, signal_842, signal_320}), .clk ( clk ), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({signal_856, signal_855, signal_854, signal_324}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_309 ( .a ({signal_1800, signal_1798, signal_1796, signal_1794}), .b ({signal_844, signal_843, signal_842, signal_320}), .clk ( clk ), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({signal_859, signal_858, signal_857, signal_325}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_310 ( .a ({signal_1808, signal_1806, signal_1804, signal_1802}), .b ({signal_853, signal_852, signal_851, signal_323}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({signal_862, signal_861, signal_860, signal_326}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_311 ( .a ({signal_1816, signal_1814, signal_1812, signal_1810}), .b ({signal_853, signal_852, signal_851, signal_323}), .clk ( clk ), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_865, signal_864, signal_863, signal_327}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_312 ( .a ({signal_856, signal_855, signal_854, signal_324}), .b ({signal_862, signal_861, signal_860, signal_326}), .c ({signal_868, signal_867, signal_866, signal_328}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_313 ( .a ({signal_847, signal_846, signal_845, signal_321}), .b ({signal_862, signal_861, signal_860, signal_326}), .c ({signal_871, signal_870, signal_869, signal_329}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_314 ( .a ({signal_859, signal_858, signal_857, signal_325}), .b ({signal_865, signal_864, signal_863, signal_327}), .c ({signal_874, signal_873, signal_872, signal_330}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_315 ( .a ({signal_850, signal_849, signal_848, signal_322}), .b ({signal_865, signal_864, signal_863, signal_327}), .c ({signal_877, signal_876, signal_875, signal_331}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_324 ( .a ({signal_874, signal_873, signal_872, signal_330}), .b ({signal_877, signal_876, signal_875, signal_331}), .c ({signal_904, signal_903, signal_902, signal_340}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_325 ( .a ({signal_868, signal_867, signal_866, signal_328}), .b ({signal_871, signal_870, signal_869, signal_329}), .c ({signal_907, signal_906, signal_905, signal_341}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_326 ( .a ({signal_871, signal_870, signal_869, signal_329}), .b ({signal_877, signal_876, signal_875, signal_331}), .c ({signal_910, signal_909, signal_908, signal_342}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_327 ( .a ({signal_868, signal_867, signal_866, signal_328}), .b ({signal_874, signal_873, signal_872, signal_330}), .c ({signal_913, signal_912, signal_911, signal_343}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_336 ( .a ({signal_910, signal_909, signal_908, signal_342}), .b ({signal_913, signal_912, signal_911, signal_343}), .c ({signal_940, signal_939, signal_938, signal_352}) ) ;
    buf_clk cell_482 ( .C ( clk ), .D ( signal_1821 ), .Q ( signal_1822 ) ) ;
    buf_clk cell_488 ( .C ( clk ), .D ( signal_1827 ), .Q ( signal_1828 ) ) ;
    buf_clk cell_494 ( .C ( clk ), .D ( signal_1833 ), .Q ( signal_1834 ) ) ;
    buf_clk cell_500 ( .C ( clk ), .D ( signal_1839 ), .Q ( signal_1840 ) ) ;
    buf_clk cell_506 ( .C ( clk ), .D ( signal_1845 ), .Q ( signal_1846 ) ) ;
    buf_clk cell_512 ( .C ( clk ), .D ( signal_1851 ), .Q ( signal_1852 ) ) ;
    buf_clk cell_518 ( .C ( clk ), .D ( signal_1857 ), .Q ( signal_1858 ) ) ;
    buf_clk cell_524 ( .C ( clk ), .D ( signal_1863 ), .Q ( signal_1864 ) ) ;
    buf_clk cell_530 ( .C ( clk ), .D ( signal_1869 ), .Q ( signal_1870 ) ) ;
    buf_clk cell_536 ( .C ( clk ), .D ( signal_1875 ), .Q ( signal_1876 ) ) ;
    buf_clk cell_542 ( .C ( clk ), .D ( signal_1881 ), .Q ( signal_1882 ) ) ;
    buf_clk cell_548 ( .C ( clk ), .D ( signal_1887 ), .Q ( signal_1888 ) ) ;
    buf_clk cell_554 ( .C ( clk ), .D ( signal_1893 ), .Q ( signal_1894 ) ) ;
    buf_clk cell_560 ( .C ( clk ), .D ( signal_1899 ), .Q ( signal_1900 ) ) ;
    buf_clk cell_566 ( .C ( clk ), .D ( signal_1905 ), .Q ( signal_1906 ) ) ;
    buf_clk cell_572 ( .C ( clk ), .D ( signal_1911 ), .Q ( signal_1912 ) ) ;
    buf_clk cell_578 ( .C ( clk ), .D ( signal_1917 ), .Q ( signal_1918 ) ) ;
    buf_clk cell_584 ( .C ( clk ), .D ( signal_1923 ), .Q ( signal_1924 ) ) ;
    buf_clk cell_590 ( .C ( clk ), .D ( signal_1929 ), .Q ( signal_1930 ) ) ;
    buf_clk cell_596 ( .C ( clk ), .D ( signal_1935 ), .Q ( signal_1936 ) ) ;
    buf_clk cell_602 ( .C ( clk ), .D ( signal_1941 ), .Q ( signal_1942 ) ) ;
    buf_clk cell_608 ( .C ( clk ), .D ( signal_1947 ), .Q ( signal_1948 ) ) ;
    buf_clk cell_614 ( .C ( clk ), .D ( signal_1953 ), .Q ( signal_1954 ) ) ;
    buf_clk cell_620 ( .C ( clk ), .D ( signal_1959 ), .Q ( signal_1960 ) ) ;
    buf_clk cell_626 ( .C ( clk ), .D ( signal_1965 ), .Q ( signal_1966 ) ) ;
    buf_clk cell_632 ( .C ( clk ), .D ( signal_1971 ), .Q ( signal_1972 ) ) ;
    buf_clk cell_638 ( .C ( clk ), .D ( signal_1977 ), .Q ( signal_1978 ) ) ;
    buf_clk cell_644 ( .C ( clk ), .D ( signal_1983 ), .Q ( signal_1984 ) ) ;
    buf_clk cell_650 ( .C ( clk ), .D ( signal_1989 ), .Q ( signal_1990 ) ) ;
    buf_clk cell_656 ( .C ( clk ), .D ( signal_1995 ), .Q ( signal_1996 ) ) ;
    buf_clk cell_662 ( .C ( clk ), .D ( signal_2001 ), .Q ( signal_2002 ) ) ;
    buf_clk cell_668 ( .C ( clk ), .D ( signal_2007 ), .Q ( signal_2008 ) ) ;
    buf_clk cell_674 ( .C ( clk ), .D ( signal_2013 ), .Q ( signal_2014 ) ) ;
    buf_clk cell_680 ( .C ( clk ), .D ( signal_2019 ), .Q ( signal_2020 ) ) ;
    buf_clk cell_686 ( .C ( clk ), .D ( signal_2025 ), .Q ( signal_2026 ) ) ;
    buf_clk cell_692 ( .C ( clk ), .D ( signal_2031 ), .Q ( signal_2032 ) ) ;
    buf_clk cell_698 ( .C ( clk ), .D ( signal_2037 ), .Q ( signal_2038 ) ) ;
    buf_clk cell_704 ( .C ( clk ), .D ( signal_2043 ), .Q ( signal_2044 ) ) ;
    buf_clk cell_710 ( .C ( clk ), .D ( signal_2049 ), .Q ( signal_2050 ) ) ;
    buf_clk cell_716 ( .C ( clk ), .D ( signal_2055 ), .Q ( signal_2056 ) ) ;
    buf_clk cell_722 ( .C ( clk ), .D ( signal_2061 ), .Q ( signal_2062 ) ) ;
    buf_clk cell_728 ( .C ( clk ), .D ( signal_2067 ), .Q ( signal_2068 ) ) ;
    buf_clk cell_734 ( .C ( clk ), .D ( signal_2073 ), .Q ( signal_2074 ) ) ;
    buf_clk cell_740 ( .C ( clk ), .D ( signal_2079 ), .Q ( signal_2080 ) ) ;
    buf_clk cell_746 ( .C ( clk ), .D ( signal_2085 ), .Q ( signal_2086 ) ) ;
    buf_clk cell_752 ( .C ( clk ), .D ( signal_2091 ), .Q ( signal_2092 ) ) ;
    buf_clk cell_758 ( .C ( clk ), .D ( signal_2097 ), .Q ( signal_2098 ) ) ;
    buf_clk cell_764 ( .C ( clk ), .D ( signal_2103 ), .Q ( signal_2104 ) ) ;
    buf_clk cell_770 ( .C ( clk ), .D ( signal_2109 ), .Q ( signal_2110 ) ) ;
    buf_clk cell_776 ( .C ( clk ), .D ( signal_2115 ), .Q ( signal_2116 ) ) ;
    buf_clk cell_782 ( .C ( clk ), .D ( signal_2121 ), .Q ( signal_2122 ) ) ;
    buf_clk cell_788 ( .C ( clk ), .D ( signal_2127 ), .Q ( signal_2128 ) ) ;
    buf_clk cell_794 ( .C ( clk ), .D ( signal_2133 ), .Q ( signal_2134 ) ) ;
    buf_clk cell_800 ( .C ( clk ), .D ( signal_2139 ), .Q ( signal_2140 ) ) ;
    buf_clk cell_806 ( .C ( clk ), .D ( signal_2145 ), .Q ( signal_2146 ) ) ;
    buf_clk cell_812 ( .C ( clk ), .D ( signal_2151 ), .Q ( signal_2152 ) ) ;
    buf_clk cell_818 ( .C ( clk ), .D ( signal_2157 ), .Q ( signal_2158 ) ) ;
    buf_clk cell_824 ( .C ( clk ), .D ( signal_2163 ), .Q ( signal_2164 ) ) ;
    buf_clk cell_830 ( .C ( clk ), .D ( signal_2169 ), .Q ( signal_2170 ) ) ;
    buf_clk cell_836 ( .C ( clk ), .D ( signal_2175 ), .Q ( signal_2176 ) ) ;
    buf_clk cell_842 ( .C ( clk ), .D ( signal_2181 ), .Q ( signal_2182 ) ) ;
    buf_clk cell_848 ( .C ( clk ), .D ( signal_2187 ), .Q ( signal_2188 ) ) ;
    buf_clk cell_854 ( .C ( clk ), .D ( signal_2193 ), .Q ( signal_2194 ) ) ;
    buf_clk cell_860 ( .C ( clk ), .D ( signal_2199 ), .Q ( signal_2200 ) ) ;
    buf_clk cell_866 ( .C ( clk ), .D ( signal_2205 ), .Q ( signal_2206 ) ) ;
    buf_clk cell_872 ( .C ( clk ), .D ( signal_2211 ), .Q ( signal_2212 ) ) ;
    buf_clk cell_878 ( .C ( clk ), .D ( signal_2217 ), .Q ( signal_2218 ) ) ;
    buf_clk cell_884 ( .C ( clk ), .D ( signal_2223 ), .Q ( signal_2224 ) ) ;
    buf_clk cell_890 ( .C ( clk ), .D ( signal_2229 ), .Q ( signal_2230 ) ) ;
    buf_clk cell_896 ( .C ( clk ), .D ( signal_2235 ), .Q ( signal_2236 ) ) ;
    buf_clk cell_902 ( .C ( clk ), .D ( signal_2241 ), .Q ( signal_2242 ) ) ;
    buf_clk cell_908 ( .C ( clk ), .D ( signal_2247 ), .Q ( signal_2248 ) ) ;
    buf_clk cell_918 ( .C ( clk ), .D ( signal_2257 ), .Q ( signal_2258 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_919 ( .C ( clk ), .D ( signal_2258 ), .Q ( signal_2259 ) ) ;

    /* cells in depth 12 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_316 ( .a ({signal_1840, signal_1834, signal_1828, signal_1822}), .b ({signal_868, signal_867, signal_866, signal_328}), .clk ( clk ), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({signal_880, signal_879, signal_878, signal_332}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_317 ( .a ({signal_1864, signal_1858, signal_1852, signal_1846}), .b ({signal_871, signal_870, signal_869, signal_329}), .clk ( clk ), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({signal_883, signal_882, signal_881, signal_333}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_318 ( .a ({signal_1888, signal_1882, signal_1876, signal_1870}), .b ({signal_874, signal_873, signal_872, signal_330}), .clk ( clk ), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({signal_886, signal_885, signal_884, signal_334}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_319 ( .a ({signal_1912, signal_1906, signal_1900, signal_1894}), .b ({signal_877, signal_876, signal_875, signal_331}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({signal_889, signal_888, signal_887, signal_335}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_320 ( .a ({signal_1936, signal_1930, signal_1924, signal_1918}), .b ({signal_868, signal_867, signal_866, signal_328}), .clk ( clk ), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_892, signal_891, signal_890, signal_336}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_321 ( .a ({signal_1960, signal_1954, signal_1948, signal_1942}), .b ({signal_871, signal_870, signal_869, signal_329}), .clk ( clk ), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({signal_895, signal_894, signal_893, signal_337}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_322 ( .a ({signal_1984, signal_1978, signal_1972, signal_1966}), .b ({signal_874, signal_873, signal_872, signal_330}), .clk ( clk ), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({signal_898, signal_897, signal_896, signal_338}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_323 ( .a ({signal_2008, signal_2002, signal_1996, signal_1990}), .b ({signal_877, signal_876, signal_875, signal_331}), .clk ( clk ), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({signal_901, signal_900, signal_899, signal_339}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_328 ( .a ({signal_2032, signal_2026, signal_2020, signal_2014}), .b ({signal_907, signal_906, signal_905, signal_341}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({signal_916, signal_915, signal_914, signal_344}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_329 ( .a ({signal_2056, signal_2050, signal_2044, signal_2038}), .b ({signal_904, signal_903, signal_902, signal_340}), .clk ( clk ), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_919, signal_918, signal_917, signal_345}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_330 ( .a ({signal_2080, signal_2074, signal_2068, signal_2062}), .b ({signal_913, signal_912, signal_911, signal_343}), .clk ( clk ), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({signal_922, signal_921, signal_920, signal_346}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_331 ( .a ({signal_2104, signal_2098, signal_2092, signal_2086}), .b ({signal_910, signal_909, signal_908, signal_342}), .clk ( clk ), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({signal_925, signal_924, signal_923, signal_347}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_332 ( .a ({signal_2128, signal_2122, signal_2116, signal_2110}), .b ({signal_907, signal_906, signal_905, signal_341}), .clk ( clk ), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({signal_928, signal_927, signal_926, signal_348}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_333 ( .a ({signal_2152, signal_2146, signal_2140, signal_2134}), .b ({signal_904, signal_903, signal_902, signal_340}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({signal_931, signal_930, signal_929, signal_349}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_334 ( .a ({signal_2176, signal_2170, signal_2164, signal_2158}), .b ({signal_913, signal_912, signal_911, signal_343}), .clk ( clk ), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_934, signal_933, signal_932, signal_350}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_335 ( .a ({signal_2200, signal_2194, signal_2188, signal_2182}), .b ({signal_910, signal_909, signal_908, signal_342}), .clk ( clk ), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({signal_937, signal_936, signal_935, signal_351}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_337 ( .a ({signal_2224, signal_2218, signal_2212, signal_2206}), .b ({signal_940, signal_939, signal_938, signal_352}), .clk ( clk ), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({signal_943, signal_942, signal_941, signal_353}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_338 ( .a ({signal_2248, signal_2242, signal_2236, signal_2230}), .b ({signal_940, signal_939, signal_938, signal_352}), .clk ( clk ), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({signal_946, signal_945, signal_944, signal_354}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_339 ( .a ({signal_880, signal_879, signal_878, signal_332}), .b ({signal_916, signal_915, signal_914, signal_344}), .c ({signal_949, signal_948, signal_947, signal_355}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_340 ( .a ({signal_883, signal_882, signal_881, signal_333}), .b ({signal_916, signal_915, signal_914, signal_344}), .c ({signal_952, signal_951, signal_950, signal_356}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_341 ( .a ({signal_886, signal_885, signal_884, signal_334}), .b ({signal_919, signal_918, signal_917, signal_345}), .c ({signal_955, signal_954, signal_953, signal_357}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_342 ( .a ({signal_889, signal_888, signal_887, signal_335}), .b ({signal_919, signal_918, signal_917, signal_345}), .c ({signal_958, signal_957, signal_956, signal_358}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_343 ( .a ({signal_922, signal_921, signal_920, signal_346}), .b ({signal_925, signal_924, signal_923, signal_347}), .c ({signal_961, signal_960, signal_959, signal_359}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_344 ( .a ({signal_892, signal_891, signal_890, signal_336}), .b ({signal_928, signal_927, signal_926, signal_348}), .c ({signal_964, signal_963, signal_962, signal_360}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_345 ( .a ({signal_895, signal_894, signal_893, signal_337}), .b ({signal_928, signal_927, signal_926, signal_348}), .c ({signal_967, signal_966, signal_965, signal_361}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_346 ( .a ({signal_898, signal_897, signal_896, signal_338}), .b ({signal_931, signal_930, signal_929, signal_349}), .c ({signal_970, signal_969, signal_968, signal_362}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_347 ( .a ({signal_901, signal_900, signal_899, signal_339}), .b ({signal_931, signal_930, signal_929, signal_349}), .c ({signal_973, signal_972, signal_971, signal_363}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_348 ( .a ({signal_934, signal_933, signal_932, signal_350}), .b ({signal_937, signal_936, signal_935, signal_351}), .c ({signal_976, signal_975, signal_974, signal_364}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_349 ( .a ({signal_952, signal_951, signal_950, signal_356}), .b ({signal_961, signal_960, signal_959, signal_359}), .c ({signal_979, signal_978, signal_977, signal_365}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_350 ( .a ({signal_958, signal_957, signal_956, signal_358}), .b ({signal_961, signal_960, signal_959, signal_359}), .c ({signal_982, signal_981, signal_980, signal_366}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_351 ( .a ({signal_925, signal_924, signal_923, signal_347}), .b ({signal_943, signal_942, signal_941, signal_353}), .c ({signal_985, signal_984, signal_983, signal_367}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_352 ( .a ({signal_967, signal_966, signal_965, signal_361}), .b ({signal_976, signal_975, signal_974, signal_364}), .c ({signal_988, signal_987, signal_986, signal_368}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_353 ( .a ({signal_973, signal_972, signal_971, signal_363}), .b ({signal_976, signal_975, signal_974, signal_364}), .c ({signal_991, signal_990, signal_989, signal_369}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_354 ( .a ({signal_937, signal_936, signal_935, signal_351}), .b ({signal_946, signal_945, signal_944, signal_354}), .c ({signal_994, signal_993, signal_992, signal_370}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_355 ( .a ({signal_988, signal_987, signal_986, signal_368}), .b ({signal_997, signal_996, signal_995, signal_371}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_356 ( .a ({signal_979, signal_978, signal_977, signal_365}), .b ({signal_991, signal_990, signal_989, signal_369}), .c ({signal_1000, signal_999, signal_998, signal_372}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_357 ( .a ({signal_979, signal_978, signal_977, signal_365}), .b ({signal_982, signal_981, signal_980, signal_366}), .c ({signal_1003, signal_1002, signal_1001, signal_373}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_358 ( .a ({signal_949, signal_948, signal_947, signal_355}), .b ({signal_985, signal_984, signal_983, signal_367}), .c ({signal_1006, signal_1005, signal_1004, signal_374}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_359 ( .a ({signal_955, signal_954, signal_953, signal_357}), .b ({signal_985, signal_984, signal_983, signal_367}), .c ({signal_1009, signal_1008, signal_1007, signal_375}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_360 ( .a ({signal_964, signal_963, signal_962, signal_360}), .b ({signal_994, signal_993, signal_992, signal_370}), .c ({signal_1012, signal_1011, signal_1010, signal_376}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_361 ( .a ({signal_970, signal_969, signal_968, signal_362}), .b ({signal_994, signal_993, signal_992, signal_370}), .c ({signal_1015, signal_1014, signal_1013, signal_377}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_364 ( .a ({signal_1009, signal_1008, signal_1007, signal_375}), .b ({signal_1015, signal_1014, signal_1013, signal_377}), .c ({signal_1024, signal_1023, signal_1022, signal_380}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_365 ( .a ({signal_982, signal_981, signal_980, signal_366}), .b ({signal_1015, signal_1014, signal_1013, signal_377}), .c ({signal_1027, signal_1026, signal_1025, signal_381}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_366 ( .a ({signal_979, signal_978, signal_977, signal_365}), .b ({signal_1015, signal_1014, signal_1013, signal_377}), .c ({signal_1030, signal_1029, signal_1028, signal_382}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_367 ( .a ({signal_1006, signal_1005, signal_1004, signal_374}), .b ({signal_1012, signal_1011, signal_1010, signal_376}), .c ({signal_1033, signal_1032, signal_1031, signal_383}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_368 ( .a ({signal_1009, signal_1008, signal_1007, signal_375}), .b ({signal_1012, signal_1011, signal_1010, signal_376}), .c ({signal_1036, signal_1035, signal_1034, signal_384}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_369 ( .a ({signal_1003, signal_1002, signal_1001, signal_373}), .b ({signal_1015, signal_1014, signal_1013, signal_377}), .c ({signal_1039, signal_1038, signal_1037, signal_385}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_370 ( .a ({signal_1024, signal_1023, signal_1022, signal_380}), .b ({signal_1042, signal_1041, signal_1040, signal_386}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_371 ( .a ({signal_1027, signal_1026, signal_1025, signal_381}), .b ({signal_1045, signal_1044, signal_1043, signal_387}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_372 ( .a ({signal_1030, signal_1029, signal_1028, signal_382}), .b ({signal_1048, signal_1047, signal_1046, signal_388}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_373 ( .a ({signal_1036, signal_1035, signal_1034, signal_384}), .b ({signal_1051, signal_1050, signal_1049, signal_389}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_378 ( .a ({signal_982, signal_981, signal_980, signal_366}), .b ({signal_1024, signal_1023, signal_1022, signal_380}), .c ({signal_1066, signal_1065, signal_1064, signal_394}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_379 ( .a ({signal_1009, signal_1008, signal_1007, signal_375}), .b ({signal_1033, signal_1032, signal_1031, signal_383}), .c ({signal_1069, signal_1068, signal_1067, signal_395}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_380 ( .a ({signal_988, signal_987, signal_986, signal_368}), .b ({signal_1036, signal_1035, signal_1034, signal_384}), .c ({signal_1072, signal_1071, signal_1070, signal_396}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_381 ( .a ({signal_1069, signal_1068, signal_1067, signal_395}), .b ({signal_1075, signal_1074, signal_1073, signal_397}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_389 ( .a ({signal_1006, signal_1005, signal_1004, signal_374}), .b ({signal_1066, signal_1065, signal_1064, signal_394}), .c ({signal_1099, signal_1098, signal_1097, signal_405}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_390 ( .a ({signal_1000, signal_999, signal_998, signal_372}), .b ({signal_1069, signal_1068, signal_1067, signal_395}), .c ({signal_1102, signal_1101, signal_1100, signal_406}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_391 ( .a ({signal_1039, signal_1038, signal_1037, signal_385}), .b ({signal_1072, signal_1071, signal_1070, signal_396}), .c ({signal_1105, signal_1104, signal_1103, signal_407}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_392 ( .a ({signal_1003, signal_1002, signal_1001, signal_373}), .b ({signal_1069, signal_1068, signal_1067, signal_395}), .c ({signal_1108, signal_1107, signal_1106, signal_408}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_393 ( .a ({signal_1000, signal_999, signal_998, signal_372}), .b ({signal_1072, signal_1071, signal_1070, signal_396}), .c ({signal_1111, signal_1110, signal_1109, signal_409}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_396 ( .a ({signal_1099, signal_1098, signal_1097, signal_405}), .b ({signal_1120, signal_1119, signal_1118, signal_412}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_397 ( .a ({signal_1105, signal_1104, signal_1103, signal_407}), .b ({signal_1123, signal_1122, signal_1121, signal_413}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_398 ( .a ({signal_1108, signal_1107, signal_1106, signal_408}), .b ({signal_1126, signal_1125, signal_1124, signal_414}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_399 ( .a ({signal_1111, signal_1110, signal_1109, signal_409}), .b ({signal_1129, signal_1128, signal_1127, signal_415}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_405 ( .a ({signal_1015, signal_1014, signal_1013, signal_377}), .b ({signal_1102, signal_1101, signal_1100, signal_406}), .c ({signal_1147, signal_1146, signal_1145, signal_420}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_406 ( .a ({signal_988, signal_987, signal_986, signal_368}), .b ({signal_1102, signal_1101, signal_1100, signal_406}), .c ({signal_1150, signal_1149, signal_1148, signal_421}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_408 ( .a ({signal_1147, signal_1146, signal_1145, signal_420}), .b ({signal_1156, signal_1155, signal_1154, signal_423}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_409 ( .a ({signal_1150, signal_1149, signal_1148, signal_421}), .b ({signal_1159, signal_1158, signal_1157, signal_424}) ) ;
    buf_clk cell_920 ( .C ( clk ), .D ( signal_2259 ), .Q ( signal_2260 ) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_362 ( .a ({1'b0, 1'b0, 1'b0, signal_2260}), .b ({signal_997, signal_996, signal_995, signal_371}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({signal_1018, signal_1017, signal_1016, signal_378}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_363 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1000, signal_999, signal_998, signal_372}), .clk ( clk ), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_1021, signal_1020, signal_1019, signal_379}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_374 ( .a ({signal_1018, signal_1017, signal_1016, signal_378}), .b ({signal_1054, signal_1053, signal_1052, signal_390}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_375 ( .a ({signal_1021, signal_1020, signal_1019, signal_379}), .b ({signal_1057, signal_1056, signal_1055, signal_391}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_376 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1039, signal_1038, signal_1037, signal_385}), .clk ( clk ), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({signal_1060, signal_1059, signal_1058, signal_392}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_377 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1033, signal_1032, signal_1031, signal_383}), .clk ( clk ), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({signal_1063, signal_1062, signal_1061, signal_393}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_382 ( .a ({signal_1060, signal_1059, signal_1058, signal_392}), .b ({signal_1078, signal_1077, signal_1076, signal_398}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_383 ( .a ({signal_1063, signal_1062, signal_1061, signal_393}), .b ({signal_1081, signal_1080, signal_1079, signal_399}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_384 ( .a ({1'b0, 1'b0, 1'b0, signal_2260}), .b ({signal_1045, signal_1044, signal_1043, signal_387}), .clk ( clk ), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({signal_1084, signal_1083, signal_1082, signal_400}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_385 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1051, signal_1050, signal_1049, signal_389}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({signal_1087, signal_1086, signal_1085, signal_401}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_386 ( .a ({1'b0, 1'b0, 1'b0, signal_2260}), .b ({signal_1048, signal_1047, signal_1046, signal_388}), .clk ( clk ), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_1090, signal_1089, signal_1088, signal_402}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_387 ( .a ({1'b0, 1'b0, 1'b0, signal_2260}), .b ({signal_1042, signal_1041, signal_1040, signal_386}), .clk ( clk ), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({signal_1093, signal_1092, signal_1091, signal_403}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_388 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1066, signal_1065, signal_1064, signal_394}), .clk ( clk ), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({signal_1096, signal_1095, signal_1094, signal_404}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_394 ( .a ({signal_1084, signal_1083, signal_1082, signal_400}), .b ({signal_1114, signal_1113, signal_1112, signal_410}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_395 ( .a ({signal_1087, signal_1086, signal_1085, signal_401}), .b ({signal_1117, signal_1116, signal_1115, signal_411}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_400 ( .a ({signal_1090, signal_1089, signal_1088, signal_402}), .b ({signal_1132, signal_1131, signal_1130, signal_416}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_401 ( .a ({signal_1093, signal_1092, signal_1091, signal_403}), .b ({signal_1135, signal_1134, signal_1133, signal_417}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_402 ( .a ({signal_1096, signal_1095, signal_1094, signal_404}), .b ({signal_1138, signal_1137, signal_1136, signal_418}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_404 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1075, signal_1074, signal_1073, signal_397}), .clk ( clk ), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({signal_1144, signal_1143, signal_1142, signal_419}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_407 ( .a ({signal_1144, signal_1143, signal_1142, signal_419}), .b ({signal_1153, signal_1152, signal_1151, signal_422}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_412 ( .a ({1'b0, 1'b0, 1'b0, signal_2260}), .b ({signal_1123, signal_1122, signal_1121, signal_413}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({signal_1168, signal_1167, signal_1166, signal_425}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_413 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1126, signal_1125, signal_1124, signal_414}), .clk ( clk ), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_1171, signal_1170, signal_1169, signal_426}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_414 ( .a ({1'b0, 1'b0, 1'b0, signal_2260}), .b ({signal_1120, signal_1119, signal_1118, signal_412}), .clk ( clk ), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({signal_1174, signal_1173, signal_1172, signal_427}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_415 ( .a ({1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1129, signal_1128, signal_1127, signal_415}), .clk ( clk ), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({signal_1177, signal_1176, signal_1175, signal_428}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_416 ( .a ({signal_1168, signal_1167, signal_1166, signal_425}), .b ({signal_1180, signal_1179, signal_1178, signal_429}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_417 ( .a ({signal_1171, signal_1170, signal_1169, signal_426}), .b ({signal_1183, signal_1182, signal_1181, signal_430}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_418 ( .a ({signal_1174, signal_1173, signal_1172, signal_427}), .b ({signal_1186, signal_1185, signal_1184, signal_431}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_419 ( .a ({signal_1177, signal_1176, signal_1175, signal_428}), .b ({signal_1189, signal_1188, signal_1187, signal_432}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_421 ( .a ({1'b0, 1'b0, 1'b0, signal_2260}), .b ({signal_1156, signal_1155, signal_1154, signal_423}), .clk ( clk ), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({signal_1195, signal_1194, signal_1193, signal_433}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_422 ( .a ({1'b0, 1'b0, 1'b0, signal_2260}), .b ({signal_1159, signal_1158, signal_1157, signal_424}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({signal_1198, signal_1197, signal_1196, signal_434}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_423 ( .a ({signal_1195, signal_1194, signal_1193, signal_433}), .b ({signal_1201, signal_1200, signal_1199, signal_435}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_424 ( .a ({signal_1198, signal_1197, signal_1196, signal_434}), .b ({signal_1204, signal_1203, signal_1202, signal_436}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_403 ( .a ({signal_1054, signal_1053, signal_1052, signal_390}), .b ({signal_1078, signal_1077, signal_1076, signal_398}), .clk ( clk ), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_1141, signal_1140, signal_1139, signal_167}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_410 ( .a ({signal_1114, signal_1113, signal_1112, signal_410}), .b ({signal_1117, signal_1116, signal_1115, signal_411}), .clk ( clk ), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({signal_1162, signal_1161, signal_1160, signal_160}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_411 ( .a ({signal_1135, signal_1134, signal_1133, signal_417}), .b ({signal_1138, signal_1137, signal_1136, signal_418}), .clk ( clk ), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({signal_1165, signal_1164, signal_1163, signal_166}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_420 ( .a ({signal_1132, signal_1131, signal_1130, signal_416}), .b ({signal_1153, signal_1152, signal_1151, signal_422}), .clk ( clk ), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({signal_1192, signal_1191, signal_1190, signal_163}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_425 ( .a ({signal_1180, signal_1179, signal_1178, signal_429}), .b ({signal_1183, signal_1182, signal_1181, signal_430}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({signal_1207, signal_1206, signal_1205, signal_164}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_426 ( .a ({signal_1186, signal_1185, signal_1184, signal_431}), .b ({signal_1189, signal_1188, signal_1187, signal_432}), .clk ( clk ), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_1210, signal_1209, signal_1208, signal_165}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_427 ( .a ({signal_1201, signal_1200, signal_1199, signal_435}), .b ({signal_1081, signal_1080, signal_1079, signal_399}), .clk ( clk ), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({signal_1213, signal_1212, signal_1211, signal_161}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_428 ( .a ({signal_1204, signal_1203, signal_1202, signal_436}), .b ({signal_1057, signal_1056, signal_1055, signal_391}), .clk ( clk ), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({signal_1216, signal_1215, signal_1214, signal_162}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_1162, signal_1161, signal_1160, signal_160}), .Q ({Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_1213, signal_1212, signal_1211, signal_161}), .Q ({Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_1216, signal_1215, signal_1214, signal_162}), .Q ({Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_1192, signal_1191, signal_1190, signal_163}), .Q ({Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_4 ( .clk ( clk ), .D ({signal_1207, signal_1206, signal_1205, signal_164}), .Q ({Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_5 ( .clk ( clk ), .D ({signal_1210, signal_1209, signal_1208, signal_165}), .Q ({Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_6 ( .clk ( clk ), .D ({signal_1165, signal_1164, signal_1163, signal_166}), .Q ({Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_7 ( .clk ( clk ), .D ({signal_1141, signal_1140, signal_1139, signal_167}), .Q ({Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
