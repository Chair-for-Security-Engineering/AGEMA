/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC1_Pipeline_d3 (X_s0, clk, X_s1, X_s2, X_s3, Fresh, Y_s0, Y_s1, Y_s2, Y_s3);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [339:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    wire T1 ;
    wire T2 ;
    wire T3 ;
    wire T4 ;
    wire T5 ;
    wire T6 ;
    wire T7 ;
    wire T8 ;
    wire T9 ;
    wire T10 ;
    wire T11 ;
    wire T12 ;
    wire T13 ;
    wire T14 ;
    wire T15 ;
    wire T16 ;
    wire T17 ;
    wire T18 ;
    wire T19 ;
    wire T20 ;
    wire T21 ;
    wire T22 ;
    wire T23 ;
    wire T24 ;
    wire T25 ;
    wire T26 ;
    wire T27 ;
    wire M1 ;
    wire M2 ;
    wire M3 ;
    wire M4 ;
    wire M5 ;
    wire M6 ;
    wire M7 ;
    wire M8 ;
    wire M9 ;
    wire M10 ;
    wire M11 ;
    wire M12 ;
    wire M13 ;
    wire M14 ;
    wire M15 ;
    wire M16 ;
    wire M17 ;
    wire M18 ;
    wire M19 ;
    wire M20 ;
    wire M21 ;
    wire M22 ;
    wire M23 ;
    wire M24 ;
    wire M25 ;
    wire M26 ;
    wire M27 ;
    wire M28 ;
    wire M29 ;
    wire M30 ;
    wire M31 ;
    wire M32 ;
    wire M33 ;
    wire M34 ;
    wire M35 ;
    wire M36 ;
    wire M37 ;
    wire M38 ;
    wire M39 ;
    wire M40 ;
    wire M41 ;
    wire M42 ;
    wire M43 ;
    wire M44 ;
    wire M45 ;
    wire M46 ;
    wire M47 ;
    wire M48 ;
    wire M49 ;
    wire M50 ;
    wire M51 ;
    wire M52 ;
    wire M53 ;
    wire M54 ;
    wire M55 ;
    wire M56 ;
    wire M57 ;
    wire M58 ;
    wire M59 ;
    wire M60 ;
    wire M61 ;
    wire M62 ;
    wire M63 ;
    wire L0 ;
    wire L1 ;
    wire L2 ;
    wire L3 ;
    wire L4 ;
    wire L5 ;
    wire L6 ;
    wire L7 ;
    wire L8 ;
    wire L9 ;
    wire L10 ;
    wire L11 ;
    wire L12 ;
    wire L13 ;
    wire L14 ;
    wire L15 ;
    wire L16 ;
    wire L17 ;
    wire L18 ;
    wire L19 ;
    wire L20 ;
    wire L21 ;
    wire L22 ;
    wire L23 ;
    wire L24 ;
    wire L25 ;
    wire L26 ;
    wire L27 ;
    wire L28 ;
    wire L29 ;
    wire [7:0] O ;
    wire new_AGEMA_signal_157 ;
    wire new_AGEMA_signal_158 ;
    wire new_AGEMA_signal_159 ;
    wire new_AGEMA_signal_163 ;
    wire new_AGEMA_signal_164 ;
    wire new_AGEMA_signal_165 ;
    wire new_AGEMA_signal_169 ;
    wire new_AGEMA_signal_170 ;
    wire new_AGEMA_signal_171 ;
    wire new_AGEMA_signal_172 ;
    wire new_AGEMA_signal_173 ;
    wire new_AGEMA_signal_174 ;
    wire new_AGEMA_signal_178 ;
    wire new_AGEMA_signal_179 ;
    wire new_AGEMA_signal_180 ;
    wire new_AGEMA_signal_187 ;
    wire new_AGEMA_signal_188 ;
    wire new_AGEMA_signal_189 ;
    wire new_AGEMA_signal_190 ;
    wire new_AGEMA_signal_191 ;
    wire new_AGEMA_signal_192 ;
    wire new_AGEMA_signal_193 ;
    wire new_AGEMA_signal_194 ;
    wire new_AGEMA_signal_195 ;
    wire new_AGEMA_signal_199 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_206 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_212 ;
    wire new_AGEMA_signal_213 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_423 ;
    wire new_AGEMA_signal_424 ;
    wire new_AGEMA_signal_425 ;
    wire new_AGEMA_signal_426 ;
    wire new_AGEMA_signal_427 ;
    wire new_AGEMA_signal_428 ;
    wire new_AGEMA_signal_429 ;
    wire new_AGEMA_signal_430 ;
    wire new_AGEMA_signal_431 ;
    wire new_AGEMA_signal_432 ;
    wire new_AGEMA_signal_433 ;
    wire new_AGEMA_signal_434 ;
    wire new_AGEMA_signal_435 ;
    wire new_AGEMA_signal_436 ;
    wire new_AGEMA_signal_437 ;
    wire new_AGEMA_signal_438 ;
    wire new_AGEMA_signal_439 ;
    wire new_AGEMA_signal_440 ;
    wire new_AGEMA_signal_441 ;
    wire new_AGEMA_signal_442 ;
    wire new_AGEMA_signal_443 ;
    wire new_AGEMA_signal_444 ;
    wire new_AGEMA_signal_445 ;
    wire new_AGEMA_signal_446 ;
    wire new_AGEMA_signal_447 ;
    wire new_AGEMA_signal_448 ;
    wire new_AGEMA_signal_449 ;
    wire new_AGEMA_signal_450 ;
    wire new_AGEMA_signal_451 ;
    wire new_AGEMA_signal_452 ;
    wire new_AGEMA_signal_453 ;
    wire new_AGEMA_signal_454 ;
    wire new_AGEMA_signal_455 ;
    wire new_AGEMA_signal_456 ;
    wire new_AGEMA_signal_457 ;
    wire new_AGEMA_signal_458 ;
    wire new_AGEMA_signal_459 ;
    wire new_AGEMA_signal_460 ;
    wire new_AGEMA_signal_461 ;
    wire new_AGEMA_signal_462 ;
    wire new_AGEMA_signal_463 ;
    wire new_AGEMA_signal_464 ;
    wire new_AGEMA_signal_465 ;
    wire new_AGEMA_signal_466 ;
    wire new_AGEMA_signal_467 ;
    wire new_AGEMA_signal_468 ;
    wire new_AGEMA_signal_469 ;
    wire new_AGEMA_signal_470 ;
    wire new_AGEMA_signal_471 ;
    wire new_AGEMA_signal_472 ;
    wire new_AGEMA_signal_473 ;
    wire new_AGEMA_signal_474 ;
    wire new_AGEMA_signal_475 ;
    wire new_AGEMA_signal_476 ;
    wire new_AGEMA_signal_477 ;
    wire new_AGEMA_signal_478 ;
    wire new_AGEMA_signal_479 ;
    wire new_AGEMA_signal_480 ;
    wire new_AGEMA_signal_481 ;
    wire new_AGEMA_signal_482 ;
    wire new_AGEMA_signal_483 ;
    wire new_AGEMA_signal_484 ;
    wire new_AGEMA_signal_485 ;
    wire new_AGEMA_signal_486 ;
    wire new_AGEMA_signal_487 ;
    wire new_AGEMA_signal_488 ;
    wire new_AGEMA_signal_489 ;
    wire new_AGEMA_signal_490 ;
    wire new_AGEMA_signal_491 ;
    wire new_AGEMA_signal_492 ;
    wire new_AGEMA_signal_493 ;
    wire new_AGEMA_signal_494 ;
    wire new_AGEMA_signal_495 ;
    wire new_AGEMA_signal_496 ;
    wire new_AGEMA_signal_497 ;
    wire new_AGEMA_signal_498 ;
    wire new_AGEMA_signal_499 ;
    wire new_AGEMA_signal_500 ;
    wire new_AGEMA_signal_501 ;
    wire new_AGEMA_signal_502 ;
    wire new_AGEMA_signal_503 ;
    wire new_AGEMA_signal_504 ;
    wire new_AGEMA_signal_505 ;
    wire new_AGEMA_signal_506 ;
    wire new_AGEMA_signal_507 ;
    wire new_AGEMA_signal_508 ;
    wire new_AGEMA_signal_509 ;
    wire new_AGEMA_signal_510 ;
    wire new_AGEMA_signal_511 ;
    wire new_AGEMA_signal_512 ;
    wire new_AGEMA_signal_513 ;
    wire new_AGEMA_signal_514 ;
    wire new_AGEMA_signal_515 ;
    wire new_AGEMA_signal_516 ;
    wire new_AGEMA_signal_517 ;
    wire new_AGEMA_signal_518 ;
    wire new_AGEMA_signal_519 ;
    wire new_AGEMA_signal_520 ;
    wire new_AGEMA_signal_521 ;
    wire new_AGEMA_signal_522 ;
    wire new_AGEMA_signal_523 ;
    wire new_AGEMA_signal_524 ;
    wire new_AGEMA_signal_525 ;
    wire new_AGEMA_signal_526 ;
    wire new_AGEMA_signal_527 ;
    wire new_AGEMA_signal_528 ;
    wire new_AGEMA_signal_529 ;
    wire new_AGEMA_signal_530 ;
    wire new_AGEMA_signal_531 ;
    wire new_AGEMA_signal_532 ;
    wire new_AGEMA_signal_533 ;
    wire new_AGEMA_signal_534 ;
    wire new_AGEMA_signal_535 ;
    wire new_AGEMA_signal_536 ;
    wire new_AGEMA_signal_537 ;
    wire new_AGEMA_signal_538 ;
    wire new_AGEMA_signal_539 ;
    wire new_AGEMA_signal_540 ;
    wire new_AGEMA_signal_541 ;
    wire new_AGEMA_signal_542 ;
    wire new_AGEMA_signal_543 ;
    wire new_AGEMA_signal_544 ;
    wire new_AGEMA_signal_545 ;
    wire new_AGEMA_signal_546 ;
    wire new_AGEMA_signal_547 ;
    wire new_AGEMA_signal_548 ;
    wire new_AGEMA_signal_549 ;
    wire new_AGEMA_signal_550 ;
    wire new_AGEMA_signal_551 ;
    wire new_AGEMA_signal_552 ;
    wire new_AGEMA_signal_553 ;
    wire new_AGEMA_signal_554 ;
    wire new_AGEMA_signal_555 ;
    wire new_AGEMA_signal_556 ;
    wire new_AGEMA_signal_557 ;
    wire new_AGEMA_signal_558 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_924 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_928 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_930 ;
    wire new_AGEMA_signal_931 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_934 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_939 ;
    wire new_AGEMA_signal_940 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_942 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;

    /* cells in depth 0 */
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T1_U1 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T2_U1 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_165, new_AGEMA_signal_164, new_AGEMA_signal_163, T2}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T3_U1 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_171, new_AGEMA_signal_170, new_AGEMA_signal_169, T3}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T4_U1 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_174, new_AGEMA_signal_173, new_AGEMA_signal_172, T4}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T5_U1 ( .a ({X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_180, new_AGEMA_signal_179, new_AGEMA_signal_178, T5}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T6_U1 ( .a ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}), .b ({new_AGEMA_signal_180, new_AGEMA_signal_179, new_AGEMA_signal_178, T5}), .c ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T7_U1 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .c ({new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T7}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T8_U1 ( .a ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}), .c ({new_AGEMA_signal_231, new_AGEMA_signal_230, new_AGEMA_signal_229, T8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T9_U1 ( .a ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T7}), .c ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, T9}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T10_U1 ( .a ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}), .b ({new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T7}), .c ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, T10}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T11_U1 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_192, new_AGEMA_signal_191, new_AGEMA_signal_190, T11}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T12_U1 ( .a ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_195, new_AGEMA_signal_194, new_AGEMA_signal_193, T12}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T13_U1 ( .a ({new_AGEMA_signal_171, new_AGEMA_signal_170, new_AGEMA_signal_169, T3}), .b ({new_AGEMA_signal_174, new_AGEMA_signal_173, new_AGEMA_signal_172, T4}), .c ({new_AGEMA_signal_213, new_AGEMA_signal_212, new_AGEMA_signal_211, T13}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T14_U1 ( .a ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}), .b ({new_AGEMA_signal_192, new_AGEMA_signal_191, new_AGEMA_signal_190, T11}), .c ({new_AGEMA_signal_237, new_AGEMA_signal_236, new_AGEMA_signal_235, T14}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T15_U1 ( .a ({new_AGEMA_signal_180, new_AGEMA_signal_179, new_AGEMA_signal_178, T5}), .b ({new_AGEMA_signal_192, new_AGEMA_signal_191, new_AGEMA_signal_190, T11}), .c ({new_AGEMA_signal_216, new_AGEMA_signal_215, new_AGEMA_signal_214, T15}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T16_U1 ( .a ({new_AGEMA_signal_180, new_AGEMA_signal_179, new_AGEMA_signal_178, T5}), .b ({new_AGEMA_signal_195, new_AGEMA_signal_194, new_AGEMA_signal_193, T12}), .c ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, T16}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T17_U1 ( .a ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, T9}), .b ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, T16}), .c ({new_AGEMA_signal_240, new_AGEMA_signal_239, new_AGEMA_signal_238, T17}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T18_U1 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T18}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T19_U1 ( .a ({new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T7}), .b ({new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T18}), .c ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, T19}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T20_U1 ( .a ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}), .b ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, T19}), .c ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, T20}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T21_U1 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_204, new_AGEMA_signal_203, new_AGEMA_signal_202, T21}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T22_U1 ( .a ({new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T7}), .b ({new_AGEMA_signal_204, new_AGEMA_signal_203, new_AGEMA_signal_202, T21}), .c ({new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T22}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T23_U1 ( .a ({new_AGEMA_signal_165, new_AGEMA_signal_164, new_AGEMA_signal_163, T2}), .b ({new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T22}), .c ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, T23}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T24_U1 ( .a ({new_AGEMA_signal_165, new_AGEMA_signal_164, new_AGEMA_signal_163, T2}), .b ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, T10}), .c ({new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, T24}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T25_U1 ( .a ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, T20}), .b ({new_AGEMA_signal_240, new_AGEMA_signal_239, new_AGEMA_signal_238, T17}), .c ({new_AGEMA_signal_273, new_AGEMA_signal_272, new_AGEMA_signal_271, T25}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T26_U1 ( .a ({new_AGEMA_signal_171, new_AGEMA_signal_170, new_AGEMA_signal_169, T3}), .b ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, T16}), .c ({new_AGEMA_signal_249, new_AGEMA_signal_248, new_AGEMA_signal_247, T26}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_T27_U1 ( .a ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}), .b ({new_AGEMA_signal_195, new_AGEMA_signal_194, new_AGEMA_signal_193, T12}), .c ({new_AGEMA_signal_228, new_AGEMA_signal_227, new_AGEMA_signal_226, T27}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_136 ( .C (clk), .D (T14), .Q (new_AGEMA_signal_923) ) ;
    buf_clk new_AGEMA_reg_buffer_138 ( .C (clk), .D (new_AGEMA_signal_235), .Q (new_AGEMA_signal_925) ) ;
    buf_clk new_AGEMA_reg_buffer_140 ( .C (clk), .D (new_AGEMA_signal_236), .Q (new_AGEMA_signal_927) ) ;
    buf_clk new_AGEMA_reg_buffer_142 ( .C (clk), .D (new_AGEMA_signal_237), .Q (new_AGEMA_signal_929) ) ;
    buf_clk new_AGEMA_reg_buffer_144 ( .C (clk), .D (T26), .Q (new_AGEMA_signal_931) ) ;
    buf_clk new_AGEMA_reg_buffer_146 ( .C (clk), .D (new_AGEMA_signal_247), .Q (new_AGEMA_signal_933) ) ;
    buf_clk new_AGEMA_reg_buffer_148 ( .C (clk), .D (new_AGEMA_signal_248), .Q (new_AGEMA_signal_935) ) ;
    buf_clk new_AGEMA_reg_buffer_150 ( .C (clk), .D (new_AGEMA_signal_249), .Q (new_AGEMA_signal_937) ) ;
    buf_clk new_AGEMA_reg_buffer_152 ( .C (clk), .D (T24), .Q (new_AGEMA_signal_939) ) ;
    buf_clk new_AGEMA_reg_buffer_154 ( .C (clk), .D (new_AGEMA_signal_268), .Q (new_AGEMA_signal_941) ) ;
    buf_clk new_AGEMA_reg_buffer_156 ( .C (clk), .D (new_AGEMA_signal_269), .Q (new_AGEMA_signal_943) ) ;
    buf_clk new_AGEMA_reg_buffer_158 ( .C (clk), .D (new_AGEMA_signal_270), .Q (new_AGEMA_signal_945) ) ;
    buf_clk new_AGEMA_reg_buffer_160 ( .C (clk), .D (T25), .Q (new_AGEMA_signal_947) ) ;
    buf_clk new_AGEMA_reg_buffer_162 ( .C (clk), .D (new_AGEMA_signal_271), .Q (new_AGEMA_signal_949) ) ;
    buf_clk new_AGEMA_reg_buffer_164 ( .C (clk), .D (new_AGEMA_signal_272), .Q (new_AGEMA_signal_951) ) ;
    buf_clk new_AGEMA_reg_buffer_166 ( .C (clk), .D (new_AGEMA_signal_273), .Q (new_AGEMA_signal_953) ) ;
    buf_clk new_AGEMA_reg_buffer_232 ( .C (clk), .D (T6), .Q (new_AGEMA_signal_1019) ) ;
    buf_clk new_AGEMA_reg_buffer_238 ( .C (clk), .D (new_AGEMA_signal_205), .Q (new_AGEMA_signal_1025) ) ;
    buf_clk new_AGEMA_reg_buffer_244 ( .C (clk), .D (new_AGEMA_signal_206), .Q (new_AGEMA_signal_1031) ) ;
    buf_clk new_AGEMA_reg_buffer_250 ( .C (clk), .D (new_AGEMA_signal_207), .Q (new_AGEMA_signal_1037) ) ;
    buf_clk new_AGEMA_reg_buffer_256 ( .C (clk), .D (T8), .Q (new_AGEMA_signal_1043) ) ;
    buf_clk new_AGEMA_reg_buffer_262 ( .C (clk), .D (new_AGEMA_signal_229), .Q (new_AGEMA_signal_1049) ) ;
    buf_clk new_AGEMA_reg_buffer_268 ( .C (clk), .D (new_AGEMA_signal_230), .Q (new_AGEMA_signal_1055) ) ;
    buf_clk new_AGEMA_reg_buffer_274 ( .C (clk), .D (new_AGEMA_signal_231), .Q (new_AGEMA_signal_1061) ) ;
    buf_clk new_AGEMA_reg_buffer_280 ( .C (clk), .D (X_s0[0]), .Q (new_AGEMA_signal_1067) ) ;
    buf_clk new_AGEMA_reg_buffer_286 ( .C (clk), .D (X_s1[0]), .Q (new_AGEMA_signal_1073) ) ;
    buf_clk new_AGEMA_reg_buffer_292 ( .C (clk), .D (X_s2[0]), .Q (new_AGEMA_signal_1079) ) ;
    buf_clk new_AGEMA_reg_buffer_298 ( .C (clk), .D (X_s3[0]), .Q (new_AGEMA_signal_1085) ) ;
    buf_clk new_AGEMA_reg_buffer_304 ( .C (clk), .D (T16), .Q (new_AGEMA_signal_1091) ) ;
    buf_clk new_AGEMA_reg_buffer_310 ( .C (clk), .D (new_AGEMA_signal_217), .Q (new_AGEMA_signal_1097) ) ;
    buf_clk new_AGEMA_reg_buffer_316 ( .C (clk), .D (new_AGEMA_signal_218), .Q (new_AGEMA_signal_1103) ) ;
    buf_clk new_AGEMA_reg_buffer_322 ( .C (clk), .D (new_AGEMA_signal_219), .Q (new_AGEMA_signal_1109) ) ;
    buf_clk new_AGEMA_reg_buffer_328 ( .C (clk), .D (T9), .Q (new_AGEMA_signal_1115) ) ;
    buf_clk new_AGEMA_reg_buffer_334 ( .C (clk), .D (new_AGEMA_signal_208), .Q (new_AGEMA_signal_1121) ) ;
    buf_clk new_AGEMA_reg_buffer_340 ( .C (clk), .D (new_AGEMA_signal_209), .Q (new_AGEMA_signal_1127) ) ;
    buf_clk new_AGEMA_reg_buffer_346 ( .C (clk), .D (new_AGEMA_signal_210), .Q (new_AGEMA_signal_1133) ) ;
    buf_clk new_AGEMA_reg_buffer_352 ( .C (clk), .D (T17), .Q (new_AGEMA_signal_1139) ) ;
    buf_clk new_AGEMA_reg_buffer_358 ( .C (clk), .D (new_AGEMA_signal_238), .Q (new_AGEMA_signal_1145) ) ;
    buf_clk new_AGEMA_reg_buffer_364 ( .C (clk), .D (new_AGEMA_signal_239), .Q (new_AGEMA_signal_1151) ) ;
    buf_clk new_AGEMA_reg_buffer_370 ( .C (clk), .D (new_AGEMA_signal_240), .Q (new_AGEMA_signal_1157) ) ;
    buf_clk new_AGEMA_reg_buffer_376 ( .C (clk), .D (T15), .Q (new_AGEMA_signal_1163) ) ;
    buf_clk new_AGEMA_reg_buffer_382 ( .C (clk), .D (new_AGEMA_signal_214), .Q (new_AGEMA_signal_1169) ) ;
    buf_clk new_AGEMA_reg_buffer_388 ( .C (clk), .D (new_AGEMA_signal_215), .Q (new_AGEMA_signal_1175) ) ;
    buf_clk new_AGEMA_reg_buffer_394 ( .C (clk), .D (new_AGEMA_signal_216), .Q (new_AGEMA_signal_1181) ) ;
    buf_clk new_AGEMA_reg_buffer_400 ( .C (clk), .D (T27), .Q (new_AGEMA_signal_1187) ) ;
    buf_clk new_AGEMA_reg_buffer_406 ( .C (clk), .D (new_AGEMA_signal_226), .Q (new_AGEMA_signal_1193) ) ;
    buf_clk new_AGEMA_reg_buffer_412 ( .C (clk), .D (new_AGEMA_signal_227), .Q (new_AGEMA_signal_1199) ) ;
    buf_clk new_AGEMA_reg_buffer_418 ( .C (clk), .D (new_AGEMA_signal_228), .Q (new_AGEMA_signal_1205) ) ;
    buf_clk new_AGEMA_reg_buffer_424 ( .C (clk), .D (T10), .Q (new_AGEMA_signal_1211) ) ;
    buf_clk new_AGEMA_reg_buffer_430 ( .C (clk), .D (new_AGEMA_signal_232), .Q (new_AGEMA_signal_1217) ) ;
    buf_clk new_AGEMA_reg_buffer_436 ( .C (clk), .D (new_AGEMA_signal_233), .Q (new_AGEMA_signal_1223) ) ;
    buf_clk new_AGEMA_reg_buffer_442 ( .C (clk), .D (new_AGEMA_signal_234), .Q (new_AGEMA_signal_1229) ) ;
    buf_clk new_AGEMA_reg_buffer_448 ( .C (clk), .D (T13), .Q (new_AGEMA_signal_1235) ) ;
    buf_clk new_AGEMA_reg_buffer_454 ( .C (clk), .D (new_AGEMA_signal_211), .Q (new_AGEMA_signal_1241) ) ;
    buf_clk new_AGEMA_reg_buffer_460 ( .C (clk), .D (new_AGEMA_signal_212), .Q (new_AGEMA_signal_1247) ) ;
    buf_clk new_AGEMA_reg_buffer_466 ( .C (clk), .D (new_AGEMA_signal_213), .Q (new_AGEMA_signal_1253) ) ;
    buf_clk new_AGEMA_reg_buffer_472 ( .C (clk), .D (T23), .Q (new_AGEMA_signal_1259) ) ;
    buf_clk new_AGEMA_reg_buffer_478 ( .C (clk), .D (new_AGEMA_signal_244), .Q (new_AGEMA_signal_1265) ) ;
    buf_clk new_AGEMA_reg_buffer_484 ( .C (clk), .D (new_AGEMA_signal_245), .Q (new_AGEMA_signal_1271) ) ;
    buf_clk new_AGEMA_reg_buffer_490 ( .C (clk), .D (new_AGEMA_signal_246), .Q (new_AGEMA_signal_1277) ) ;
    buf_clk new_AGEMA_reg_buffer_496 ( .C (clk), .D (T19), .Q (new_AGEMA_signal_1283) ) ;
    buf_clk new_AGEMA_reg_buffer_502 ( .C (clk), .D (new_AGEMA_signal_220), .Q (new_AGEMA_signal_1289) ) ;
    buf_clk new_AGEMA_reg_buffer_508 ( .C (clk), .D (new_AGEMA_signal_221), .Q (new_AGEMA_signal_1295) ) ;
    buf_clk new_AGEMA_reg_buffer_514 ( .C (clk), .D (new_AGEMA_signal_222), .Q (new_AGEMA_signal_1301) ) ;
    buf_clk new_AGEMA_reg_buffer_520 ( .C (clk), .D (T3), .Q (new_AGEMA_signal_1307) ) ;
    buf_clk new_AGEMA_reg_buffer_526 ( .C (clk), .D (new_AGEMA_signal_169), .Q (new_AGEMA_signal_1313) ) ;
    buf_clk new_AGEMA_reg_buffer_532 ( .C (clk), .D (new_AGEMA_signal_170), .Q (new_AGEMA_signal_1319) ) ;
    buf_clk new_AGEMA_reg_buffer_538 ( .C (clk), .D (new_AGEMA_signal_171), .Q (new_AGEMA_signal_1325) ) ;
    buf_clk new_AGEMA_reg_buffer_544 ( .C (clk), .D (T22), .Q (new_AGEMA_signal_1331) ) ;
    buf_clk new_AGEMA_reg_buffer_550 ( .C (clk), .D (new_AGEMA_signal_223), .Q (new_AGEMA_signal_1337) ) ;
    buf_clk new_AGEMA_reg_buffer_556 ( .C (clk), .D (new_AGEMA_signal_224), .Q (new_AGEMA_signal_1343) ) ;
    buf_clk new_AGEMA_reg_buffer_562 ( .C (clk), .D (new_AGEMA_signal_225), .Q (new_AGEMA_signal_1349) ) ;
    buf_clk new_AGEMA_reg_buffer_568 ( .C (clk), .D (T20), .Q (new_AGEMA_signal_1355) ) ;
    buf_clk new_AGEMA_reg_buffer_574 ( .C (clk), .D (new_AGEMA_signal_241), .Q (new_AGEMA_signal_1361) ) ;
    buf_clk new_AGEMA_reg_buffer_580 ( .C (clk), .D (new_AGEMA_signal_242), .Q (new_AGEMA_signal_1367) ) ;
    buf_clk new_AGEMA_reg_buffer_586 ( .C (clk), .D (new_AGEMA_signal_243), .Q (new_AGEMA_signal_1373) ) ;
    buf_clk new_AGEMA_reg_buffer_592 ( .C (clk), .D (T1), .Q (new_AGEMA_signal_1379) ) ;
    buf_clk new_AGEMA_reg_buffer_598 ( .C (clk), .D (new_AGEMA_signal_157), .Q (new_AGEMA_signal_1385) ) ;
    buf_clk new_AGEMA_reg_buffer_604 ( .C (clk), .D (new_AGEMA_signal_158), .Q (new_AGEMA_signal_1391) ) ;
    buf_clk new_AGEMA_reg_buffer_610 ( .C (clk), .D (new_AGEMA_signal_159), .Q (new_AGEMA_signal_1397) ) ;
    buf_clk new_AGEMA_reg_buffer_616 ( .C (clk), .D (T4), .Q (new_AGEMA_signal_1403) ) ;
    buf_clk new_AGEMA_reg_buffer_622 ( .C (clk), .D (new_AGEMA_signal_172), .Q (new_AGEMA_signal_1409) ) ;
    buf_clk new_AGEMA_reg_buffer_628 ( .C (clk), .D (new_AGEMA_signal_173), .Q (new_AGEMA_signal_1415) ) ;
    buf_clk new_AGEMA_reg_buffer_634 ( .C (clk), .D (new_AGEMA_signal_174), .Q (new_AGEMA_signal_1421) ) ;
    buf_clk new_AGEMA_reg_buffer_640 ( .C (clk), .D (T2), .Q (new_AGEMA_signal_1427) ) ;
    buf_clk new_AGEMA_reg_buffer_646 ( .C (clk), .D (new_AGEMA_signal_163), .Q (new_AGEMA_signal_1433) ) ;
    buf_clk new_AGEMA_reg_buffer_652 ( .C (clk), .D (new_AGEMA_signal_164), .Q (new_AGEMA_signal_1439) ) ;
    buf_clk new_AGEMA_reg_buffer_658 ( .C (clk), .D (new_AGEMA_signal_165), .Q (new_AGEMA_signal_1445) ) ;

    /* cells in depth 2 */
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M1_U1 ( .ina ({new_AGEMA_signal_213, new_AGEMA_signal_212, new_AGEMA_signal_211, T13}), .inb ({new_AGEMA_signal_207, new_AGEMA_signal_206, new_AGEMA_signal_205, T6}), .clk (clk), .rnd ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .outt ({new_AGEMA_signal_252, new_AGEMA_signal_251, new_AGEMA_signal_250, M1}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M2_U1 ( .ina ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, T23}), .inb ({new_AGEMA_signal_231, new_AGEMA_signal_230, new_AGEMA_signal_229, T8}), .clk (clk), .rnd ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .outt ({new_AGEMA_signal_276, new_AGEMA_signal_275, new_AGEMA_signal_274, M2}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M3_U1 ( .a ({new_AGEMA_signal_930, new_AGEMA_signal_928, new_AGEMA_signal_926, new_AGEMA_signal_924}), .b ({new_AGEMA_signal_252, new_AGEMA_signal_251, new_AGEMA_signal_250, M1}), .c ({new_AGEMA_signal_279, new_AGEMA_signal_278, new_AGEMA_signal_277, M3}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M4_U1 ( .ina ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, T19}), .inb ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .clk (clk), .rnd ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .outt ({new_AGEMA_signal_255, new_AGEMA_signal_254, new_AGEMA_signal_253, M4}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M5_U1 ( .a ({new_AGEMA_signal_255, new_AGEMA_signal_254, new_AGEMA_signal_253, M4}), .b ({new_AGEMA_signal_252, new_AGEMA_signal_251, new_AGEMA_signal_250, M1}), .c ({new_AGEMA_signal_282, new_AGEMA_signal_281, new_AGEMA_signal_280, M5}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M6_U1 ( .ina ({new_AGEMA_signal_171, new_AGEMA_signal_170, new_AGEMA_signal_169, T3}), .inb ({new_AGEMA_signal_219, new_AGEMA_signal_218, new_AGEMA_signal_217, T16}), .clk (clk), .rnd ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .outt ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, M6}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M7_U1 ( .ina ({new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T22}), .inb ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, T9}), .clk (clk), .rnd ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .outt ({new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, M7}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M8_U1 ( .a ({new_AGEMA_signal_938, new_AGEMA_signal_936, new_AGEMA_signal_934, new_AGEMA_signal_932}), .b ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, M6}), .c ({new_AGEMA_signal_285, new_AGEMA_signal_284, new_AGEMA_signal_283, M8}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M9_U1 ( .ina ({new_AGEMA_signal_243, new_AGEMA_signal_242, new_AGEMA_signal_241, T20}), .inb ({new_AGEMA_signal_240, new_AGEMA_signal_239, new_AGEMA_signal_238, T17}), .clk (clk), .rnd ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .outt ({new_AGEMA_signal_288, new_AGEMA_signal_287, new_AGEMA_signal_286, M9}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M10_U1 ( .a ({new_AGEMA_signal_288, new_AGEMA_signal_287, new_AGEMA_signal_286, M9}), .b ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, M6}), .c ({new_AGEMA_signal_297, new_AGEMA_signal_296, new_AGEMA_signal_295, M10}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M11_U1 ( .ina ({new_AGEMA_signal_159, new_AGEMA_signal_158, new_AGEMA_signal_157, T1}), .inb ({new_AGEMA_signal_216, new_AGEMA_signal_215, new_AGEMA_signal_214, T15}), .clk (clk), .rnd ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .outt ({new_AGEMA_signal_264, new_AGEMA_signal_263, new_AGEMA_signal_262, M11}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M12_U1 ( .ina ({new_AGEMA_signal_174, new_AGEMA_signal_173, new_AGEMA_signal_172, T4}), .inb ({new_AGEMA_signal_228, new_AGEMA_signal_227, new_AGEMA_signal_226, T27}), .clk (clk), .rnd ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .outt ({new_AGEMA_signal_267, new_AGEMA_signal_266, new_AGEMA_signal_265, M12}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M13_U1 ( .a ({new_AGEMA_signal_267, new_AGEMA_signal_266, new_AGEMA_signal_265, M12}), .b ({new_AGEMA_signal_264, new_AGEMA_signal_263, new_AGEMA_signal_262, M11}), .c ({new_AGEMA_signal_291, new_AGEMA_signal_290, new_AGEMA_signal_289, M13}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M14_U1 ( .ina ({new_AGEMA_signal_165, new_AGEMA_signal_164, new_AGEMA_signal_163, T2}), .inb ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, T10}), .clk (clk), .rnd ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .outt ({new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, M14}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M15_U1 ( .a ({new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, M14}), .b ({new_AGEMA_signal_264, new_AGEMA_signal_263, new_AGEMA_signal_262, M11}), .c ({new_AGEMA_signal_300, new_AGEMA_signal_299, new_AGEMA_signal_298, M15}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M16_U1 ( .a ({new_AGEMA_signal_279, new_AGEMA_signal_278, new_AGEMA_signal_277, M3}), .b ({new_AGEMA_signal_276, new_AGEMA_signal_275, new_AGEMA_signal_274, M2}), .c ({new_AGEMA_signal_303, new_AGEMA_signal_302, new_AGEMA_signal_301, M16}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M17_U1 ( .a ({new_AGEMA_signal_282, new_AGEMA_signal_281, new_AGEMA_signal_280, M5}), .b ({new_AGEMA_signal_946, new_AGEMA_signal_944, new_AGEMA_signal_942, new_AGEMA_signal_940}), .c ({new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, M17}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M18_U1 ( .a ({new_AGEMA_signal_285, new_AGEMA_signal_284, new_AGEMA_signal_283, M8}), .b ({new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, M7}), .c ({new_AGEMA_signal_309, new_AGEMA_signal_308, new_AGEMA_signal_307, M18}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M19_U1 ( .a ({new_AGEMA_signal_297, new_AGEMA_signal_296, new_AGEMA_signal_295, M10}), .b ({new_AGEMA_signal_300, new_AGEMA_signal_299, new_AGEMA_signal_298, M15}), .c ({new_AGEMA_signal_312, new_AGEMA_signal_311, new_AGEMA_signal_310, M19}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M20_U1 ( .a ({new_AGEMA_signal_303, new_AGEMA_signal_302, new_AGEMA_signal_301, M16}), .b ({new_AGEMA_signal_291, new_AGEMA_signal_290, new_AGEMA_signal_289, M13}), .c ({new_AGEMA_signal_315, new_AGEMA_signal_314, new_AGEMA_signal_313, M20}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M21_U1 ( .a ({new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, M17}), .b ({new_AGEMA_signal_300, new_AGEMA_signal_299, new_AGEMA_signal_298, M15}), .c ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, M21}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M22_U1 ( .a ({new_AGEMA_signal_309, new_AGEMA_signal_308, new_AGEMA_signal_307, M18}), .b ({new_AGEMA_signal_291, new_AGEMA_signal_290, new_AGEMA_signal_289, M13}), .c ({new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M22}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M23_U1 ( .a ({new_AGEMA_signal_312, new_AGEMA_signal_311, new_AGEMA_signal_310, M19}), .b ({new_AGEMA_signal_954, new_AGEMA_signal_952, new_AGEMA_signal_950, new_AGEMA_signal_948}), .c ({new_AGEMA_signal_324, new_AGEMA_signal_323, new_AGEMA_signal_322, M23}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M24_U1 ( .a ({new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M22}), .b ({new_AGEMA_signal_324, new_AGEMA_signal_323, new_AGEMA_signal_322, M23}), .c ({new_AGEMA_signal_336, new_AGEMA_signal_335, new_AGEMA_signal_334, M24}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M27_U1 ( .a ({new_AGEMA_signal_315, new_AGEMA_signal_314, new_AGEMA_signal_313, M20}), .b ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, M21}), .c ({new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, M27}) ) ;
    buf_clk new_AGEMA_reg_buffer_137 ( .C (clk), .D (new_AGEMA_signal_923), .Q (new_AGEMA_signal_924) ) ;
    buf_clk new_AGEMA_reg_buffer_139 ( .C (clk), .D (new_AGEMA_signal_925), .Q (new_AGEMA_signal_926) ) ;
    buf_clk new_AGEMA_reg_buffer_141 ( .C (clk), .D (new_AGEMA_signal_927), .Q (new_AGEMA_signal_928) ) ;
    buf_clk new_AGEMA_reg_buffer_143 ( .C (clk), .D (new_AGEMA_signal_929), .Q (new_AGEMA_signal_930) ) ;
    buf_clk new_AGEMA_reg_buffer_145 ( .C (clk), .D (new_AGEMA_signal_931), .Q (new_AGEMA_signal_932) ) ;
    buf_clk new_AGEMA_reg_buffer_147 ( .C (clk), .D (new_AGEMA_signal_933), .Q (new_AGEMA_signal_934) ) ;
    buf_clk new_AGEMA_reg_buffer_149 ( .C (clk), .D (new_AGEMA_signal_935), .Q (new_AGEMA_signal_936) ) ;
    buf_clk new_AGEMA_reg_buffer_151 ( .C (clk), .D (new_AGEMA_signal_937), .Q (new_AGEMA_signal_938) ) ;
    buf_clk new_AGEMA_reg_buffer_153 ( .C (clk), .D (new_AGEMA_signal_939), .Q (new_AGEMA_signal_940) ) ;
    buf_clk new_AGEMA_reg_buffer_155 ( .C (clk), .D (new_AGEMA_signal_941), .Q (new_AGEMA_signal_942) ) ;
    buf_clk new_AGEMA_reg_buffer_157 ( .C (clk), .D (new_AGEMA_signal_943), .Q (new_AGEMA_signal_944) ) ;
    buf_clk new_AGEMA_reg_buffer_159 ( .C (clk), .D (new_AGEMA_signal_945), .Q (new_AGEMA_signal_946) ) ;
    buf_clk new_AGEMA_reg_buffer_161 ( .C (clk), .D (new_AGEMA_signal_947), .Q (new_AGEMA_signal_948) ) ;
    buf_clk new_AGEMA_reg_buffer_163 ( .C (clk), .D (new_AGEMA_signal_949), .Q (new_AGEMA_signal_950) ) ;
    buf_clk new_AGEMA_reg_buffer_165 ( .C (clk), .D (new_AGEMA_signal_951), .Q (new_AGEMA_signal_952) ) ;
    buf_clk new_AGEMA_reg_buffer_167 ( .C (clk), .D (new_AGEMA_signal_953), .Q (new_AGEMA_signal_954) ) ;
    buf_clk new_AGEMA_reg_buffer_233 ( .C (clk), .D (new_AGEMA_signal_1019), .Q (new_AGEMA_signal_1020) ) ;
    buf_clk new_AGEMA_reg_buffer_239 ( .C (clk), .D (new_AGEMA_signal_1025), .Q (new_AGEMA_signal_1026) ) ;
    buf_clk new_AGEMA_reg_buffer_245 ( .C (clk), .D (new_AGEMA_signal_1031), .Q (new_AGEMA_signal_1032) ) ;
    buf_clk new_AGEMA_reg_buffer_251 ( .C (clk), .D (new_AGEMA_signal_1037), .Q (new_AGEMA_signal_1038) ) ;
    buf_clk new_AGEMA_reg_buffer_257 ( .C (clk), .D (new_AGEMA_signal_1043), .Q (new_AGEMA_signal_1044) ) ;
    buf_clk new_AGEMA_reg_buffer_263 ( .C (clk), .D (new_AGEMA_signal_1049), .Q (new_AGEMA_signal_1050) ) ;
    buf_clk new_AGEMA_reg_buffer_269 ( .C (clk), .D (new_AGEMA_signal_1055), .Q (new_AGEMA_signal_1056) ) ;
    buf_clk new_AGEMA_reg_buffer_275 ( .C (clk), .D (new_AGEMA_signal_1061), .Q (new_AGEMA_signal_1062) ) ;
    buf_clk new_AGEMA_reg_buffer_281 ( .C (clk), .D (new_AGEMA_signal_1067), .Q (new_AGEMA_signal_1068) ) ;
    buf_clk new_AGEMA_reg_buffer_287 ( .C (clk), .D (new_AGEMA_signal_1073), .Q (new_AGEMA_signal_1074) ) ;
    buf_clk new_AGEMA_reg_buffer_293 ( .C (clk), .D (new_AGEMA_signal_1079), .Q (new_AGEMA_signal_1080) ) ;
    buf_clk new_AGEMA_reg_buffer_299 ( .C (clk), .D (new_AGEMA_signal_1085), .Q (new_AGEMA_signal_1086) ) ;
    buf_clk new_AGEMA_reg_buffer_305 ( .C (clk), .D (new_AGEMA_signal_1091), .Q (new_AGEMA_signal_1092) ) ;
    buf_clk new_AGEMA_reg_buffer_311 ( .C (clk), .D (new_AGEMA_signal_1097), .Q (new_AGEMA_signal_1098) ) ;
    buf_clk new_AGEMA_reg_buffer_317 ( .C (clk), .D (new_AGEMA_signal_1103), .Q (new_AGEMA_signal_1104) ) ;
    buf_clk new_AGEMA_reg_buffer_323 ( .C (clk), .D (new_AGEMA_signal_1109), .Q (new_AGEMA_signal_1110) ) ;
    buf_clk new_AGEMA_reg_buffer_329 ( .C (clk), .D (new_AGEMA_signal_1115), .Q (new_AGEMA_signal_1116) ) ;
    buf_clk new_AGEMA_reg_buffer_335 ( .C (clk), .D (new_AGEMA_signal_1121), .Q (new_AGEMA_signal_1122) ) ;
    buf_clk new_AGEMA_reg_buffer_341 ( .C (clk), .D (new_AGEMA_signal_1127), .Q (new_AGEMA_signal_1128) ) ;
    buf_clk new_AGEMA_reg_buffer_347 ( .C (clk), .D (new_AGEMA_signal_1133), .Q (new_AGEMA_signal_1134) ) ;
    buf_clk new_AGEMA_reg_buffer_353 ( .C (clk), .D (new_AGEMA_signal_1139), .Q (new_AGEMA_signal_1140) ) ;
    buf_clk new_AGEMA_reg_buffer_359 ( .C (clk), .D (new_AGEMA_signal_1145), .Q (new_AGEMA_signal_1146) ) ;
    buf_clk new_AGEMA_reg_buffer_365 ( .C (clk), .D (new_AGEMA_signal_1151), .Q (new_AGEMA_signal_1152) ) ;
    buf_clk new_AGEMA_reg_buffer_371 ( .C (clk), .D (new_AGEMA_signal_1157), .Q (new_AGEMA_signal_1158) ) ;
    buf_clk new_AGEMA_reg_buffer_377 ( .C (clk), .D (new_AGEMA_signal_1163), .Q (new_AGEMA_signal_1164) ) ;
    buf_clk new_AGEMA_reg_buffer_383 ( .C (clk), .D (new_AGEMA_signal_1169), .Q (new_AGEMA_signal_1170) ) ;
    buf_clk new_AGEMA_reg_buffer_389 ( .C (clk), .D (new_AGEMA_signal_1175), .Q (new_AGEMA_signal_1176) ) ;
    buf_clk new_AGEMA_reg_buffer_395 ( .C (clk), .D (new_AGEMA_signal_1181), .Q (new_AGEMA_signal_1182) ) ;
    buf_clk new_AGEMA_reg_buffer_401 ( .C (clk), .D (new_AGEMA_signal_1187), .Q (new_AGEMA_signal_1188) ) ;
    buf_clk new_AGEMA_reg_buffer_407 ( .C (clk), .D (new_AGEMA_signal_1193), .Q (new_AGEMA_signal_1194) ) ;
    buf_clk new_AGEMA_reg_buffer_413 ( .C (clk), .D (new_AGEMA_signal_1199), .Q (new_AGEMA_signal_1200) ) ;
    buf_clk new_AGEMA_reg_buffer_419 ( .C (clk), .D (new_AGEMA_signal_1205), .Q (new_AGEMA_signal_1206) ) ;
    buf_clk new_AGEMA_reg_buffer_425 ( .C (clk), .D (new_AGEMA_signal_1211), .Q (new_AGEMA_signal_1212) ) ;
    buf_clk new_AGEMA_reg_buffer_431 ( .C (clk), .D (new_AGEMA_signal_1217), .Q (new_AGEMA_signal_1218) ) ;
    buf_clk new_AGEMA_reg_buffer_437 ( .C (clk), .D (new_AGEMA_signal_1223), .Q (new_AGEMA_signal_1224) ) ;
    buf_clk new_AGEMA_reg_buffer_443 ( .C (clk), .D (new_AGEMA_signal_1229), .Q (new_AGEMA_signal_1230) ) ;
    buf_clk new_AGEMA_reg_buffer_449 ( .C (clk), .D (new_AGEMA_signal_1235), .Q (new_AGEMA_signal_1236) ) ;
    buf_clk new_AGEMA_reg_buffer_455 ( .C (clk), .D (new_AGEMA_signal_1241), .Q (new_AGEMA_signal_1242) ) ;
    buf_clk new_AGEMA_reg_buffer_461 ( .C (clk), .D (new_AGEMA_signal_1247), .Q (new_AGEMA_signal_1248) ) ;
    buf_clk new_AGEMA_reg_buffer_467 ( .C (clk), .D (new_AGEMA_signal_1253), .Q (new_AGEMA_signal_1254) ) ;
    buf_clk new_AGEMA_reg_buffer_473 ( .C (clk), .D (new_AGEMA_signal_1259), .Q (new_AGEMA_signal_1260) ) ;
    buf_clk new_AGEMA_reg_buffer_479 ( .C (clk), .D (new_AGEMA_signal_1265), .Q (new_AGEMA_signal_1266) ) ;
    buf_clk new_AGEMA_reg_buffer_485 ( .C (clk), .D (new_AGEMA_signal_1271), .Q (new_AGEMA_signal_1272) ) ;
    buf_clk new_AGEMA_reg_buffer_491 ( .C (clk), .D (new_AGEMA_signal_1277), .Q (new_AGEMA_signal_1278) ) ;
    buf_clk new_AGEMA_reg_buffer_497 ( .C (clk), .D (new_AGEMA_signal_1283), .Q (new_AGEMA_signal_1284) ) ;
    buf_clk new_AGEMA_reg_buffer_503 ( .C (clk), .D (new_AGEMA_signal_1289), .Q (new_AGEMA_signal_1290) ) ;
    buf_clk new_AGEMA_reg_buffer_509 ( .C (clk), .D (new_AGEMA_signal_1295), .Q (new_AGEMA_signal_1296) ) ;
    buf_clk new_AGEMA_reg_buffer_515 ( .C (clk), .D (new_AGEMA_signal_1301), .Q (new_AGEMA_signal_1302) ) ;
    buf_clk new_AGEMA_reg_buffer_521 ( .C (clk), .D (new_AGEMA_signal_1307), .Q (new_AGEMA_signal_1308) ) ;
    buf_clk new_AGEMA_reg_buffer_527 ( .C (clk), .D (new_AGEMA_signal_1313), .Q (new_AGEMA_signal_1314) ) ;
    buf_clk new_AGEMA_reg_buffer_533 ( .C (clk), .D (new_AGEMA_signal_1319), .Q (new_AGEMA_signal_1320) ) ;
    buf_clk new_AGEMA_reg_buffer_539 ( .C (clk), .D (new_AGEMA_signal_1325), .Q (new_AGEMA_signal_1326) ) ;
    buf_clk new_AGEMA_reg_buffer_545 ( .C (clk), .D (new_AGEMA_signal_1331), .Q (new_AGEMA_signal_1332) ) ;
    buf_clk new_AGEMA_reg_buffer_551 ( .C (clk), .D (new_AGEMA_signal_1337), .Q (new_AGEMA_signal_1338) ) ;
    buf_clk new_AGEMA_reg_buffer_557 ( .C (clk), .D (new_AGEMA_signal_1343), .Q (new_AGEMA_signal_1344) ) ;
    buf_clk new_AGEMA_reg_buffer_563 ( .C (clk), .D (new_AGEMA_signal_1349), .Q (new_AGEMA_signal_1350) ) ;
    buf_clk new_AGEMA_reg_buffer_569 ( .C (clk), .D (new_AGEMA_signal_1355), .Q (new_AGEMA_signal_1356) ) ;
    buf_clk new_AGEMA_reg_buffer_575 ( .C (clk), .D (new_AGEMA_signal_1361), .Q (new_AGEMA_signal_1362) ) ;
    buf_clk new_AGEMA_reg_buffer_581 ( .C (clk), .D (new_AGEMA_signal_1367), .Q (new_AGEMA_signal_1368) ) ;
    buf_clk new_AGEMA_reg_buffer_587 ( .C (clk), .D (new_AGEMA_signal_1373), .Q (new_AGEMA_signal_1374) ) ;
    buf_clk new_AGEMA_reg_buffer_593 ( .C (clk), .D (new_AGEMA_signal_1379), .Q (new_AGEMA_signal_1380) ) ;
    buf_clk new_AGEMA_reg_buffer_599 ( .C (clk), .D (new_AGEMA_signal_1385), .Q (new_AGEMA_signal_1386) ) ;
    buf_clk new_AGEMA_reg_buffer_605 ( .C (clk), .D (new_AGEMA_signal_1391), .Q (new_AGEMA_signal_1392) ) ;
    buf_clk new_AGEMA_reg_buffer_611 ( .C (clk), .D (new_AGEMA_signal_1397), .Q (new_AGEMA_signal_1398) ) ;
    buf_clk new_AGEMA_reg_buffer_617 ( .C (clk), .D (new_AGEMA_signal_1403), .Q (new_AGEMA_signal_1404) ) ;
    buf_clk new_AGEMA_reg_buffer_623 ( .C (clk), .D (new_AGEMA_signal_1409), .Q (new_AGEMA_signal_1410) ) ;
    buf_clk new_AGEMA_reg_buffer_629 ( .C (clk), .D (new_AGEMA_signal_1415), .Q (new_AGEMA_signal_1416) ) ;
    buf_clk new_AGEMA_reg_buffer_635 ( .C (clk), .D (new_AGEMA_signal_1421), .Q (new_AGEMA_signal_1422) ) ;
    buf_clk new_AGEMA_reg_buffer_641 ( .C (clk), .D (new_AGEMA_signal_1427), .Q (new_AGEMA_signal_1428) ) ;
    buf_clk new_AGEMA_reg_buffer_647 ( .C (clk), .D (new_AGEMA_signal_1433), .Q (new_AGEMA_signal_1434) ) ;
    buf_clk new_AGEMA_reg_buffer_653 ( .C (clk), .D (new_AGEMA_signal_1439), .Q (new_AGEMA_signal_1440) ) ;
    buf_clk new_AGEMA_reg_buffer_659 ( .C (clk), .D (new_AGEMA_signal_1445), .Q (new_AGEMA_signal_1446) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_168 ( .C (clk), .D (M21), .Q (new_AGEMA_signal_955) ) ;
    buf_clk new_AGEMA_reg_buffer_170 ( .C (clk), .D (new_AGEMA_signal_316), .Q (new_AGEMA_signal_957) ) ;
    buf_clk new_AGEMA_reg_buffer_172 ( .C (clk), .D (new_AGEMA_signal_317), .Q (new_AGEMA_signal_959) ) ;
    buf_clk new_AGEMA_reg_buffer_174 ( .C (clk), .D (new_AGEMA_signal_318), .Q (new_AGEMA_signal_961) ) ;
    buf_clk new_AGEMA_reg_buffer_176 ( .C (clk), .D (M23), .Q (new_AGEMA_signal_963) ) ;
    buf_clk new_AGEMA_reg_buffer_178 ( .C (clk), .D (new_AGEMA_signal_322), .Q (new_AGEMA_signal_965) ) ;
    buf_clk new_AGEMA_reg_buffer_180 ( .C (clk), .D (new_AGEMA_signal_323), .Q (new_AGEMA_signal_967) ) ;
    buf_clk new_AGEMA_reg_buffer_182 ( .C (clk), .D (new_AGEMA_signal_324), .Q (new_AGEMA_signal_969) ) ;
    buf_clk new_AGEMA_reg_buffer_184 ( .C (clk), .D (M27), .Q (new_AGEMA_signal_971) ) ;
    buf_clk new_AGEMA_reg_buffer_186 ( .C (clk), .D (new_AGEMA_signal_328), .Q (new_AGEMA_signal_973) ) ;
    buf_clk new_AGEMA_reg_buffer_188 ( .C (clk), .D (new_AGEMA_signal_329), .Q (new_AGEMA_signal_975) ) ;
    buf_clk new_AGEMA_reg_buffer_190 ( .C (clk), .D (new_AGEMA_signal_330), .Q (new_AGEMA_signal_977) ) ;
    buf_clk new_AGEMA_reg_buffer_192 ( .C (clk), .D (M24), .Q (new_AGEMA_signal_979) ) ;
    buf_clk new_AGEMA_reg_buffer_194 ( .C (clk), .D (new_AGEMA_signal_334), .Q (new_AGEMA_signal_981) ) ;
    buf_clk new_AGEMA_reg_buffer_196 ( .C (clk), .D (new_AGEMA_signal_335), .Q (new_AGEMA_signal_983) ) ;
    buf_clk new_AGEMA_reg_buffer_198 ( .C (clk), .D (new_AGEMA_signal_336), .Q (new_AGEMA_signal_985) ) ;
    buf_clk new_AGEMA_reg_buffer_234 ( .C (clk), .D (new_AGEMA_signal_1020), .Q (new_AGEMA_signal_1021) ) ;
    buf_clk new_AGEMA_reg_buffer_240 ( .C (clk), .D (new_AGEMA_signal_1026), .Q (new_AGEMA_signal_1027) ) ;
    buf_clk new_AGEMA_reg_buffer_246 ( .C (clk), .D (new_AGEMA_signal_1032), .Q (new_AGEMA_signal_1033) ) ;
    buf_clk new_AGEMA_reg_buffer_252 ( .C (clk), .D (new_AGEMA_signal_1038), .Q (new_AGEMA_signal_1039) ) ;
    buf_clk new_AGEMA_reg_buffer_258 ( .C (clk), .D (new_AGEMA_signal_1044), .Q (new_AGEMA_signal_1045) ) ;
    buf_clk new_AGEMA_reg_buffer_264 ( .C (clk), .D (new_AGEMA_signal_1050), .Q (new_AGEMA_signal_1051) ) ;
    buf_clk new_AGEMA_reg_buffer_270 ( .C (clk), .D (new_AGEMA_signal_1056), .Q (new_AGEMA_signal_1057) ) ;
    buf_clk new_AGEMA_reg_buffer_276 ( .C (clk), .D (new_AGEMA_signal_1062), .Q (new_AGEMA_signal_1063) ) ;
    buf_clk new_AGEMA_reg_buffer_282 ( .C (clk), .D (new_AGEMA_signal_1068), .Q (new_AGEMA_signal_1069) ) ;
    buf_clk new_AGEMA_reg_buffer_288 ( .C (clk), .D (new_AGEMA_signal_1074), .Q (new_AGEMA_signal_1075) ) ;
    buf_clk new_AGEMA_reg_buffer_294 ( .C (clk), .D (new_AGEMA_signal_1080), .Q (new_AGEMA_signal_1081) ) ;
    buf_clk new_AGEMA_reg_buffer_300 ( .C (clk), .D (new_AGEMA_signal_1086), .Q (new_AGEMA_signal_1087) ) ;
    buf_clk new_AGEMA_reg_buffer_306 ( .C (clk), .D (new_AGEMA_signal_1092), .Q (new_AGEMA_signal_1093) ) ;
    buf_clk new_AGEMA_reg_buffer_312 ( .C (clk), .D (new_AGEMA_signal_1098), .Q (new_AGEMA_signal_1099) ) ;
    buf_clk new_AGEMA_reg_buffer_318 ( .C (clk), .D (new_AGEMA_signal_1104), .Q (new_AGEMA_signal_1105) ) ;
    buf_clk new_AGEMA_reg_buffer_324 ( .C (clk), .D (new_AGEMA_signal_1110), .Q (new_AGEMA_signal_1111) ) ;
    buf_clk new_AGEMA_reg_buffer_330 ( .C (clk), .D (new_AGEMA_signal_1116), .Q (new_AGEMA_signal_1117) ) ;
    buf_clk new_AGEMA_reg_buffer_336 ( .C (clk), .D (new_AGEMA_signal_1122), .Q (new_AGEMA_signal_1123) ) ;
    buf_clk new_AGEMA_reg_buffer_342 ( .C (clk), .D (new_AGEMA_signal_1128), .Q (new_AGEMA_signal_1129) ) ;
    buf_clk new_AGEMA_reg_buffer_348 ( .C (clk), .D (new_AGEMA_signal_1134), .Q (new_AGEMA_signal_1135) ) ;
    buf_clk new_AGEMA_reg_buffer_354 ( .C (clk), .D (new_AGEMA_signal_1140), .Q (new_AGEMA_signal_1141) ) ;
    buf_clk new_AGEMA_reg_buffer_360 ( .C (clk), .D (new_AGEMA_signal_1146), .Q (new_AGEMA_signal_1147) ) ;
    buf_clk new_AGEMA_reg_buffer_366 ( .C (clk), .D (new_AGEMA_signal_1152), .Q (new_AGEMA_signal_1153) ) ;
    buf_clk new_AGEMA_reg_buffer_372 ( .C (clk), .D (new_AGEMA_signal_1158), .Q (new_AGEMA_signal_1159) ) ;
    buf_clk new_AGEMA_reg_buffer_378 ( .C (clk), .D (new_AGEMA_signal_1164), .Q (new_AGEMA_signal_1165) ) ;
    buf_clk new_AGEMA_reg_buffer_384 ( .C (clk), .D (new_AGEMA_signal_1170), .Q (new_AGEMA_signal_1171) ) ;
    buf_clk new_AGEMA_reg_buffer_390 ( .C (clk), .D (new_AGEMA_signal_1176), .Q (new_AGEMA_signal_1177) ) ;
    buf_clk new_AGEMA_reg_buffer_396 ( .C (clk), .D (new_AGEMA_signal_1182), .Q (new_AGEMA_signal_1183) ) ;
    buf_clk new_AGEMA_reg_buffer_402 ( .C (clk), .D (new_AGEMA_signal_1188), .Q (new_AGEMA_signal_1189) ) ;
    buf_clk new_AGEMA_reg_buffer_408 ( .C (clk), .D (new_AGEMA_signal_1194), .Q (new_AGEMA_signal_1195) ) ;
    buf_clk new_AGEMA_reg_buffer_414 ( .C (clk), .D (new_AGEMA_signal_1200), .Q (new_AGEMA_signal_1201) ) ;
    buf_clk new_AGEMA_reg_buffer_420 ( .C (clk), .D (new_AGEMA_signal_1206), .Q (new_AGEMA_signal_1207) ) ;
    buf_clk new_AGEMA_reg_buffer_426 ( .C (clk), .D (new_AGEMA_signal_1212), .Q (new_AGEMA_signal_1213) ) ;
    buf_clk new_AGEMA_reg_buffer_432 ( .C (clk), .D (new_AGEMA_signal_1218), .Q (new_AGEMA_signal_1219) ) ;
    buf_clk new_AGEMA_reg_buffer_438 ( .C (clk), .D (new_AGEMA_signal_1224), .Q (new_AGEMA_signal_1225) ) ;
    buf_clk new_AGEMA_reg_buffer_444 ( .C (clk), .D (new_AGEMA_signal_1230), .Q (new_AGEMA_signal_1231) ) ;
    buf_clk new_AGEMA_reg_buffer_450 ( .C (clk), .D (new_AGEMA_signal_1236), .Q (new_AGEMA_signal_1237) ) ;
    buf_clk new_AGEMA_reg_buffer_456 ( .C (clk), .D (new_AGEMA_signal_1242), .Q (new_AGEMA_signal_1243) ) ;
    buf_clk new_AGEMA_reg_buffer_462 ( .C (clk), .D (new_AGEMA_signal_1248), .Q (new_AGEMA_signal_1249) ) ;
    buf_clk new_AGEMA_reg_buffer_468 ( .C (clk), .D (new_AGEMA_signal_1254), .Q (new_AGEMA_signal_1255) ) ;
    buf_clk new_AGEMA_reg_buffer_474 ( .C (clk), .D (new_AGEMA_signal_1260), .Q (new_AGEMA_signal_1261) ) ;
    buf_clk new_AGEMA_reg_buffer_480 ( .C (clk), .D (new_AGEMA_signal_1266), .Q (new_AGEMA_signal_1267) ) ;
    buf_clk new_AGEMA_reg_buffer_486 ( .C (clk), .D (new_AGEMA_signal_1272), .Q (new_AGEMA_signal_1273) ) ;
    buf_clk new_AGEMA_reg_buffer_492 ( .C (clk), .D (new_AGEMA_signal_1278), .Q (new_AGEMA_signal_1279) ) ;
    buf_clk new_AGEMA_reg_buffer_498 ( .C (clk), .D (new_AGEMA_signal_1284), .Q (new_AGEMA_signal_1285) ) ;
    buf_clk new_AGEMA_reg_buffer_504 ( .C (clk), .D (new_AGEMA_signal_1290), .Q (new_AGEMA_signal_1291) ) ;
    buf_clk new_AGEMA_reg_buffer_510 ( .C (clk), .D (new_AGEMA_signal_1296), .Q (new_AGEMA_signal_1297) ) ;
    buf_clk new_AGEMA_reg_buffer_516 ( .C (clk), .D (new_AGEMA_signal_1302), .Q (new_AGEMA_signal_1303) ) ;
    buf_clk new_AGEMA_reg_buffer_522 ( .C (clk), .D (new_AGEMA_signal_1308), .Q (new_AGEMA_signal_1309) ) ;
    buf_clk new_AGEMA_reg_buffer_528 ( .C (clk), .D (new_AGEMA_signal_1314), .Q (new_AGEMA_signal_1315) ) ;
    buf_clk new_AGEMA_reg_buffer_534 ( .C (clk), .D (new_AGEMA_signal_1320), .Q (new_AGEMA_signal_1321) ) ;
    buf_clk new_AGEMA_reg_buffer_540 ( .C (clk), .D (new_AGEMA_signal_1326), .Q (new_AGEMA_signal_1327) ) ;
    buf_clk new_AGEMA_reg_buffer_546 ( .C (clk), .D (new_AGEMA_signal_1332), .Q (new_AGEMA_signal_1333) ) ;
    buf_clk new_AGEMA_reg_buffer_552 ( .C (clk), .D (new_AGEMA_signal_1338), .Q (new_AGEMA_signal_1339) ) ;
    buf_clk new_AGEMA_reg_buffer_558 ( .C (clk), .D (new_AGEMA_signal_1344), .Q (new_AGEMA_signal_1345) ) ;
    buf_clk new_AGEMA_reg_buffer_564 ( .C (clk), .D (new_AGEMA_signal_1350), .Q (new_AGEMA_signal_1351) ) ;
    buf_clk new_AGEMA_reg_buffer_570 ( .C (clk), .D (new_AGEMA_signal_1356), .Q (new_AGEMA_signal_1357) ) ;
    buf_clk new_AGEMA_reg_buffer_576 ( .C (clk), .D (new_AGEMA_signal_1362), .Q (new_AGEMA_signal_1363) ) ;
    buf_clk new_AGEMA_reg_buffer_582 ( .C (clk), .D (new_AGEMA_signal_1368), .Q (new_AGEMA_signal_1369) ) ;
    buf_clk new_AGEMA_reg_buffer_588 ( .C (clk), .D (new_AGEMA_signal_1374), .Q (new_AGEMA_signal_1375) ) ;
    buf_clk new_AGEMA_reg_buffer_594 ( .C (clk), .D (new_AGEMA_signal_1380), .Q (new_AGEMA_signal_1381) ) ;
    buf_clk new_AGEMA_reg_buffer_600 ( .C (clk), .D (new_AGEMA_signal_1386), .Q (new_AGEMA_signal_1387) ) ;
    buf_clk new_AGEMA_reg_buffer_606 ( .C (clk), .D (new_AGEMA_signal_1392), .Q (new_AGEMA_signal_1393) ) ;
    buf_clk new_AGEMA_reg_buffer_612 ( .C (clk), .D (new_AGEMA_signal_1398), .Q (new_AGEMA_signal_1399) ) ;
    buf_clk new_AGEMA_reg_buffer_618 ( .C (clk), .D (new_AGEMA_signal_1404), .Q (new_AGEMA_signal_1405) ) ;
    buf_clk new_AGEMA_reg_buffer_624 ( .C (clk), .D (new_AGEMA_signal_1410), .Q (new_AGEMA_signal_1411) ) ;
    buf_clk new_AGEMA_reg_buffer_630 ( .C (clk), .D (new_AGEMA_signal_1416), .Q (new_AGEMA_signal_1417) ) ;
    buf_clk new_AGEMA_reg_buffer_636 ( .C (clk), .D (new_AGEMA_signal_1422), .Q (new_AGEMA_signal_1423) ) ;
    buf_clk new_AGEMA_reg_buffer_642 ( .C (clk), .D (new_AGEMA_signal_1428), .Q (new_AGEMA_signal_1429) ) ;
    buf_clk new_AGEMA_reg_buffer_648 ( .C (clk), .D (new_AGEMA_signal_1434), .Q (new_AGEMA_signal_1435) ) ;
    buf_clk new_AGEMA_reg_buffer_654 ( .C (clk), .D (new_AGEMA_signal_1440), .Q (new_AGEMA_signal_1441) ) ;
    buf_clk new_AGEMA_reg_buffer_660 ( .C (clk), .D (new_AGEMA_signal_1446), .Q (new_AGEMA_signal_1447) ) ;

    /* cells in depth 4 */
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M25_U1 ( .ina ({new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M22}), .inb ({new_AGEMA_signal_315, new_AGEMA_signal_314, new_AGEMA_signal_313, M20}), .clk (clk), .rnd ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .outt ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, M25}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M26_U1 ( .a ({new_AGEMA_signal_962, new_AGEMA_signal_960, new_AGEMA_signal_958, new_AGEMA_signal_956}), .b ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, M25}), .c ({new_AGEMA_signal_339, new_AGEMA_signal_338, new_AGEMA_signal_337, M26}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M28_U1 ( .a ({new_AGEMA_signal_970, new_AGEMA_signal_968, new_AGEMA_signal_966, new_AGEMA_signal_964}), .b ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, M25}), .c ({new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, M28}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M31_U1 ( .ina ({new_AGEMA_signal_315, new_AGEMA_signal_314, new_AGEMA_signal_313, M20}), .inb ({new_AGEMA_signal_324, new_AGEMA_signal_323, new_AGEMA_signal_322, M23}), .clk (clk), .rnd ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .outt ({new_AGEMA_signal_345, new_AGEMA_signal_344, new_AGEMA_signal_343, M31}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M33_U1 ( .a ({new_AGEMA_signal_978, new_AGEMA_signal_976, new_AGEMA_signal_974, new_AGEMA_signal_972}), .b ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, M25}), .c ({new_AGEMA_signal_348, new_AGEMA_signal_347, new_AGEMA_signal_346, M33}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M34_U1 ( .ina ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, M21}), .inb ({new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M22}), .clk (clk), .rnd ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .outt ({new_AGEMA_signal_333, new_AGEMA_signal_332, new_AGEMA_signal_331, M34}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M36_U1 ( .a ({new_AGEMA_signal_986, new_AGEMA_signal_984, new_AGEMA_signal_982, new_AGEMA_signal_980}), .b ({new_AGEMA_signal_327, new_AGEMA_signal_326, new_AGEMA_signal_325, M25}), .c ({new_AGEMA_signal_363, new_AGEMA_signal_362, new_AGEMA_signal_361, M36}) ) ;
    buf_clk new_AGEMA_reg_buffer_169 ( .C (clk), .D (new_AGEMA_signal_955), .Q (new_AGEMA_signal_956) ) ;
    buf_clk new_AGEMA_reg_buffer_171 ( .C (clk), .D (new_AGEMA_signal_957), .Q (new_AGEMA_signal_958) ) ;
    buf_clk new_AGEMA_reg_buffer_173 ( .C (clk), .D (new_AGEMA_signal_959), .Q (new_AGEMA_signal_960) ) ;
    buf_clk new_AGEMA_reg_buffer_175 ( .C (clk), .D (new_AGEMA_signal_961), .Q (new_AGEMA_signal_962) ) ;
    buf_clk new_AGEMA_reg_buffer_177 ( .C (clk), .D (new_AGEMA_signal_963), .Q (new_AGEMA_signal_964) ) ;
    buf_clk new_AGEMA_reg_buffer_179 ( .C (clk), .D (new_AGEMA_signal_965), .Q (new_AGEMA_signal_966) ) ;
    buf_clk new_AGEMA_reg_buffer_181 ( .C (clk), .D (new_AGEMA_signal_967), .Q (new_AGEMA_signal_968) ) ;
    buf_clk new_AGEMA_reg_buffer_183 ( .C (clk), .D (new_AGEMA_signal_969), .Q (new_AGEMA_signal_970) ) ;
    buf_clk new_AGEMA_reg_buffer_185 ( .C (clk), .D (new_AGEMA_signal_971), .Q (new_AGEMA_signal_972) ) ;
    buf_clk new_AGEMA_reg_buffer_187 ( .C (clk), .D (new_AGEMA_signal_973), .Q (new_AGEMA_signal_974) ) ;
    buf_clk new_AGEMA_reg_buffer_189 ( .C (clk), .D (new_AGEMA_signal_975), .Q (new_AGEMA_signal_976) ) ;
    buf_clk new_AGEMA_reg_buffer_191 ( .C (clk), .D (new_AGEMA_signal_977), .Q (new_AGEMA_signal_978) ) ;
    buf_clk new_AGEMA_reg_buffer_193 ( .C (clk), .D (new_AGEMA_signal_979), .Q (new_AGEMA_signal_980) ) ;
    buf_clk new_AGEMA_reg_buffer_195 ( .C (clk), .D (new_AGEMA_signal_981), .Q (new_AGEMA_signal_982) ) ;
    buf_clk new_AGEMA_reg_buffer_197 ( .C (clk), .D (new_AGEMA_signal_983), .Q (new_AGEMA_signal_984) ) ;
    buf_clk new_AGEMA_reg_buffer_199 ( .C (clk), .D (new_AGEMA_signal_985), .Q (new_AGEMA_signal_986) ) ;
    buf_clk new_AGEMA_reg_buffer_235 ( .C (clk), .D (new_AGEMA_signal_1021), .Q (new_AGEMA_signal_1022) ) ;
    buf_clk new_AGEMA_reg_buffer_241 ( .C (clk), .D (new_AGEMA_signal_1027), .Q (new_AGEMA_signal_1028) ) ;
    buf_clk new_AGEMA_reg_buffer_247 ( .C (clk), .D (new_AGEMA_signal_1033), .Q (new_AGEMA_signal_1034) ) ;
    buf_clk new_AGEMA_reg_buffer_253 ( .C (clk), .D (new_AGEMA_signal_1039), .Q (new_AGEMA_signal_1040) ) ;
    buf_clk new_AGEMA_reg_buffer_259 ( .C (clk), .D (new_AGEMA_signal_1045), .Q (new_AGEMA_signal_1046) ) ;
    buf_clk new_AGEMA_reg_buffer_265 ( .C (clk), .D (new_AGEMA_signal_1051), .Q (new_AGEMA_signal_1052) ) ;
    buf_clk new_AGEMA_reg_buffer_271 ( .C (clk), .D (new_AGEMA_signal_1057), .Q (new_AGEMA_signal_1058) ) ;
    buf_clk new_AGEMA_reg_buffer_277 ( .C (clk), .D (new_AGEMA_signal_1063), .Q (new_AGEMA_signal_1064) ) ;
    buf_clk new_AGEMA_reg_buffer_283 ( .C (clk), .D (new_AGEMA_signal_1069), .Q (new_AGEMA_signal_1070) ) ;
    buf_clk new_AGEMA_reg_buffer_289 ( .C (clk), .D (new_AGEMA_signal_1075), .Q (new_AGEMA_signal_1076) ) ;
    buf_clk new_AGEMA_reg_buffer_295 ( .C (clk), .D (new_AGEMA_signal_1081), .Q (new_AGEMA_signal_1082) ) ;
    buf_clk new_AGEMA_reg_buffer_301 ( .C (clk), .D (new_AGEMA_signal_1087), .Q (new_AGEMA_signal_1088) ) ;
    buf_clk new_AGEMA_reg_buffer_307 ( .C (clk), .D (new_AGEMA_signal_1093), .Q (new_AGEMA_signal_1094) ) ;
    buf_clk new_AGEMA_reg_buffer_313 ( .C (clk), .D (new_AGEMA_signal_1099), .Q (new_AGEMA_signal_1100) ) ;
    buf_clk new_AGEMA_reg_buffer_319 ( .C (clk), .D (new_AGEMA_signal_1105), .Q (new_AGEMA_signal_1106) ) ;
    buf_clk new_AGEMA_reg_buffer_325 ( .C (clk), .D (new_AGEMA_signal_1111), .Q (new_AGEMA_signal_1112) ) ;
    buf_clk new_AGEMA_reg_buffer_331 ( .C (clk), .D (new_AGEMA_signal_1117), .Q (new_AGEMA_signal_1118) ) ;
    buf_clk new_AGEMA_reg_buffer_337 ( .C (clk), .D (new_AGEMA_signal_1123), .Q (new_AGEMA_signal_1124) ) ;
    buf_clk new_AGEMA_reg_buffer_343 ( .C (clk), .D (new_AGEMA_signal_1129), .Q (new_AGEMA_signal_1130) ) ;
    buf_clk new_AGEMA_reg_buffer_349 ( .C (clk), .D (new_AGEMA_signal_1135), .Q (new_AGEMA_signal_1136) ) ;
    buf_clk new_AGEMA_reg_buffer_355 ( .C (clk), .D (new_AGEMA_signal_1141), .Q (new_AGEMA_signal_1142) ) ;
    buf_clk new_AGEMA_reg_buffer_361 ( .C (clk), .D (new_AGEMA_signal_1147), .Q (new_AGEMA_signal_1148) ) ;
    buf_clk new_AGEMA_reg_buffer_367 ( .C (clk), .D (new_AGEMA_signal_1153), .Q (new_AGEMA_signal_1154) ) ;
    buf_clk new_AGEMA_reg_buffer_373 ( .C (clk), .D (new_AGEMA_signal_1159), .Q (new_AGEMA_signal_1160) ) ;
    buf_clk new_AGEMA_reg_buffer_379 ( .C (clk), .D (new_AGEMA_signal_1165), .Q (new_AGEMA_signal_1166) ) ;
    buf_clk new_AGEMA_reg_buffer_385 ( .C (clk), .D (new_AGEMA_signal_1171), .Q (new_AGEMA_signal_1172) ) ;
    buf_clk new_AGEMA_reg_buffer_391 ( .C (clk), .D (new_AGEMA_signal_1177), .Q (new_AGEMA_signal_1178) ) ;
    buf_clk new_AGEMA_reg_buffer_397 ( .C (clk), .D (new_AGEMA_signal_1183), .Q (new_AGEMA_signal_1184) ) ;
    buf_clk new_AGEMA_reg_buffer_403 ( .C (clk), .D (new_AGEMA_signal_1189), .Q (new_AGEMA_signal_1190) ) ;
    buf_clk new_AGEMA_reg_buffer_409 ( .C (clk), .D (new_AGEMA_signal_1195), .Q (new_AGEMA_signal_1196) ) ;
    buf_clk new_AGEMA_reg_buffer_415 ( .C (clk), .D (new_AGEMA_signal_1201), .Q (new_AGEMA_signal_1202) ) ;
    buf_clk new_AGEMA_reg_buffer_421 ( .C (clk), .D (new_AGEMA_signal_1207), .Q (new_AGEMA_signal_1208) ) ;
    buf_clk new_AGEMA_reg_buffer_427 ( .C (clk), .D (new_AGEMA_signal_1213), .Q (new_AGEMA_signal_1214) ) ;
    buf_clk new_AGEMA_reg_buffer_433 ( .C (clk), .D (new_AGEMA_signal_1219), .Q (new_AGEMA_signal_1220) ) ;
    buf_clk new_AGEMA_reg_buffer_439 ( .C (clk), .D (new_AGEMA_signal_1225), .Q (new_AGEMA_signal_1226) ) ;
    buf_clk new_AGEMA_reg_buffer_445 ( .C (clk), .D (new_AGEMA_signal_1231), .Q (new_AGEMA_signal_1232) ) ;
    buf_clk new_AGEMA_reg_buffer_451 ( .C (clk), .D (new_AGEMA_signal_1237), .Q (new_AGEMA_signal_1238) ) ;
    buf_clk new_AGEMA_reg_buffer_457 ( .C (clk), .D (new_AGEMA_signal_1243), .Q (new_AGEMA_signal_1244) ) ;
    buf_clk new_AGEMA_reg_buffer_463 ( .C (clk), .D (new_AGEMA_signal_1249), .Q (new_AGEMA_signal_1250) ) ;
    buf_clk new_AGEMA_reg_buffer_469 ( .C (clk), .D (new_AGEMA_signal_1255), .Q (new_AGEMA_signal_1256) ) ;
    buf_clk new_AGEMA_reg_buffer_475 ( .C (clk), .D (new_AGEMA_signal_1261), .Q (new_AGEMA_signal_1262) ) ;
    buf_clk new_AGEMA_reg_buffer_481 ( .C (clk), .D (new_AGEMA_signal_1267), .Q (new_AGEMA_signal_1268) ) ;
    buf_clk new_AGEMA_reg_buffer_487 ( .C (clk), .D (new_AGEMA_signal_1273), .Q (new_AGEMA_signal_1274) ) ;
    buf_clk new_AGEMA_reg_buffer_493 ( .C (clk), .D (new_AGEMA_signal_1279), .Q (new_AGEMA_signal_1280) ) ;
    buf_clk new_AGEMA_reg_buffer_499 ( .C (clk), .D (new_AGEMA_signal_1285), .Q (new_AGEMA_signal_1286) ) ;
    buf_clk new_AGEMA_reg_buffer_505 ( .C (clk), .D (new_AGEMA_signal_1291), .Q (new_AGEMA_signal_1292) ) ;
    buf_clk new_AGEMA_reg_buffer_511 ( .C (clk), .D (new_AGEMA_signal_1297), .Q (new_AGEMA_signal_1298) ) ;
    buf_clk new_AGEMA_reg_buffer_517 ( .C (clk), .D (new_AGEMA_signal_1303), .Q (new_AGEMA_signal_1304) ) ;
    buf_clk new_AGEMA_reg_buffer_523 ( .C (clk), .D (new_AGEMA_signal_1309), .Q (new_AGEMA_signal_1310) ) ;
    buf_clk new_AGEMA_reg_buffer_529 ( .C (clk), .D (new_AGEMA_signal_1315), .Q (new_AGEMA_signal_1316) ) ;
    buf_clk new_AGEMA_reg_buffer_535 ( .C (clk), .D (new_AGEMA_signal_1321), .Q (new_AGEMA_signal_1322) ) ;
    buf_clk new_AGEMA_reg_buffer_541 ( .C (clk), .D (new_AGEMA_signal_1327), .Q (new_AGEMA_signal_1328) ) ;
    buf_clk new_AGEMA_reg_buffer_547 ( .C (clk), .D (new_AGEMA_signal_1333), .Q (new_AGEMA_signal_1334) ) ;
    buf_clk new_AGEMA_reg_buffer_553 ( .C (clk), .D (new_AGEMA_signal_1339), .Q (new_AGEMA_signal_1340) ) ;
    buf_clk new_AGEMA_reg_buffer_559 ( .C (clk), .D (new_AGEMA_signal_1345), .Q (new_AGEMA_signal_1346) ) ;
    buf_clk new_AGEMA_reg_buffer_565 ( .C (clk), .D (new_AGEMA_signal_1351), .Q (new_AGEMA_signal_1352) ) ;
    buf_clk new_AGEMA_reg_buffer_571 ( .C (clk), .D (new_AGEMA_signal_1357), .Q (new_AGEMA_signal_1358) ) ;
    buf_clk new_AGEMA_reg_buffer_577 ( .C (clk), .D (new_AGEMA_signal_1363), .Q (new_AGEMA_signal_1364) ) ;
    buf_clk new_AGEMA_reg_buffer_583 ( .C (clk), .D (new_AGEMA_signal_1369), .Q (new_AGEMA_signal_1370) ) ;
    buf_clk new_AGEMA_reg_buffer_589 ( .C (clk), .D (new_AGEMA_signal_1375), .Q (new_AGEMA_signal_1376) ) ;
    buf_clk new_AGEMA_reg_buffer_595 ( .C (clk), .D (new_AGEMA_signal_1381), .Q (new_AGEMA_signal_1382) ) ;
    buf_clk new_AGEMA_reg_buffer_601 ( .C (clk), .D (new_AGEMA_signal_1387), .Q (new_AGEMA_signal_1388) ) ;
    buf_clk new_AGEMA_reg_buffer_607 ( .C (clk), .D (new_AGEMA_signal_1393), .Q (new_AGEMA_signal_1394) ) ;
    buf_clk new_AGEMA_reg_buffer_613 ( .C (clk), .D (new_AGEMA_signal_1399), .Q (new_AGEMA_signal_1400) ) ;
    buf_clk new_AGEMA_reg_buffer_619 ( .C (clk), .D (new_AGEMA_signal_1405), .Q (new_AGEMA_signal_1406) ) ;
    buf_clk new_AGEMA_reg_buffer_625 ( .C (clk), .D (new_AGEMA_signal_1411), .Q (new_AGEMA_signal_1412) ) ;
    buf_clk new_AGEMA_reg_buffer_631 ( .C (clk), .D (new_AGEMA_signal_1417), .Q (new_AGEMA_signal_1418) ) ;
    buf_clk new_AGEMA_reg_buffer_637 ( .C (clk), .D (new_AGEMA_signal_1423), .Q (new_AGEMA_signal_1424) ) ;
    buf_clk new_AGEMA_reg_buffer_643 ( .C (clk), .D (new_AGEMA_signal_1429), .Q (new_AGEMA_signal_1430) ) ;
    buf_clk new_AGEMA_reg_buffer_649 ( .C (clk), .D (new_AGEMA_signal_1435), .Q (new_AGEMA_signal_1436) ) ;
    buf_clk new_AGEMA_reg_buffer_655 ( .C (clk), .D (new_AGEMA_signal_1441), .Q (new_AGEMA_signal_1442) ) ;
    buf_clk new_AGEMA_reg_buffer_661 ( .C (clk), .D (new_AGEMA_signal_1447), .Q (new_AGEMA_signal_1448) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_200 ( .C (clk), .D (new_AGEMA_signal_956), .Q (new_AGEMA_signal_987) ) ;
    buf_clk new_AGEMA_reg_buffer_202 ( .C (clk), .D (new_AGEMA_signal_958), .Q (new_AGEMA_signal_989) ) ;
    buf_clk new_AGEMA_reg_buffer_204 ( .C (clk), .D (new_AGEMA_signal_960), .Q (new_AGEMA_signal_991) ) ;
    buf_clk new_AGEMA_reg_buffer_206 ( .C (clk), .D (new_AGEMA_signal_962), .Q (new_AGEMA_signal_993) ) ;
    buf_clk new_AGEMA_reg_buffer_208 ( .C (clk), .D (M33), .Q (new_AGEMA_signal_995) ) ;
    buf_clk new_AGEMA_reg_buffer_210 ( .C (clk), .D (new_AGEMA_signal_346), .Q (new_AGEMA_signal_997) ) ;
    buf_clk new_AGEMA_reg_buffer_212 ( .C (clk), .D (new_AGEMA_signal_347), .Q (new_AGEMA_signal_999) ) ;
    buf_clk new_AGEMA_reg_buffer_214 ( .C (clk), .D (new_AGEMA_signal_348), .Q (new_AGEMA_signal_1001) ) ;
    buf_clk new_AGEMA_reg_buffer_216 ( .C (clk), .D (new_AGEMA_signal_964), .Q (new_AGEMA_signal_1003) ) ;
    buf_clk new_AGEMA_reg_buffer_218 ( .C (clk), .D (new_AGEMA_signal_966), .Q (new_AGEMA_signal_1005) ) ;
    buf_clk new_AGEMA_reg_buffer_220 ( .C (clk), .D (new_AGEMA_signal_968), .Q (new_AGEMA_signal_1007) ) ;
    buf_clk new_AGEMA_reg_buffer_222 ( .C (clk), .D (new_AGEMA_signal_970), .Q (new_AGEMA_signal_1009) ) ;
    buf_clk new_AGEMA_reg_buffer_224 ( .C (clk), .D (M36), .Q (new_AGEMA_signal_1011) ) ;
    buf_clk new_AGEMA_reg_buffer_226 ( .C (clk), .D (new_AGEMA_signal_361), .Q (new_AGEMA_signal_1013) ) ;
    buf_clk new_AGEMA_reg_buffer_228 ( .C (clk), .D (new_AGEMA_signal_362), .Q (new_AGEMA_signal_1015) ) ;
    buf_clk new_AGEMA_reg_buffer_230 ( .C (clk), .D (new_AGEMA_signal_363), .Q (new_AGEMA_signal_1017) ) ;
    buf_clk new_AGEMA_reg_buffer_236 ( .C (clk), .D (new_AGEMA_signal_1022), .Q (new_AGEMA_signal_1023) ) ;
    buf_clk new_AGEMA_reg_buffer_242 ( .C (clk), .D (new_AGEMA_signal_1028), .Q (new_AGEMA_signal_1029) ) ;
    buf_clk new_AGEMA_reg_buffer_248 ( .C (clk), .D (new_AGEMA_signal_1034), .Q (new_AGEMA_signal_1035) ) ;
    buf_clk new_AGEMA_reg_buffer_254 ( .C (clk), .D (new_AGEMA_signal_1040), .Q (new_AGEMA_signal_1041) ) ;
    buf_clk new_AGEMA_reg_buffer_260 ( .C (clk), .D (new_AGEMA_signal_1046), .Q (new_AGEMA_signal_1047) ) ;
    buf_clk new_AGEMA_reg_buffer_266 ( .C (clk), .D (new_AGEMA_signal_1052), .Q (new_AGEMA_signal_1053) ) ;
    buf_clk new_AGEMA_reg_buffer_272 ( .C (clk), .D (new_AGEMA_signal_1058), .Q (new_AGEMA_signal_1059) ) ;
    buf_clk new_AGEMA_reg_buffer_278 ( .C (clk), .D (new_AGEMA_signal_1064), .Q (new_AGEMA_signal_1065) ) ;
    buf_clk new_AGEMA_reg_buffer_284 ( .C (clk), .D (new_AGEMA_signal_1070), .Q (new_AGEMA_signal_1071) ) ;
    buf_clk new_AGEMA_reg_buffer_290 ( .C (clk), .D (new_AGEMA_signal_1076), .Q (new_AGEMA_signal_1077) ) ;
    buf_clk new_AGEMA_reg_buffer_296 ( .C (clk), .D (new_AGEMA_signal_1082), .Q (new_AGEMA_signal_1083) ) ;
    buf_clk new_AGEMA_reg_buffer_302 ( .C (clk), .D (new_AGEMA_signal_1088), .Q (new_AGEMA_signal_1089) ) ;
    buf_clk new_AGEMA_reg_buffer_308 ( .C (clk), .D (new_AGEMA_signal_1094), .Q (new_AGEMA_signal_1095) ) ;
    buf_clk new_AGEMA_reg_buffer_314 ( .C (clk), .D (new_AGEMA_signal_1100), .Q (new_AGEMA_signal_1101) ) ;
    buf_clk new_AGEMA_reg_buffer_320 ( .C (clk), .D (new_AGEMA_signal_1106), .Q (new_AGEMA_signal_1107) ) ;
    buf_clk new_AGEMA_reg_buffer_326 ( .C (clk), .D (new_AGEMA_signal_1112), .Q (new_AGEMA_signal_1113) ) ;
    buf_clk new_AGEMA_reg_buffer_332 ( .C (clk), .D (new_AGEMA_signal_1118), .Q (new_AGEMA_signal_1119) ) ;
    buf_clk new_AGEMA_reg_buffer_338 ( .C (clk), .D (new_AGEMA_signal_1124), .Q (new_AGEMA_signal_1125) ) ;
    buf_clk new_AGEMA_reg_buffer_344 ( .C (clk), .D (new_AGEMA_signal_1130), .Q (new_AGEMA_signal_1131) ) ;
    buf_clk new_AGEMA_reg_buffer_350 ( .C (clk), .D (new_AGEMA_signal_1136), .Q (new_AGEMA_signal_1137) ) ;
    buf_clk new_AGEMA_reg_buffer_356 ( .C (clk), .D (new_AGEMA_signal_1142), .Q (new_AGEMA_signal_1143) ) ;
    buf_clk new_AGEMA_reg_buffer_362 ( .C (clk), .D (new_AGEMA_signal_1148), .Q (new_AGEMA_signal_1149) ) ;
    buf_clk new_AGEMA_reg_buffer_368 ( .C (clk), .D (new_AGEMA_signal_1154), .Q (new_AGEMA_signal_1155) ) ;
    buf_clk new_AGEMA_reg_buffer_374 ( .C (clk), .D (new_AGEMA_signal_1160), .Q (new_AGEMA_signal_1161) ) ;
    buf_clk new_AGEMA_reg_buffer_380 ( .C (clk), .D (new_AGEMA_signal_1166), .Q (new_AGEMA_signal_1167) ) ;
    buf_clk new_AGEMA_reg_buffer_386 ( .C (clk), .D (new_AGEMA_signal_1172), .Q (new_AGEMA_signal_1173) ) ;
    buf_clk new_AGEMA_reg_buffer_392 ( .C (clk), .D (new_AGEMA_signal_1178), .Q (new_AGEMA_signal_1179) ) ;
    buf_clk new_AGEMA_reg_buffer_398 ( .C (clk), .D (new_AGEMA_signal_1184), .Q (new_AGEMA_signal_1185) ) ;
    buf_clk new_AGEMA_reg_buffer_404 ( .C (clk), .D (new_AGEMA_signal_1190), .Q (new_AGEMA_signal_1191) ) ;
    buf_clk new_AGEMA_reg_buffer_410 ( .C (clk), .D (new_AGEMA_signal_1196), .Q (new_AGEMA_signal_1197) ) ;
    buf_clk new_AGEMA_reg_buffer_416 ( .C (clk), .D (new_AGEMA_signal_1202), .Q (new_AGEMA_signal_1203) ) ;
    buf_clk new_AGEMA_reg_buffer_422 ( .C (clk), .D (new_AGEMA_signal_1208), .Q (new_AGEMA_signal_1209) ) ;
    buf_clk new_AGEMA_reg_buffer_428 ( .C (clk), .D (new_AGEMA_signal_1214), .Q (new_AGEMA_signal_1215) ) ;
    buf_clk new_AGEMA_reg_buffer_434 ( .C (clk), .D (new_AGEMA_signal_1220), .Q (new_AGEMA_signal_1221) ) ;
    buf_clk new_AGEMA_reg_buffer_440 ( .C (clk), .D (new_AGEMA_signal_1226), .Q (new_AGEMA_signal_1227) ) ;
    buf_clk new_AGEMA_reg_buffer_446 ( .C (clk), .D (new_AGEMA_signal_1232), .Q (new_AGEMA_signal_1233) ) ;
    buf_clk new_AGEMA_reg_buffer_452 ( .C (clk), .D (new_AGEMA_signal_1238), .Q (new_AGEMA_signal_1239) ) ;
    buf_clk new_AGEMA_reg_buffer_458 ( .C (clk), .D (new_AGEMA_signal_1244), .Q (new_AGEMA_signal_1245) ) ;
    buf_clk new_AGEMA_reg_buffer_464 ( .C (clk), .D (new_AGEMA_signal_1250), .Q (new_AGEMA_signal_1251) ) ;
    buf_clk new_AGEMA_reg_buffer_470 ( .C (clk), .D (new_AGEMA_signal_1256), .Q (new_AGEMA_signal_1257) ) ;
    buf_clk new_AGEMA_reg_buffer_476 ( .C (clk), .D (new_AGEMA_signal_1262), .Q (new_AGEMA_signal_1263) ) ;
    buf_clk new_AGEMA_reg_buffer_482 ( .C (clk), .D (new_AGEMA_signal_1268), .Q (new_AGEMA_signal_1269) ) ;
    buf_clk new_AGEMA_reg_buffer_488 ( .C (clk), .D (new_AGEMA_signal_1274), .Q (new_AGEMA_signal_1275) ) ;
    buf_clk new_AGEMA_reg_buffer_494 ( .C (clk), .D (new_AGEMA_signal_1280), .Q (new_AGEMA_signal_1281) ) ;
    buf_clk new_AGEMA_reg_buffer_500 ( .C (clk), .D (new_AGEMA_signal_1286), .Q (new_AGEMA_signal_1287) ) ;
    buf_clk new_AGEMA_reg_buffer_506 ( .C (clk), .D (new_AGEMA_signal_1292), .Q (new_AGEMA_signal_1293) ) ;
    buf_clk new_AGEMA_reg_buffer_512 ( .C (clk), .D (new_AGEMA_signal_1298), .Q (new_AGEMA_signal_1299) ) ;
    buf_clk new_AGEMA_reg_buffer_518 ( .C (clk), .D (new_AGEMA_signal_1304), .Q (new_AGEMA_signal_1305) ) ;
    buf_clk new_AGEMA_reg_buffer_524 ( .C (clk), .D (new_AGEMA_signal_1310), .Q (new_AGEMA_signal_1311) ) ;
    buf_clk new_AGEMA_reg_buffer_530 ( .C (clk), .D (new_AGEMA_signal_1316), .Q (new_AGEMA_signal_1317) ) ;
    buf_clk new_AGEMA_reg_buffer_536 ( .C (clk), .D (new_AGEMA_signal_1322), .Q (new_AGEMA_signal_1323) ) ;
    buf_clk new_AGEMA_reg_buffer_542 ( .C (clk), .D (new_AGEMA_signal_1328), .Q (new_AGEMA_signal_1329) ) ;
    buf_clk new_AGEMA_reg_buffer_548 ( .C (clk), .D (new_AGEMA_signal_1334), .Q (new_AGEMA_signal_1335) ) ;
    buf_clk new_AGEMA_reg_buffer_554 ( .C (clk), .D (new_AGEMA_signal_1340), .Q (new_AGEMA_signal_1341) ) ;
    buf_clk new_AGEMA_reg_buffer_560 ( .C (clk), .D (new_AGEMA_signal_1346), .Q (new_AGEMA_signal_1347) ) ;
    buf_clk new_AGEMA_reg_buffer_566 ( .C (clk), .D (new_AGEMA_signal_1352), .Q (new_AGEMA_signal_1353) ) ;
    buf_clk new_AGEMA_reg_buffer_572 ( .C (clk), .D (new_AGEMA_signal_1358), .Q (new_AGEMA_signal_1359) ) ;
    buf_clk new_AGEMA_reg_buffer_578 ( .C (clk), .D (new_AGEMA_signal_1364), .Q (new_AGEMA_signal_1365) ) ;
    buf_clk new_AGEMA_reg_buffer_584 ( .C (clk), .D (new_AGEMA_signal_1370), .Q (new_AGEMA_signal_1371) ) ;
    buf_clk new_AGEMA_reg_buffer_590 ( .C (clk), .D (new_AGEMA_signal_1376), .Q (new_AGEMA_signal_1377) ) ;
    buf_clk new_AGEMA_reg_buffer_596 ( .C (clk), .D (new_AGEMA_signal_1382), .Q (new_AGEMA_signal_1383) ) ;
    buf_clk new_AGEMA_reg_buffer_602 ( .C (clk), .D (new_AGEMA_signal_1388), .Q (new_AGEMA_signal_1389) ) ;
    buf_clk new_AGEMA_reg_buffer_608 ( .C (clk), .D (new_AGEMA_signal_1394), .Q (new_AGEMA_signal_1395) ) ;
    buf_clk new_AGEMA_reg_buffer_614 ( .C (clk), .D (new_AGEMA_signal_1400), .Q (new_AGEMA_signal_1401) ) ;
    buf_clk new_AGEMA_reg_buffer_620 ( .C (clk), .D (new_AGEMA_signal_1406), .Q (new_AGEMA_signal_1407) ) ;
    buf_clk new_AGEMA_reg_buffer_626 ( .C (clk), .D (new_AGEMA_signal_1412), .Q (new_AGEMA_signal_1413) ) ;
    buf_clk new_AGEMA_reg_buffer_632 ( .C (clk), .D (new_AGEMA_signal_1418), .Q (new_AGEMA_signal_1419) ) ;
    buf_clk new_AGEMA_reg_buffer_638 ( .C (clk), .D (new_AGEMA_signal_1424), .Q (new_AGEMA_signal_1425) ) ;
    buf_clk new_AGEMA_reg_buffer_644 ( .C (clk), .D (new_AGEMA_signal_1430), .Q (new_AGEMA_signal_1431) ) ;
    buf_clk new_AGEMA_reg_buffer_650 ( .C (clk), .D (new_AGEMA_signal_1436), .Q (new_AGEMA_signal_1437) ) ;
    buf_clk new_AGEMA_reg_buffer_656 ( .C (clk), .D (new_AGEMA_signal_1442), .Q (new_AGEMA_signal_1443) ) ;
    buf_clk new_AGEMA_reg_buffer_662 ( .C (clk), .D (new_AGEMA_signal_1448), .Q (new_AGEMA_signal_1449) ) ;

    /* cells in depth 6 */
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M29_U1 ( .ina ({new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, M28}), .inb ({new_AGEMA_signal_978, new_AGEMA_signal_976, new_AGEMA_signal_974, new_AGEMA_signal_972}), .clk (clk), .rnd ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .outt ({new_AGEMA_signal_351, new_AGEMA_signal_350, new_AGEMA_signal_349, M29}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M30_U1 ( .ina ({new_AGEMA_signal_339, new_AGEMA_signal_338, new_AGEMA_signal_337, M26}), .inb ({new_AGEMA_signal_986, new_AGEMA_signal_984, new_AGEMA_signal_982, new_AGEMA_signal_980}), .clk (clk), .rnd ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .outt ({new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, M30}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M32_U1 ( .ina ({new_AGEMA_signal_978, new_AGEMA_signal_976, new_AGEMA_signal_974, new_AGEMA_signal_972}), .inb ({new_AGEMA_signal_345, new_AGEMA_signal_344, new_AGEMA_signal_343, M31}), .clk (clk), .rnd ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .outt ({new_AGEMA_signal_357, new_AGEMA_signal_356, new_AGEMA_signal_355, M32}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M35_U1 ( .ina ({new_AGEMA_signal_986, new_AGEMA_signal_984, new_AGEMA_signal_982, new_AGEMA_signal_980}), .inb ({new_AGEMA_signal_333, new_AGEMA_signal_332, new_AGEMA_signal_331, M34}), .clk (clk), .rnd ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .outt ({new_AGEMA_signal_360, new_AGEMA_signal_359, new_AGEMA_signal_358, M35}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M37_U1 ( .a ({new_AGEMA_signal_994, new_AGEMA_signal_992, new_AGEMA_signal_990, new_AGEMA_signal_988}), .b ({new_AGEMA_signal_351, new_AGEMA_signal_350, new_AGEMA_signal_349, M29}), .c ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, M37}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M38_U1 ( .a ({new_AGEMA_signal_357, new_AGEMA_signal_356, new_AGEMA_signal_355, M32}), .b ({new_AGEMA_signal_1002, new_AGEMA_signal_1000, new_AGEMA_signal_998, new_AGEMA_signal_996}), .c ({new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M38}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M39_U1 ( .a ({new_AGEMA_signal_1010, new_AGEMA_signal_1008, new_AGEMA_signal_1006, new_AGEMA_signal_1004}), .b ({new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, M30}), .c ({new_AGEMA_signal_372, new_AGEMA_signal_371, new_AGEMA_signal_370, M39}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M40_U1 ( .a ({new_AGEMA_signal_360, new_AGEMA_signal_359, new_AGEMA_signal_358, M35}), .b ({new_AGEMA_signal_1018, new_AGEMA_signal_1016, new_AGEMA_signal_1014, new_AGEMA_signal_1012}), .c ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, M40}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M41_U1 ( .a ({new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M38}), .b ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, M40}), .c ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, M41}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M42_U1 ( .a ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, M37}), .b ({new_AGEMA_signal_372, new_AGEMA_signal_371, new_AGEMA_signal_370, M39}), .c ({new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M42}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M43_U1 ( .a ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, M37}), .b ({new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M38}), .c ({new_AGEMA_signal_384, new_AGEMA_signal_383, new_AGEMA_signal_382, M43}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M44_U1 ( .a ({new_AGEMA_signal_372, new_AGEMA_signal_371, new_AGEMA_signal_370, M39}), .b ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, M40}), .c ({new_AGEMA_signal_387, new_AGEMA_signal_386, new_AGEMA_signal_385, M44}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_M45_U1 ( .a ({new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M42}), .b ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, M41}), .c ({new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, M45}) ) ;
    buf_clk new_AGEMA_reg_buffer_201 ( .C (clk), .D (new_AGEMA_signal_987), .Q (new_AGEMA_signal_988) ) ;
    buf_clk new_AGEMA_reg_buffer_203 ( .C (clk), .D (new_AGEMA_signal_989), .Q (new_AGEMA_signal_990) ) ;
    buf_clk new_AGEMA_reg_buffer_205 ( .C (clk), .D (new_AGEMA_signal_991), .Q (new_AGEMA_signal_992) ) ;
    buf_clk new_AGEMA_reg_buffer_207 ( .C (clk), .D (new_AGEMA_signal_993), .Q (new_AGEMA_signal_994) ) ;
    buf_clk new_AGEMA_reg_buffer_209 ( .C (clk), .D (new_AGEMA_signal_995), .Q (new_AGEMA_signal_996) ) ;
    buf_clk new_AGEMA_reg_buffer_211 ( .C (clk), .D (new_AGEMA_signal_997), .Q (new_AGEMA_signal_998) ) ;
    buf_clk new_AGEMA_reg_buffer_213 ( .C (clk), .D (new_AGEMA_signal_999), .Q (new_AGEMA_signal_1000) ) ;
    buf_clk new_AGEMA_reg_buffer_215 ( .C (clk), .D (new_AGEMA_signal_1001), .Q (new_AGEMA_signal_1002) ) ;
    buf_clk new_AGEMA_reg_buffer_217 ( .C (clk), .D (new_AGEMA_signal_1003), .Q (new_AGEMA_signal_1004) ) ;
    buf_clk new_AGEMA_reg_buffer_219 ( .C (clk), .D (new_AGEMA_signal_1005), .Q (new_AGEMA_signal_1006) ) ;
    buf_clk new_AGEMA_reg_buffer_221 ( .C (clk), .D (new_AGEMA_signal_1007), .Q (new_AGEMA_signal_1008) ) ;
    buf_clk new_AGEMA_reg_buffer_223 ( .C (clk), .D (new_AGEMA_signal_1009), .Q (new_AGEMA_signal_1010) ) ;
    buf_clk new_AGEMA_reg_buffer_225 ( .C (clk), .D (new_AGEMA_signal_1011), .Q (new_AGEMA_signal_1012) ) ;
    buf_clk new_AGEMA_reg_buffer_227 ( .C (clk), .D (new_AGEMA_signal_1013), .Q (new_AGEMA_signal_1014) ) ;
    buf_clk new_AGEMA_reg_buffer_229 ( .C (clk), .D (new_AGEMA_signal_1015), .Q (new_AGEMA_signal_1016) ) ;
    buf_clk new_AGEMA_reg_buffer_231 ( .C (clk), .D (new_AGEMA_signal_1017), .Q (new_AGEMA_signal_1018) ) ;
    buf_clk new_AGEMA_reg_buffer_237 ( .C (clk), .D (new_AGEMA_signal_1023), .Q (new_AGEMA_signal_1024) ) ;
    buf_clk new_AGEMA_reg_buffer_243 ( .C (clk), .D (new_AGEMA_signal_1029), .Q (new_AGEMA_signal_1030) ) ;
    buf_clk new_AGEMA_reg_buffer_249 ( .C (clk), .D (new_AGEMA_signal_1035), .Q (new_AGEMA_signal_1036) ) ;
    buf_clk new_AGEMA_reg_buffer_255 ( .C (clk), .D (new_AGEMA_signal_1041), .Q (new_AGEMA_signal_1042) ) ;
    buf_clk new_AGEMA_reg_buffer_261 ( .C (clk), .D (new_AGEMA_signal_1047), .Q (new_AGEMA_signal_1048) ) ;
    buf_clk new_AGEMA_reg_buffer_267 ( .C (clk), .D (new_AGEMA_signal_1053), .Q (new_AGEMA_signal_1054) ) ;
    buf_clk new_AGEMA_reg_buffer_273 ( .C (clk), .D (new_AGEMA_signal_1059), .Q (new_AGEMA_signal_1060) ) ;
    buf_clk new_AGEMA_reg_buffer_279 ( .C (clk), .D (new_AGEMA_signal_1065), .Q (new_AGEMA_signal_1066) ) ;
    buf_clk new_AGEMA_reg_buffer_285 ( .C (clk), .D (new_AGEMA_signal_1071), .Q (new_AGEMA_signal_1072) ) ;
    buf_clk new_AGEMA_reg_buffer_291 ( .C (clk), .D (new_AGEMA_signal_1077), .Q (new_AGEMA_signal_1078) ) ;
    buf_clk new_AGEMA_reg_buffer_297 ( .C (clk), .D (new_AGEMA_signal_1083), .Q (new_AGEMA_signal_1084) ) ;
    buf_clk new_AGEMA_reg_buffer_303 ( .C (clk), .D (new_AGEMA_signal_1089), .Q (new_AGEMA_signal_1090) ) ;
    buf_clk new_AGEMA_reg_buffer_309 ( .C (clk), .D (new_AGEMA_signal_1095), .Q (new_AGEMA_signal_1096) ) ;
    buf_clk new_AGEMA_reg_buffer_315 ( .C (clk), .D (new_AGEMA_signal_1101), .Q (new_AGEMA_signal_1102) ) ;
    buf_clk new_AGEMA_reg_buffer_321 ( .C (clk), .D (new_AGEMA_signal_1107), .Q (new_AGEMA_signal_1108) ) ;
    buf_clk new_AGEMA_reg_buffer_327 ( .C (clk), .D (new_AGEMA_signal_1113), .Q (new_AGEMA_signal_1114) ) ;
    buf_clk new_AGEMA_reg_buffer_333 ( .C (clk), .D (new_AGEMA_signal_1119), .Q (new_AGEMA_signal_1120) ) ;
    buf_clk new_AGEMA_reg_buffer_339 ( .C (clk), .D (new_AGEMA_signal_1125), .Q (new_AGEMA_signal_1126) ) ;
    buf_clk new_AGEMA_reg_buffer_345 ( .C (clk), .D (new_AGEMA_signal_1131), .Q (new_AGEMA_signal_1132) ) ;
    buf_clk new_AGEMA_reg_buffer_351 ( .C (clk), .D (new_AGEMA_signal_1137), .Q (new_AGEMA_signal_1138) ) ;
    buf_clk new_AGEMA_reg_buffer_357 ( .C (clk), .D (new_AGEMA_signal_1143), .Q (new_AGEMA_signal_1144) ) ;
    buf_clk new_AGEMA_reg_buffer_363 ( .C (clk), .D (new_AGEMA_signal_1149), .Q (new_AGEMA_signal_1150) ) ;
    buf_clk new_AGEMA_reg_buffer_369 ( .C (clk), .D (new_AGEMA_signal_1155), .Q (new_AGEMA_signal_1156) ) ;
    buf_clk new_AGEMA_reg_buffer_375 ( .C (clk), .D (new_AGEMA_signal_1161), .Q (new_AGEMA_signal_1162) ) ;
    buf_clk new_AGEMA_reg_buffer_381 ( .C (clk), .D (new_AGEMA_signal_1167), .Q (new_AGEMA_signal_1168) ) ;
    buf_clk new_AGEMA_reg_buffer_387 ( .C (clk), .D (new_AGEMA_signal_1173), .Q (new_AGEMA_signal_1174) ) ;
    buf_clk new_AGEMA_reg_buffer_393 ( .C (clk), .D (new_AGEMA_signal_1179), .Q (new_AGEMA_signal_1180) ) ;
    buf_clk new_AGEMA_reg_buffer_399 ( .C (clk), .D (new_AGEMA_signal_1185), .Q (new_AGEMA_signal_1186) ) ;
    buf_clk new_AGEMA_reg_buffer_405 ( .C (clk), .D (new_AGEMA_signal_1191), .Q (new_AGEMA_signal_1192) ) ;
    buf_clk new_AGEMA_reg_buffer_411 ( .C (clk), .D (new_AGEMA_signal_1197), .Q (new_AGEMA_signal_1198) ) ;
    buf_clk new_AGEMA_reg_buffer_417 ( .C (clk), .D (new_AGEMA_signal_1203), .Q (new_AGEMA_signal_1204) ) ;
    buf_clk new_AGEMA_reg_buffer_423 ( .C (clk), .D (new_AGEMA_signal_1209), .Q (new_AGEMA_signal_1210) ) ;
    buf_clk new_AGEMA_reg_buffer_429 ( .C (clk), .D (new_AGEMA_signal_1215), .Q (new_AGEMA_signal_1216) ) ;
    buf_clk new_AGEMA_reg_buffer_435 ( .C (clk), .D (new_AGEMA_signal_1221), .Q (new_AGEMA_signal_1222) ) ;
    buf_clk new_AGEMA_reg_buffer_441 ( .C (clk), .D (new_AGEMA_signal_1227), .Q (new_AGEMA_signal_1228) ) ;
    buf_clk new_AGEMA_reg_buffer_447 ( .C (clk), .D (new_AGEMA_signal_1233), .Q (new_AGEMA_signal_1234) ) ;
    buf_clk new_AGEMA_reg_buffer_453 ( .C (clk), .D (new_AGEMA_signal_1239), .Q (new_AGEMA_signal_1240) ) ;
    buf_clk new_AGEMA_reg_buffer_459 ( .C (clk), .D (new_AGEMA_signal_1245), .Q (new_AGEMA_signal_1246) ) ;
    buf_clk new_AGEMA_reg_buffer_465 ( .C (clk), .D (new_AGEMA_signal_1251), .Q (new_AGEMA_signal_1252) ) ;
    buf_clk new_AGEMA_reg_buffer_471 ( .C (clk), .D (new_AGEMA_signal_1257), .Q (new_AGEMA_signal_1258) ) ;
    buf_clk new_AGEMA_reg_buffer_477 ( .C (clk), .D (new_AGEMA_signal_1263), .Q (new_AGEMA_signal_1264) ) ;
    buf_clk new_AGEMA_reg_buffer_483 ( .C (clk), .D (new_AGEMA_signal_1269), .Q (new_AGEMA_signal_1270) ) ;
    buf_clk new_AGEMA_reg_buffer_489 ( .C (clk), .D (new_AGEMA_signal_1275), .Q (new_AGEMA_signal_1276) ) ;
    buf_clk new_AGEMA_reg_buffer_495 ( .C (clk), .D (new_AGEMA_signal_1281), .Q (new_AGEMA_signal_1282) ) ;
    buf_clk new_AGEMA_reg_buffer_501 ( .C (clk), .D (new_AGEMA_signal_1287), .Q (new_AGEMA_signal_1288) ) ;
    buf_clk new_AGEMA_reg_buffer_507 ( .C (clk), .D (new_AGEMA_signal_1293), .Q (new_AGEMA_signal_1294) ) ;
    buf_clk new_AGEMA_reg_buffer_513 ( .C (clk), .D (new_AGEMA_signal_1299), .Q (new_AGEMA_signal_1300) ) ;
    buf_clk new_AGEMA_reg_buffer_519 ( .C (clk), .D (new_AGEMA_signal_1305), .Q (new_AGEMA_signal_1306) ) ;
    buf_clk new_AGEMA_reg_buffer_525 ( .C (clk), .D (new_AGEMA_signal_1311), .Q (new_AGEMA_signal_1312) ) ;
    buf_clk new_AGEMA_reg_buffer_531 ( .C (clk), .D (new_AGEMA_signal_1317), .Q (new_AGEMA_signal_1318) ) ;
    buf_clk new_AGEMA_reg_buffer_537 ( .C (clk), .D (new_AGEMA_signal_1323), .Q (new_AGEMA_signal_1324) ) ;
    buf_clk new_AGEMA_reg_buffer_543 ( .C (clk), .D (new_AGEMA_signal_1329), .Q (new_AGEMA_signal_1330) ) ;
    buf_clk new_AGEMA_reg_buffer_549 ( .C (clk), .D (new_AGEMA_signal_1335), .Q (new_AGEMA_signal_1336) ) ;
    buf_clk new_AGEMA_reg_buffer_555 ( .C (clk), .D (new_AGEMA_signal_1341), .Q (new_AGEMA_signal_1342) ) ;
    buf_clk new_AGEMA_reg_buffer_561 ( .C (clk), .D (new_AGEMA_signal_1347), .Q (new_AGEMA_signal_1348) ) ;
    buf_clk new_AGEMA_reg_buffer_567 ( .C (clk), .D (new_AGEMA_signal_1353), .Q (new_AGEMA_signal_1354) ) ;
    buf_clk new_AGEMA_reg_buffer_573 ( .C (clk), .D (new_AGEMA_signal_1359), .Q (new_AGEMA_signal_1360) ) ;
    buf_clk new_AGEMA_reg_buffer_579 ( .C (clk), .D (new_AGEMA_signal_1365), .Q (new_AGEMA_signal_1366) ) ;
    buf_clk new_AGEMA_reg_buffer_585 ( .C (clk), .D (new_AGEMA_signal_1371), .Q (new_AGEMA_signal_1372) ) ;
    buf_clk new_AGEMA_reg_buffer_591 ( .C (clk), .D (new_AGEMA_signal_1377), .Q (new_AGEMA_signal_1378) ) ;
    buf_clk new_AGEMA_reg_buffer_597 ( .C (clk), .D (new_AGEMA_signal_1383), .Q (new_AGEMA_signal_1384) ) ;
    buf_clk new_AGEMA_reg_buffer_603 ( .C (clk), .D (new_AGEMA_signal_1389), .Q (new_AGEMA_signal_1390) ) ;
    buf_clk new_AGEMA_reg_buffer_609 ( .C (clk), .D (new_AGEMA_signal_1395), .Q (new_AGEMA_signal_1396) ) ;
    buf_clk new_AGEMA_reg_buffer_615 ( .C (clk), .D (new_AGEMA_signal_1401), .Q (new_AGEMA_signal_1402) ) ;
    buf_clk new_AGEMA_reg_buffer_621 ( .C (clk), .D (new_AGEMA_signal_1407), .Q (new_AGEMA_signal_1408) ) ;
    buf_clk new_AGEMA_reg_buffer_627 ( .C (clk), .D (new_AGEMA_signal_1413), .Q (new_AGEMA_signal_1414) ) ;
    buf_clk new_AGEMA_reg_buffer_633 ( .C (clk), .D (new_AGEMA_signal_1419), .Q (new_AGEMA_signal_1420) ) ;
    buf_clk new_AGEMA_reg_buffer_639 ( .C (clk), .D (new_AGEMA_signal_1425), .Q (new_AGEMA_signal_1426) ) ;
    buf_clk new_AGEMA_reg_buffer_645 ( .C (clk), .D (new_AGEMA_signal_1431), .Q (new_AGEMA_signal_1432) ) ;
    buf_clk new_AGEMA_reg_buffer_651 ( .C (clk), .D (new_AGEMA_signal_1437), .Q (new_AGEMA_signal_1438) ) ;
    buf_clk new_AGEMA_reg_buffer_657 ( .C (clk), .D (new_AGEMA_signal_1443), .Q (new_AGEMA_signal_1444) ) ;
    buf_clk new_AGEMA_reg_buffer_663 ( .C (clk), .D (new_AGEMA_signal_1449), .Q (new_AGEMA_signal_1450) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M46_U1 ( .ina ({new_AGEMA_signal_387, new_AGEMA_signal_386, new_AGEMA_signal_385, M44}), .inb ({new_AGEMA_signal_1042, new_AGEMA_signal_1036, new_AGEMA_signal_1030, new_AGEMA_signal_1024}), .clk (clk), .rnd ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .outt ({new_AGEMA_signal_417, new_AGEMA_signal_416, new_AGEMA_signal_415, M46}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M47_U1 ( .ina ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, M40}), .inb ({new_AGEMA_signal_1066, new_AGEMA_signal_1060, new_AGEMA_signal_1054, new_AGEMA_signal_1048}), .clk (clk), .rnd ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .outt ({new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, M47}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M48_U1 ( .ina ({new_AGEMA_signal_372, new_AGEMA_signal_371, new_AGEMA_signal_370, M39}), .inb ({new_AGEMA_signal_1090, new_AGEMA_signal_1084, new_AGEMA_signal_1078, new_AGEMA_signal_1072}), .clk (clk), .rnd ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .outt ({new_AGEMA_signal_393, new_AGEMA_signal_392, new_AGEMA_signal_391, M48}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M49_U1 ( .ina ({new_AGEMA_signal_384, new_AGEMA_signal_383, new_AGEMA_signal_382, M43}), .inb ({new_AGEMA_signal_1114, new_AGEMA_signal_1108, new_AGEMA_signal_1102, new_AGEMA_signal_1096}), .clk (clk), .rnd ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .outt ({new_AGEMA_signal_420, new_AGEMA_signal_419, new_AGEMA_signal_418, M49}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M50_U1 ( .ina ({new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M38}), .inb ({new_AGEMA_signal_1138, new_AGEMA_signal_1132, new_AGEMA_signal_1126, new_AGEMA_signal_1120}), .clk (clk), .rnd ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .outt ({new_AGEMA_signal_396, new_AGEMA_signal_395, new_AGEMA_signal_394, M50}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M51_U1 ( .ina ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, M37}), .inb ({new_AGEMA_signal_1162, new_AGEMA_signal_1156, new_AGEMA_signal_1150, new_AGEMA_signal_1144}), .clk (clk), .rnd ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .outt ({new_AGEMA_signal_399, new_AGEMA_signal_398, new_AGEMA_signal_397, M51}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M52_U1 ( .ina ({new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M42}), .inb ({new_AGEMA_signal_1186, new_AGEMA_signal_1180, new_AGEMA_signal_1174, new_AGEMA_signal_1168}), .clk (clk), .rnd ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .outt ({new_AGEMA_signal_423, new_AGEMA_signal_422, new_AGEMA_signal_421, M52}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M53_U1 ( .ina ({new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, M45}), .inb ({new_AGEMA_signal_1210, new_AGEMA_signal_1204, new_AGEMA_signal_1198, new_AGEMA_signal_1192}), .clk (clk), .rnd ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .outt ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, M53}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M54_U1 ( .ina ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, M41}), .inb ({new_AGEMA_signal_1234, new_AGEMA_signal_1228, new_AGEMA_signal_1222, new_AGEMA_signal_1216}), .clk (clk), .rnd ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .outt ({new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, M54}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M55_U1 ( .ina ({new_AGEMA_signal_387, new_AGEMA_signal_386, new_AGEMA_signal_385, M44}), .inb ({new_AGEMA_signal_1258, new_AGEMA_signal_1252, new_AGEMA_signal_1246, new_AGEMA_signal_1240}), .clk (clk), .rnd ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .outt ({new_AGEMA_signal_429, new_AGEMA_signal_428, new_AGEMA_signal_427, M55}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M56_U1 ( .ina ({new_AGEMA_signal_375, new_AGEMA_signal_374, new_AGEMA_signal_373, M40}), .inb ({new_AGEMA_signal_1282, new_AGEMA_signal_1276, new_AGEMA_signal_1270, new_AGEMA_signal_1264}), .clk (clk), .rnd ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .outt ({new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, M56}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M57_U1 ( .ina ({new_AGEMA_signal_372, new_AGEMA_signal_371, new_AGEMA_signal_370, M39}), .inb ({new_AGEMA_signal_1306, new_AGEMA_signal_1300, new_AGEMA_signal_1294, new_AGEMA_signal_1288}), .clk (clk), .rnd ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .outt ({new_AGEMA_signal_405, new_AGEMA_signal_404, new_AGEMA_signal_403, M57}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M58_U1 ( .ina ({new_AGEMA_signal_384, new_AGEMA_signal_383, new_AGEMA_signal_382, M43}), .inb ({new_AGEMA_signal_1330, new_AGEMA_signal_1324, new_AGEMA_signal_1318, new_AGEMA_signal_1312}), .clk (clk), .rnd ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .outt ({new_AGEMA_signal_432, new_AGEMA_signal_431, new_AGEMA_signal_430, M58}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M59_U1 ( .ina ({new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M38}), .inb ({new_AGEMA_signal_1354, new_AGEMA_signal_1348, new_AGEMA_signal_1342, new_AGEMA_signal_1336}), .clk (clk), .rnd ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .outt ({new_AGEMA_signal_408, new_AGEMA_signal_407, new_AGEMA_signal_406, M59}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M60_U1 ( .ina ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, M37}), .inb ({new_AGEMA_signal_1378, new_AGEMA_signal_1372, new_AGEMA_signal_1366, new_AGEMA_signal_1360}), .clk (clk), .rnd ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .outt ({new_AGEMA_signal_411, new_AGEMA_signal_410, new_AGEMA_signal_409, M60}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M61_U1 ( .ina ({new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M42}), .inb ({new_AGEMA_signal_1402, new_AGEMA_signal_1396, new_AGEMA_signal_1390, new_AGEMA_signal_1384}), .clk (clk), .rnd ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .outt ({new_AGEMA_signal_435, new_AGEMA_signal_434, new_AGEMA_signal_433, M61}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M62_U1 ( .ina ({new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, M45}), .inb ({new_AGEMA_signal_1426, new_AGEMA_signal_1420, new_AGEMA_signal_1414, new_AGEMA_signal_1408}), .clk (clk), .rnd ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .outt ({new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M62}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) AND_M63_U1 ( .ina ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, M41}), .inb ({new_AGEMA_signal_1450, new_AGEMA_signal_1444, new_AGEMA_signal_1438, new_AGEMA_signal_1432}), .clk (clk), .rnd ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .outt ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, M63}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L0_U1 ( .a ({new_AGEMA_signal_435, new_AGEMA_signal_434, new_AGEMA_signal_433, M61}), .b ({new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M62}), .c ({new_AGEMA_signal_480, new_AGEMA_signal_479, new_AGEMA_signal_478, L0}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L1_U1 ( .a ({new_AGEMA_signal_396, new_AGEMA_signal_395, new_AGEMA_signal_394, M50}), .b ({new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, M56}), .c ({new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, L1}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L2_U1 ( .a ({new_AGEMA_signal_417, new_AGEMA_signal_416, new_AGEMA_signal_415, M46}), .b ({new_AGEMA_signal_393, new_AGEMA_signal_392, new_AGEMA_signal_391, M48}), .c ({new_AGEMA_signal_456, new_AGEMA_signal_455, new_AGEMA_signal_454, L2}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L3_U1 ( .a ({new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, M47}), .b ({new_AGEMA_signal_429, new_AGEMA_signal_428, new_AGEMA_signal_427, M55}), .c ({new_AGEMA_signal_459, new_AGEMA_signal_458, new_AGEMA_signal_457, L3}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L4_U1 ( .a ({new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, M54}), .b ({new_AGEMA_signal_432, new_AGEMA_signal_431, new_AGEMA_signal_430, M58}), .c ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, L4}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L5_U1 ( .a ({new_AGEMA_signal_420, new_AGEMA_signal_419, new_AGEMA_signal_418, M49}), .b ({new_AGEMA_signal_435, new_AGEMA_signal_434, new_AGEMA_signal_433, M61}), .c ({new_AGEMA_signal_465, new_AGEMA_signal_464, new_AGEMA_signal_463, L5}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L6_U1 ( .a ({new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M62}), .b ({new_AGEMA_signal_465, new_AGEMA_signal_464, new_AGEMA_signal_463, L5}), .c ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, L6}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L7_U1 ( .a ({new_AGEMA_signal_417, new_AGEMA_signal_416, new_AGEMA_signal_415, M46}), .b ({new_AGEMA_signal_459, new_AGEMA_signal_458, new_AGEMA_signal_457, L3}), .c ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, L7}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L8_U1 ( .a ({new_AGEMA_signal_399, new_AGEMA_signal_398, new_AGEMA_signal_397, M51}), .b ({new_AGEMA_signal_408, new_AGEMA_signal_407, new_AGEMA_signal_406, M59}), .c ({new_AGEMA_signal_444, new_AGEMA_signal_443, new_AGEMA_signal_442, L8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L9_U1 ( .a ({new_AGEMA_signal_423, new_AGEMA_signal_422, new_AGEMA_signal_421, M52}), .b ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, M53}), .c ({new_AGEMA_signal_489, new_AGEMA_signal_488, new_AGEMA_signal_487, L9}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L10_U1 ( .a ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, M53}), .b ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, L4}), .c ({new_AGEMA_signal_492, new_AGEMA_signal_491, new_AGEMA_signal_490, L10}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L11_U1 ( .a ({new_AGEMA_signal_411, new_AGEMA_signal_410, new_AGEMA_signal_409, M60}), .b ({new_AGEMA_signal_456, new_AGEMA_signal_455, new_AGEMA_signal_454, L2}), .c ({new_AGEMA_signal_495, new_AGEMA_signal_494, new_AGEMA_signal_493, L11}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L12_U1 ( .a ({new_AGEMA_signal_393, new_AGEMA_signal_392, new_AGEMA_signal_391, M48}), .b ({new_AGEMA_signal_399, new_AGEMA_signal_398, new_AGEMA_signal_397, M51}), .c ({new_AGEMA_signal_447, new_AGEMA_signal_446, new_AGEMA_signal_445, L12}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L13_U1 ( .a ({new_AGEMA_signal_396, new_AGEMA_signal_395, new_AGEMA_signal_394, M50}), .b ({new_AGEMA_signal_480, new_AGEMA_signal_479, new_AGEMA_signal_478, L0}), .c ({new_AGEMA_signal_507, new_AGEMA_signal_506, new_AGEMA_signal_505, L13}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L14_U1 ( .a ({new_AGEMA_signal_423, new_AGEMA_signal_422, new_AGEMA_signal_421, M52}), .b ({new_AGEMA_signal_435, new_AGEMA_signal_434, new_AGEMA_signal_433, M61}), .c ({new_AGEMA_signal_468, new_AGEMA_signal_467, new_AGEMA_signal_466, L14}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L15_U1 ( .a ({new_AGEMA_signal_429, new_AGEMA_signal_428, new_AGEMA_signal_427, M55}), .b ({new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, L1}), .c ({new_AGEMA_signal_471, new_AGEMA_signal_470, new_AGEMA_signal_469, L15}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L16_U1 ( .a ({new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, M56}), .b ({new_AGEMA_signal_480, new_AGEMA_signal_479, new_AGEMA_signal_478, L0}), .c ({new_AGEMA_signal_510, new_AGEMA_signal_509, new_AGEMA_signal_508, L16}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L17_U1 ( .a ({new_AGEMA_signal_405, new_AGEMA_signal_404, new_AGEMA_signal_403, M57}), .b ({new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, L1}), .c ({new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, L17}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L18_U1 ( .a ({new_AGEMA_signal_432, new_AGEMA_signal_431, new_AGEMA_signal_430, M58}), .b ({new_AGEMA_signal_444, new_AGEMA_signal_443, new_AGEMA_signal_442, L8}), .c ({new_AGEMA_signal_477, new_AGEMA_signal_476, new_AGEMA_signal_475, L18}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L19_U1 ( .a ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, M63}), .b ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, L4}), .c ({new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, L19}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L20_U1 ( .a ({new_AGEMA_signal_480, new_AGEMA_signal_479, new_AGEMA_signal_478, L0}), .b ({new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, L1}), .c ({new_AGEMA_signal_513, new_AGEMA_signal_512, new_AGEMA_signal_511, L20}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L21_U1 ( .a ({new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, L1}), .b ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, L7}), .c ({new_AGEMA_signal_516, new_AGEMA_signal_515, new_AGEMA_signal_514, L21}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L22_U1 ( .a ({new_AGEMA_signal_459, new_AGEMA_signal_458, new_AGEMA_signal_457, L3}), .b ({new_AGEMA_signal_447, new_AGEMA_signal_446, new_AGEMA_signal_445, L12}), .c ({new_AGEMA_signal_501, new_AGEMA_signal_500, new_AGEMA_signal_499, L22}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L23_U1 ( .a ({new_AGEMA_signal_477, new_AGEMA_signal_476, new_AGEMA_signal_475, L18}), .b ({new_AGEMA_signal_456, new_AGEMA_signal_455, new_AGEMA_signal_454, L2}), .c ({new_AGEMA_signal_504, new_AGEMA_signal_503, new_AGEMA_signal_502, L23}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L24_U1 ( .a ({new_AGEMA_signal_471, new_AGEMA_signal_470, new_AGEMA_signal_469, L15}), .b ({new_AGEMA_signal_489, new_AGEMA_signal_488, new_AGEMA_signal_487, L9}), .c ({new_AGEMA_signal_519, new_AGEMA_signal_518, new_AGEMA_signal_517, L24}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L25_U1 ( .a ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, L6}), .b ({new_AGEMA_signal_492, new_AGEMA_signal_491, new_AGEMA_signal_490, L10}), .c ({new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, L25}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L26_U1 ( .a ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, L7}), .b ({new_AGEMA_signal_489, new_AGEMA_signal_488, new_AGEMA_signal_487, L9}), .c ({new_AGEMA_signal_525, new_AGEMA_signal_524, new_AGEMA_signal_523, L26}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L27_U1 ( .a ({new_AGEMA_signal_444, new_AGEMA_signal_443, new_AGEMA_signal_442, L8}), .b ({new_AGEMA_signal_492, new_AGEMA_signal_491, new_AGEMA_signal_490, L10}), .c ({new_AGEMA_signal_528, new_AGEMA_signal_527, new_AGEMA_signal_526, L27}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L28_U1 ( .a ({new_AGEMA_signal_495, new_AGEMA_signal_494, new_AGEMA_signal_493, L11}), .b ({new_AGEMA_signal_468, new_AGEMA_signal_467, new_AGEMA_signal_466, L14}), .c ({new_AGEMA_signal_531, new_AGEMA_signal_530, new_AGEMA_signal_529, L28}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_L29_U1 ( .a ({new_AGEMA_signal_495, new_AGEMA_signal_494, new_AGEMA_signal_493, L11}), .b ({new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, L17}), .c ({new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, L29}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_S0_U1 ( .a ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, L6}), .b ({new_AGEMA_signal_519, new_AGEMA_signal_518, new_AGEMA_signal_517, L24}), .c ({new_AGEMA_signal_540, new_AGEMA_signal_539, new_AGEMA_signal_538, O[7]}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(1)) XOR_S1_U1 ( .a ({new_AGEMA_signal_510, new_AGEMA_signal_509, new_AGEMA_signal_508, L16}), .b ({new_AGEMA_signal_525, new_AGEMA_signal_524, new_AGEMA_signal_523, L26}), .c ({new_AGEMA_signal_543, new_AGEMA_signal_542, new_AGEMA_signal_541, O[6]}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(1)) XOR_S2_U1 ( .a ({new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, L19}), .b ({new_AGEMA_signal_531, new_AGEMA_signal_530, new_AGEMA_signal_529, L28}), .c ({new_AGEMA_signal_546, new_AGEMA_signal_545, new_AGEMA_signal_544, O[5]}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_S3_U1 ( .a ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, L6}), .b ({new_AGEMA_signal_516, new_AGEMA_signal_515, new_AGEMA_signal_514, L21}), .c ({new_AGEMA_signal_549, new_AGEMA_signal_548, new_AGEMA_signal_547, O[4]}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_S4_U1 ( .a ({new_AGEMA_signal_513, new_AGEMA_signal_512, new_AGEMA_signal_511, L20}), .b ({new_AGEMA_signal_501, new_AGEMA_signal_500, new_AGEMA_signal_499, L22}), .c ({new_AGEMA_signal_552, new_AGEMA_signal_551, new_AGEMA_signal_550, O[3]}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(1)) XOR_S5_U1 ( .a ({new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, L25}), .b ({new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, L29}), .c ({new_AGEMA_signal_555, new_AGEMA_signal_554, new_AGEMA_signal_553, O[2]}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(1)) XOR_S6_U1 ( .a ({new_AGEMA_signal_507, new_AGEMA_signal_506, new_AGEMA_signal_505, L13}), .b ({new_AGEMA_signal_528, new_AGEMA_signal_527, new_AGEMA_signal_526, L27}), .c ({new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, O[1]}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(1)) XOR_S7_U1 ( .a ({new_AGEMA_signal_483, new_AGEMA_signal_482, new_AGEMA_signal_481, L6}), .b ({new_AGEMA_signal_504, new_AGEMA_signal_503, new_AGEMA_signal_502, L23}), .c ({new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, O[0]}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_7_ ( .clk (clk), .D ({new_AGEMA_signal_540, new_AGEMA_signal_539, new_AGEMA_signal_538, O[7]}), .Q ({Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_6_ ( .clk (clk), .D ({new_AGEMA_signal_543, new_AGEMA_signal_542, new_AGEMA_signal_541, O[6]}), .Q ({Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_5_ ( .clk (clk), .D ({new_AGEMA_signal_546, new_AGEMA_signal_545, new_AGEMA_signal_544, O[5]}), .Q ({Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_4_ ( .clk (clk), .D ({new_AGEMA_signal_549, new_AGEMA_signal_548, new_AGEMA_signal_547, O[4]}), .Q ({Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_3_ ( .clk (clk), .D ({new_AGEMA_signal_552, new_AGEMA_signal_551, new_AGEMA_signal_550, O[3]}), .Q ({Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_2_ ( .clk (clk), .D ({new_AGEMA_signal_555, new_AGEMA_signal_554, new_AGEMA_signal_553, O[2]}), .Q ({Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_1_ ( .clk (clk), .D ({new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, O[1]}), .Q ({Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_0_ ( .clk (clk), .D ({new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, O[0]}), .Q ({Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
