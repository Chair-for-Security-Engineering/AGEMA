/* modified netlist. Source: module sbox in file Designs/SkinnySbox/AGEMA/sbox_opt_correct/sbox.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d4 (X_s0, clk, X_s1, X_s2, X_s3, X_s4, Fresh, Y_s0, Y_s1, Y_s2, Y_s3, Y_s4);
    input [3:0] X_s0 ;
    input clk ;
    input [3:0] X_s1 ;
    input [3:0] X_s2 ;
    input [3:0] X_s3 ;
    input [3:0] X_s4 ;
    input [39:0] Fresh ;
    output [3:0] Y_s0 ;
    output [3:0] Y_s1 ;
    output [3:0] Y_s2 ;
    output [3:0] Y_s3 ;
    output [3:0] Y_s4 ;
    wire signal_33 ;
    wire signal_34 ;
    wire signal_35 ;
    wire signal_36 ;
    wire signal_37 ;
    wire signal_38 ;
    wire signal_39 ;
    wire signal_40 ;
    wire signal_41 ;
    wire signal_42 ;
    wire signal_43 ;
    wire signal_44 ;
    wire signal_45 ;
    wire signal_46 ;
    wire signal_47 ;
    wire signal_48 ;
    wire signal_49 ;
    wire signal_50 ;
    wire signal_51 ;
    wire signal_52 ;
    wire signal_53 ;
    wire signal_54 ;
    wire signal_55 ;
    wire signal_56 ;
    wire signal_61 ;
    wire signal_62 ;
    wire signal_63 ;
    wire signal_64 ;
    wire signal_69 ;
    wire signal_70 ;
    wire signal_71 ;
    wire signal_72 ;
    wire signal_77 ;
    wire signal_78 ;
    wire signal_79 ;
    wire signal_80 ;
    wire signal_85 ;
    wire signal_86 ;
    wire signal_87 ;
    wire signal_88 ;
    wire signal_89 ;
    wire signal_90 ;
    wire signal_91 ;
    wire signal_92 ;
    wire signal_93 ;
    wire signal_94 ;
    wire signal_95 ;
    wire signal_96 ;
    wire signal_97 ;
    wire signal_98 ;
    wire signal_99 ;
    wire signal_100 ;
    wire signal_101 ;
    wire signal_102 ;
    wire signal_103 ;
    wire signal_104 ;
    wire signal_105 ;
    wire signal_106 ;
    wire signal_107 ;
    wire signal_108 ;
    wire signal_109 ;
    wire signal_110 ;
    wire signal_111 ;
    wire signal_112 ;
    wire signal_113 ;
    wire signal_114 ;
    wire signal_115 ;
    wire signal_116 ;
    wire signal_117 ;
    wire signal_118 ;
    wire signal_119 ;
    wire signal_120 ;
    wire signal_121 ;
    wire signal_122 ;
    wire signal_123 ;
    wire signal_124 ;
    wire signal_125 ;
    wire signal_126 ;
    wire signal_127 ;
    wire signal_128 ;
    wire signal_129 ;
    wire signal_130 ;
    wire signal_131 ;
    wire signal_132 ;
    wire signal_133 ;
    wire signal_134 ;
    wire signal_135 ;
    wire signal_136 ;
    wire signal_137 ;
    wire signal_138 ;
    wire signal_139 ;
    wire signal_140 ;
    wire signal_141 ;
    wire signal_142 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;

    /* cells in depth 0 */
    not_masked #(.security_order(4), .pipeline(1)) cell_26 ( .a ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_64, signal_63, signal_62, signal_61, signal_37}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_27 ( .a ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_72, signal_71, signal_70, signal_69, signal_38}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_28 ( .a ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_80, signal_79, signal_78, signal_77, signal_39}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_29 ( .a ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_88, signal_87, signal_86, signal_85, signal_40}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_31 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_80, signal_79, signal_78, signal_77, signal_39}), .c ({signal_96, signal_95, signal_94, signal_93, signal_42}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_32 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_72, signal_71, signal_70, signal_69, signal_38}), .c ({signal_100, signal_99, signal_98, signal_97, signal_43}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_33 ( .a ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_80, signal_79, signal_78, signal_77, signal_39}), .c ({signal_104, signal_103, signal_102, signal_101, signal_44}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_34 ( .a ({signal_104, signal_103, signal_102, signal_101, signal_44}), .b ({signal_108, signal_107, signal_106, signal_105, signal_45}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_36 ( .a ({signal_100, signal_99, signal_98, signal_97, signal_43}), .b ({signal_104, signal_103, signal_102, signal_101, signal_44}), .c ({signal_116, signal_115, signal_114, signal_113, signal_47}) ) ;

    /* cells in depth 1 */
    buf_clk cell_50 ( .C (clk), .D (signal_38), .Q (signal_225) ) ;
    buf_clk cell_52 ( .C (clk), .D (signal_69), .Q (signal_227) ) ;
    buf_clk cell_54 ( .C (clk), .D (signal_70), .Q (signal_229) ) ;
    buf_clk cell_56 ( .C (clk), .D (signal_71), .Q (signal_231) ) ;
    buf_clk cell_58 ( .C (clk), .D (signal_72), .Q (signal_233) ) ;
    buf_clk cell_60 ( .C (clk), .D (signal_42), .Q (signal_235) ) ;
    buf_clk cell_62 ( .C (clk), .D (signal_93), .Q (signal_237) ) ;
    buf_clk cell_64 ( .C (clk), .D (signal_94), .Q (signal_239) ) ;
    buf_clk cell_66 ( .C (clk), .D (signal_95), .Q (signal_241) ) ;
    buf_clk cell_68 ( .C (clk), .D (signal_96), .Q (signal_243) ) ;
    buf_clk cell_70 ( .C (clk), .D (signal_47), .Q (signal_245) ) ;
    buf_clk cell_72 ( .C (clk), .D (signal_113), .Q (signal_247) ) ;
    buf_clk cell_74 ( .C (clk), .D (signal_114), .Q (signal_249) ) ;
    buf_clk cell_76 ( .C (clk), .D (signal_115), .Q (signal_251) ) ;
    buf_clk cell_78 ( .C (clk), .D (signal_116), .Q (signal_253) ) ;
    buf_clk cell_80 ( .C (clk), .D (signal_39), .Q (signal_255) ) ;
    buf_clk cell_82 ( .C (clk), .D (signal_77), .Q (signal_257) ) ;
    buf_clk cell_84 ( .C (clk), .D (signal_78), .Q (signal_259) ) ;
    buf_clk cell_86 ( .C (clk), .D (signal_79), .Q (signal_261) ) ;
    buf_clk cell_88 ( .C (clk), .D (signal_80), .Q (signal_263) ) ;
    buf_clk cell_90 ( .C (clk), .D (X_s0[1]), .Q (signal_265) ) ;
    buf_clk cell_92 ( .C (clk), .D (X_s1[1]), .Q (signal_267) ) ;
    buf_clk cell_94 ( .C (clk), .D (X_s2[1]), .Q (signal_269) ) ;
    buf_clk cell_96 ( .C (clk), .D (X_s3[1]), .Q (signal_271) ) ;
    buf_clk cell_98 ( .C (clk), .D (X_s4[1]), .Q (signal_273) ) ;
    buf_clk cell_100 ( .C (clk), .D (signal_45), .Q (signal_275) ) ;
    buf_clk cell_102 ( .C (clk), .D (signal_105), .Q (signal_277) ) ;
    buf_clk cell_104 ( .C (clk), .D (signal_106), .Q (signal_279) ) ;
    buf_clk cell_106 ( .C (clk), .D (signal_107), .Q (signal_281) ) ;
    buf_clk cell_108 ( .C (clk), .D (signal_108), .Q (signal_283) ) ;
    buf_clk cell_120 ( .C (clk), .D (signal_40), .Q (signal_295) ) ;
    buf_clk cell_124 ( .C (clk), .D (signal_85), .Q (signal_299) ) ;
    buf_clk cell_128 ( .C (clk), .D (signal_86), .Q (signal_303) ) ;
    buf_clk cell_132 ( .C (clk), .D (signal_87), .Q (signal_307) ) ;
    buf_clk cell_136 ( .C (clk), .D (signal_88), .Q (signal_311) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_30 ( .a ({signal_64, signal_63, signal_62, signal_61, signal_37}), .b ({signal_88, signal_87, signal_86, signal_85, signal_40}), .clk (clk), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_92, signal_91, signal_90, signal_89, signal_41}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_35 ( .a ({signal_64, signal_63, signal_62, signal_61, signal_37}), .b ({signal_100, signal_99, signal_98, signal_97, signal_43}), .clk (clk), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({signal_112, signal_111, signal_110, signal_109, signal_46}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_37 ( .a ({signal_234, signal_232, signal_230, signal_228, signal_226}), .b ({signal_92, signal_91, signal_90, signal_89, signal_41}), .c ({signal_120, signal_119, signal_118, signal_117, signal_48}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_38 ( .a ({signal_120, signal_119, signal_118, signal_117, signal_48}), .b ({signal_124, signal_123, signal_122, signal_121, signal_36}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_39 ( .a ({signal_244, signal_242, signal_240, signal_238, signal_236}), .b ({signal_112, signal_111, signal_110, signal_109, signal_46}), .c ({signal_128, signal_127, signal_126, signal_125, signal_49}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_40 ( .a ({signal_92, signal_91, signal_90, signal_89, signal_41}), .b ({signal_254, signal_252, signal_250, signal_248, signal_246}), .c ({signal_132, signal_131, signal_130, signal_129, signal_50}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_41 ( .a ({signal_264, signal_262, signal_260, signal_258, signal_256}), .b ({signal_112, signal_111, signal_110, signal_109, signal_46}), .c ({signal_136, signal_135, signal_134, signal_133, signal_51}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_44 ( .a ({signal_92, signal_91, signal_90, signal_89, signal_41}), .b ({signal_136, signal_135, signal_134, signal_133, signal_51}), .c ({signal_148, signal_147, signal_146, signal_145, signal_54}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_45 ( .a ({signal_148, signal_147, signal_146, signal_145, signal_54}), .b ({signal_152, signal_151, signal_150, signal_149, signal_35}) ) ;
    buf_clk cell_51 ( .C (clk), .D (signal_225), .Q (signal_226) ) ;
    buf_clk cell_53 ( .C (clk), .D (signal_227), .Q (signal_228) ) ;
    buf_clk cell_55 ( .C (clk), .D (signal_229), .Q (signal_230) ) ;
    buf_clk cell_57 ( .C (clk), .D (signal_231), .Q (signal_232) ) ;
    buf_clk cell_59 ( .C (clk), .D (signal_233), .Q (signal_234) ) ;
    buf_clk cell_61 ( .C (clk), .D (signal_235), .Q (signal_236) ) ;
    buf_clk cell_63 ( .C (clk), .D (signal_237), .Q (signal_238) ) ;
    buf_clk cell_65 ( .C (clk), .D (signal_239), .Q (signal_240) ) ;
    buf_clk cell_67 ( .C (clk), .D (signal_241), .Q (signal_242) ) ;
    buf_clk cell_69 ( .C (clk), .D (signal_243), .Q (signal_244) ) ;
    buf_clk cell_71 ( .C (clk), .D (signal_245), .Q (signal_246) ) ;
    buf_clk cell_73 ( .C (clk), .D (signal_247), .Q (signal_248) ) ;
    buf_clk cell_75 ( .C (clk), .D (signal_249), .Q (signal_250) ) ;
    buf_clk cell_77 ( .C (clk), .D (signal_251), .Q (signal_252) ) ;
    buf_clk cell_79 ( .C (clk), .D (signal_253), .Q (signal_254) ) ;
    buf_clk cell_81 ( .C (clk), .D (signal_255), .Q (signal_256) ) ;
    buf_clk cell_83 ( .C (clk), .D (signal_257), .Q (signal_258) ) ;
    buf_clk cell_85 ( .C (clk), .D (signal_259), .Q (signal_260) ) ;
    buf_clk cell_87 ( .C (clk), .D (signal_261), .Q (signal_262) ) ;
    buf_clk cell_89 ( .C (clk), .D (signal_263), .Q (signal_264) ) ;
    buf_clk cell_91 ( .C (clk), .D (signal_265), .Q (signal_266) ) ;
    buf_clk cell_93 ( .C (clk), .D (signal_267), .Q (signal_268) ) ;
    buf_clk cell_95 ( .C (clk), .D (signal_269), .Q (signal_270) ) ;
    buf_clk cell_97 ( .C (clk), .D (signal_271), .Q (signal_272) ) ;
    buf_clk cell_99 ( .C (clk), .D (signal_273), .Q (signal_274) ) ;
    buf_clk cell_101 ( .C (clk), .D (signal_275), .Q (signal_276) ) ;
    buf_clk cell_103 ( .C (clk), .D (signal_277), .Q (signal_278) ) ;
    buf_clk cell_105 ( .C (clk), .D (signal_279), .Q (signal_280) ) ;
    buf_clk cell_107 ( .C (clk), .D (signal_281), .Q (signal_282) ) ;
    buf_clk cell_109 ( .C (clk), .D (signal_283), .Q (signal_284) ) ;
    buf_clk cell_121 ( .C (clk), .D (signal_295), .Q (signal_296) ) ;
    buf_clk cell_125 ( .C (clk), .D (signal_299), .Q (signal_300) ) ;
    buf_clk cell_129 ( .C (clk), .D (signal_303), .Q (signal_304) ) ;
    buf_clk cell_133 ( .C (clk), .D (signal_307), .Q (signal_308) ) ;
    buf_clk cell_137 ( .C (clk), .D (signal_311), .Q (signal_312) ) ;

    /* cells in depth 3 */
    buf_clk cell_110 ( .C (clk), .D (signal_41), .Q (signal_285) ) ;
    buf_clk cell_112 ( .C (clk), .D (signal_89), .Q (signal_287) ) ;
    buf_clk cell_114 ( .C (clk), .D (signal_90), .Q (signal_289) ) ;
    buf_clk cell_116 ( .C (clk), .D (signal_91), .Q (signal_291) ) ;
    buf_clk cell_118 ( .C (clk), .D (signal_92), .Q (signal_293) ) ;
    buf_clk cell_122 ( .C (clk), .D (signal_296), .Q (signal_297) ) ;
    buf_clk cell_126 ( .C (clk), .D (signal_300), .Q (signal_301) ) ;
    buf_clk cell_130 ( .C (clk), .D (signal_304), .Q (signal_305) ) ;
    buf_clk cell_134 ( .C (clk), .D (signal_308), .Q (signal_309) ) ;
    buf_clk cell_138 ( .C (clk), .D (signal_312), .Q (signal_313) ) ;
    buf_clk cell_140 ( .C (clk), .D (signal_51), .Q (signal_315) ) ;
    buf_clk cell_142 ( .C (clk), .D (signal_133), .Q (signal_317) ) ;
    buf_clk cell_144 ( .C (clk), .D (signal_134), .Q (signal_319) ) ;
    buf_clk cell_146 ( .C (clk), .D (signal_135), .Q (signal_321) ) ;
    buf_clk cell_148 ( .C (clk), .D (signal_136), .Q (signal_323) ) ;
    buf_clk cell_150 ( .C (clk), .D (signal_35), .Q (signal_325) ) ;
    buf_clk cell_152 ( .C (clk), .D (signal_149), .Q (signal_327) ) ;
    buf_clk cell_154 ( .C (clk), .D (signal_150), .Q (signal_329) ) ;
    buf_clk cell_156 ( .C (clk), .D (signal_151), .Q (signal_331) ) ;
    buf_clk cell_158 ( .C (clk), .D (signal_152), .Q (signal_333) ) ;
    buf_clk cell_160 ( .C (clk), .D (signal_36), .Q (signal_335) ) ;
    buf_clk cell_162 ( .C (clk), .D (signal_121), .Q (signal_337) ) ;
    buf_clk cell_164 ( .C (clk), .D (signal_122), .Q (signal_339) ) ;
    buf_clk cell_166 ( .C (clk), .D (signal_123), .Q (signal_341) ) ;
    buf_clk cell_168 ( .C (clk), .D (signal_124), .Q (signal_343) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_42 ( .a ({signal_274, signal_272, signal_270, signal_268, signal_266}), .b ({signal_128, signal_127, signal_126, signal_125, signal_49}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({signal_140, signal_139, signal_138, signal_137, signal_52}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_43 ( .a ({signal_284, signal_282, signal_280, signal_278, signal_276}), .b ({signal_132, signal_131, signal_130, signal_129, signal_50}), .clk (clk), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_144, signal_143, signal_142, signal_141, signal_53}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_46 ( .a ({signal_294, signal_292, signal_290, signal_288, signal_286}), .b ({signal_140, signal_139, signal_138, signal_137, signal_52}), .c ({signal_156, signal_155, signal_154, signal_153, signal_55}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_47 ( .a ({signal_314, signal_310, signal_306, signal_302, signal_298}), .b ({signal_140, signal_139, signal_138, signal_137, signal_52}), .c ({signal_160, signal_159, signal_158, signal_157, signal_56}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_48 ( .a ({signal_324, signal_322, signal_320, signal_318, signal_316}), .b ({signal_160, signal_159, signal_158, signal_157, signal_56}), .c ({signal_164, signal_163, signal_162, signal_161, signal_33}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_49 ( .a ({signal_144, signal_143, signal_142, signal_141, signal_53}), .b ({signal_156, signal_155, signal_154, signal_153, signal_55}), .c ({signal_168, signal_167, signal_166, signal_165, signal_34}) ) ;
    buf_clk cell_111 ( .C (clk), .D (signal_285), .Q (signal_286) ) ;
    buf_clk cell_113 ( .C (clk), .D (signal_287), .Q (signal_288) ) ;
    buf_clk cell_115 ( .C (clk), .D (signal_289), .Q (signal_290) ) ;
    buf_clk cell_117 ( .C (clk), .D (signal_291), .Q (signal_292) ) ;
    buf_clk cell_119 ( .C (clk), .D (signal_293), .Q (signal_294) ) ;
    buf_clk cell_123 ( .C (clk), .D (signal_297), .Q (signal_298) ) ;
    buf_clk cell_127 ( .C (clk), .D (signal_301), .Q (signal_302) ) ;
    buf_clk cell_131 ( .C (clk), .D (signal_305), .Q (signal_306) ) ;
    buf_clk cell_135 ( .C (clk), .D (signal_309), .Q (signal_310) ) ;
    buf_clk cell_139 ( .C (clk), .D (signal_313), .Q (signal_314) ) ;
    buf_clk cell_141 ( .C (clk), .D (signal_315), .Q (signal_316) ) ;
    buf_clk cell_143 ( .C (clk), .D (signal_317), .Q (signal_318) ) ;
    buf_clk cell_145 ( .C (clk), .D (signal_319), .Q (signal_320) ) ;
    buf_clk cell_147 ( .C (clk), .D (signal_321), .Q (signal_322) ) ;
    buf_clk cell_149 ( .C (clk), .D (signal_323), .Q (signal_324) ) ;
    buf_clk cell_151 ( .C (clk), .D (signal_325), .Q (signal_326) ) ;
    buf_clk cell_153 ( .C (clk), .D (signal_327), .Q (signal_328) ) ;
    buf_clk cell_155 ( .C (clk), .D (signal_329), .Q (signal_330) ) ;
    buf_clk cell_157 ( .C (clk), .D (signal_331), .Q (signal_332) ) ;
    buf_clk cell_159 ( .C (clk), .D (signal_333), .Q (signal_334) ) ;
    buf_clk cell_161 ( .C (clk), .D (signal_335), .Q (signal_336) ) ;
    buf_clk cell_163 ( .C (clk), .D (signal_337), .Q (signal_338) ) ;
    buf_clk cell_165 ( .C (clk), .D (signal_339), .Q (signal_340) ) ;
    buf_clk cell_167 ( .C (clk), .D (signal_341), .Q (signal_342) ) ;
    buf_clk cell_169 ( .C (clk), .D (signal_343), .Q (signal_344) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_334, signal_332, signal_330, signal_328, signal_326}), .Q ({Y_s4[3], Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_344, signal_342, signal_340, signal_338, signal_336}), .Q ({Y_s4[2], Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_164, signal_163, signal_162, signal_161, signal_33}), .Q ({Y_s4[1], Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_168, signal_167, signal_166, signal_165, signal_34}), .Q ({Y_s4[0], Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
