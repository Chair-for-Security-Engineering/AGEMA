/* modified netlist. Source: module Midori64 in file ../CaseStudies/12_Midori64_round_based_enc_dec/FPGA_based/Midori_synthesis.v */
/* clock gating is added to the circuit, the latency increased 1 time(s)  */

module Midori64_GHPCLL_ClockGating_d1 (clk, reset, enc_dec, input_0_s0, key_s0, key_s1, input_0_s1, Fresh, done, output_1_s0, output_1_s1, Synch);
    input clk ;
    input reset ;
    input enc_dec ;
    input [63:0] input_0_s0 ;
    input [127:0] key_s0 ;
    input [127:0] key_s1 ;
    input [63:0] input_0_s1 ;
    input [1023:0] Fresh ;
    output done ;
    output [63:0] output_1_s0 ;
    output [63:0] output_1_s1 ;
    output Synch ;
    wire \Midori/rounds/constant_MUX/Mram_roundConstant15 ;
    wire \Midori/rounds/constant_MUX/Mram_roundConstant11 ;
    wire \Midori/rounds/constant_MUX/Mram_roundConstant8 ;
    wire \Midori/rounds/constant_MUX/Mram_roundConstant7 ;
    wire \Midori/rounds/constant_MUX/Mram_roundConstant6 ;
    wire \Midori/rounds/constant_MUX/Mram_roundConstant5 ;
    wire \Midori/rounds/constant_MUX/Mram_roundConstant3 ;
    wire \Midori/rounds/constant_MUX/Mram_roundConstant2 ;
    wire \Midori/rounds/constant_MUX/Mram_roundConstant1 ;
    wire [60:0] \Midori/rounds/ProcessedKey ;
    wire [63:1] \Midori/rounds/SelectedKey ;
    wire \Midori/rounds/roundResult_Reg/GEN[0].SFF/Q_663 ;
    wire \Midori/rounds/roundResult_Reg/GEN[1].SFF/Q_664 ;
    wire \Midori/rounds/roundResult_Reg/GEN[2].SFF/Q_665 ;
    wire \Midori/rounds/roundResult_Reg/GEN[3].SFF/Q_666 ;
    wire \Midori/rounds/roundResult_Reg/GEN[4].SFF/Q_667 ;
    wire \Midori/rounds/roundResult_Reg/GEN[5].SFF/Q_668 ;
    wire \Midori/rounds/roundResult_Reg/GEN[6].SFF/Q_669 ;
    wire \Midori/rounds/roundResult_Reg/GEN[7].SFF/Q_670 ;
    wire \Midori/rounds/roundResult_Reg/GEN[8].SFF/Q_671 ;
    wire \Midori/rounds/roundResult_Reg/GEN[9].SFF/Q_672 ;
    wire \Midori/rounds/roundResult_Reg/GEN[10].SFF/Q_673 ;
    wire \Midori/rounds/roundResult_Reg/GEN[11].SFF/Q_674 ;
    wire \Midori/rounds/roundResult_Reg/GEN[12].SFF/Q_675 ;
    wire \Midori/rounds/roundResult_Reg/GEN[13].SFF/Q_676 ;
    wire \Midori/rounds/roundResult_Reg/GEN[14].SFF/Q_677 ;
    wire \Midori/rounds/roundResult_Reg/GEN[15].SFF/Q_678 ;
    wire \Midori/rounds/roundResult_Reg/GEN[16].SFF/Q_679 ;
    wire \Midori/rounds/roundResult_Reg/GEN[17].SFF/Q_680 ;
    wire \Midori/rounds/roundResult_Reg/GEN[18].SFF/Q_681 ;
    wire \Midori/rounds/roundResult_Reg/GEN[19].SFF/Q_682 ;
    wire \Midori/rounds/roundResult_Reg/GEN[20].SFF/Q_683 ;
    wire \Midori/rounds/roundResult_Reg/GEN[21].SFF/Q_684 ;
    wire \Midori/rounds/roundResult_Reg/GEN[22].SFF/Q_685 ;
    wire \Midori/rounds/roundResult_Reg/GEN[23].SFF/Q_686 ;
    wire \Midori/rounds/roundResult_Reg/GEN[24].SFF/Q_687 ;
    wire \Midori/rounds/roundResult_Reg/GEN[25].SFF/Q_688 ;
    wire \Midori/rounds/roundResult_Reg/GEN[26].SFF/Q_689 ;
    wire \Midori/rounds/roundResult_Reg/GEN[27].SFF/Q_690 ;
    wire \Midori/rounds/roundResult_Reg/GEN[28].SFF/Q_691 ;
    wire \Midori/rounds/roundResult_Reg/GEN[29].SFF/Q_692 ;
    wire \Midori/rounds/roundResult_Reg/GEN[30].SFF/Q_693 ;
    wire \Midori/rounds/roundResult_Reg/GEN[31].SFF/Q_694 ;
    wire \Midori/rounds/roundResult_Reg/GEN[32].SFF/Q_695 ;
    wire \Midori/rounds/roundResult_Reg/GEN[33].SFF/Q_696 ;
    wire \Midori/rounds/roundResult_Reg/GEN[34].SFF/Q_697 ;
    wire \Midori/rounds/roundResult_Reg/GEN[35].SFF/Q_698 ;
    wire \Midori/rounds/roundResult_Reg/GEN[36].SFF/Q_699 ;
    wire \Midori/rounds/roundResult_Reg/GEN[37].SFF/Q_700 ;
    wire \Midori/rounds/roundResult_Reg/GEN[38].SFF/Q_701 ;
    wire \Midori/rounds/roundResult_Reg/GEN[39].SFF/Q_702 ;
    wire \Midori/rounds/roundResult_Reg/GEN[40].SFF/Q_703 ;
    wire \Midori/rounds/roundResult_Reg/GEN[41].SFF/Q_704 ;
    wire \Midori/rounds/roundResult_Reg/GEN[42].SFF/Q_705 ;
    wire \Midori/rounds/roundResult_Reg/GEN[43].SFF/Q_706 ;
    wire \Midori/rounds/roundResult_Reg/GEN[44].SFF/Q_707 ;
    wire \Midori/rounds/roundResult_Reg/GEN[45].SFF/Q_708 ;
    wire \Midori/rounds/roundResult_Reg/GEN[46].SFF/Q_709 ;
    wire \Midori/rounds/roundResult_Reg/GEN[47].SFF/Q_710 ;
    wire \Midori/rounds/roundResult_Reg/GEN[48].SFF/Q_711 ;
    wire \Midori/rounds/roundResult_Reg/GEN[49].SFF/Q_712 ;
    wire \Midori/rounds/roundResult_Reg/GEN[50].SFF/Q_713 ;
    wire \Midori/rounds/roundResult_Reg/GEN[51].SFF/Q_714 ;
    wire \Midori/rounds/roundResult_Reg/GEN[52].SFF/Q_715 ;
    wire \Midori/rounds/roundResult_Reg/GEN[53].SFF/Q_716 ;
    wire \Midori/rounds/roundResult_Reg/GEN[54].SFF/Q_717 ;
    wire \Midori/rounds/roundResult_Reg/GEN[55].SFF/Q_718 ;
    wire \Midori/rounds/roundResult_Reg/GEN[56].SFF/Q_719 ;
    wire \Midori/rounds/roundResult_Reg/GEN[57].SFF/Q_720 ;
    wire \Midori/rounds/roundResult_Reg/GEN[58].SFF/Q_721 ;
    wire \Midori/rounds/roundResult_Reg/GEN[59].SFF/Q_722 ;
    wire \Midori/rounds/roundResult_Reg/GEN[60].SFF/Q_723 ;
    wire \Midori/rounds/roundResult_Reg/GEN[61].SFF/Q_724 ;
    wire \Midori/rounds/roundResult_Reg/GEN[62].SFF/Q_725 ;
    wire \Midori/rounds/roundResult_Reg/GEN[63].SFF/Q_726 ;
    wire \Midori/rounds/roundResult_Reg/GEN[0].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[1].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[2].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[3].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[4].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[5].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[6].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[7].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[8].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[9].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[10].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[11].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[12].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[13].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[14].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[15].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[16].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[17].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[18].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[19].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[20].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[21].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[22].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[23].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[24].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[25].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[26].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[27].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[28].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[29].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[30].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[31].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[32].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[33].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[34].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[35].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[36].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[37].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[38].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[39].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[40].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[41].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[42].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[43].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[44].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[45].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[46].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[47].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[48].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[49].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[50].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[51].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[52].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[53].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[54].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[55].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[56].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[57].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[58].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[59].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[60].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[61].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[62].SFF/DQ ;
    wire \Midori/rounds/roundResult_Reg/GEN[63].SFF/DQ ;
    wire \Midori/rounds/Mxor_ProcessedKey<36>_xo<0> ;
    wire \Midori/rounds/Mxor_ProcessedKey<52>_xo<0> ;
    wire \Midori/rounds/Mxor_ProcessedKey<48>_xo<0> ;
    wire N9 ;
    wire N111 ;
    wire N13 ;
    wire N15 ;
    wire N17 ;
    wire N19 ;
    wire N21 ;
    wire N23 ;
    wire N25 ;
    wire N27 ;
    wire N29 ;
    wire N34 ;
    wire \controller/roundCounter/count_3_1_1066 ;
    wire \controller/roundCounter/count_2_1_1067 ;
    wire \controller/roundCounter/count_0_1_1068 ;
    wire \controller/roundCounter/count_1_1_1069 ;
    wire \controller/roundCounter/count_2_2_1070 ;
    wire \controller/roundCounter/count_3_2_1071 ;
    wire \controller/roundCounter/count_1_2_1072 ;
    wire N36 ;
    wire N37 ;
    wire N38 ;
    wire N39 ;
    wire N40 ;
    wire N41 ;
    wire [63:0] \Midori/add_Result_Start ;
    wire [63:0] \Midori/rounds_Output ;
    wire [3:0] Result ;
    wire [3:0] \controller/roundCounter/count ;
    wire [63:0] \Midori/rounds/mul_Result ;
    wire [63:0] \Midori/rounds/mul_ResultXORkey ;
    wire [63:0] \Midori/rounds/mul_input ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire clk_gated ;

    /* cells in depth 0 */
    LUT4 #( .INIT ( 16'h8000 ) ) \controller/done<3>1 ( .I0 (\controller/roundCounter/count [3]), .I1 (\controller/roundCounter/count [2]), .I2 (\controller/roundCounter/count [1]), .I3 (\controller/roundCounter/count [0]), .O (done) ) ;
    LUT2 #( .INIT ( 4'h6 ) ) \controller/roundCounter/Mcount_count_xor<1>11 ( .I0 (\controller/roundCounter/count [1]), .I1 (\controller/roundCounter/count [0]), .O (Result[1]) ) ;
    LUT4 #( .INIT ( 16'h6CCC ) ) \Result<3>1 ( .I0 (\controller/roundCounter/count [2]), .I1 (\controller/roundCounter/count [3]), .I2 (\controller/roundCounter/count [0]), .I3 (\controller/roundCounter/count [1]), .O (Result[3]) ) ;
    LUT3 #( .INIT ( 8'h6A ) ) \Result<2>1 ( .I0 (\controller/roundCounter/count [2]), .I1 (\controller/roundCounter/count [0]), .I2 (\controller/roundCounter/count [1]), .O (Result[2]) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<9>1 ( .I0 ({key_s1[73], key_s0[73]}), .I1 ({input_0_s1[9], input_0_s0[9]}), .I2 ({key_s1[9], key_s0[9]}), .O ({new_AGEMA_signal_1214, \Midori/add_Result_Start [9]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<8>1 ( .I0 ({key_s1[72], key_s0[72]}), .I1 ({input_0_s1[8], input_0_s0[8]}), .I2 ({key_s1[8], key_s0[8]}), .O ({new_AGEMA_signal_1218, \Midori/add_Result_Start [8]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<7>1 ( .I0 ({key_s1[71], key_s0[71]}), .I1 ({input_0_s1[7], input_0_s0[7]}), .I2 ({key_s1[7], key_s0[7]}), .O ({new_AGEMA_signal_1222, \Midori/add_Result_Start [7]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<63>1 ( .I0 ({input_0_s1[63], input_0_s0[63]}), .I1 ({key_s1[63], key_s0[63]}), .I2 ({key_s1[127], key_s0[127]}), .O ({new_AGEMA_signal_1226, \Midori/add_Result_Start [63]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<62>1 ( .I0 ({input_0_s1[62], input_0_s0[62]}), .I1 ({key_s1[62], key_s0[62]}), .I2 ({key_s1[126], key_s0[126]}), .O ({new_AGEMA_signal_1230, \Midori/add_Result_Start [62]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<61>1 ( .I0 ({input_0_s1[61], input_0_s0[61]}), .I1 ({key_s1[61], key_s0[61]}), .I2 ({key_s1[125], key_s0[125]}), .O ({new_AGEMA_signal_1234, \Midori/add_Result_Start [61]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<60>1 ( .I0 ({input_0_s1[60], input_0_s0[60]}), .I1 ({key_s1[60], key_s0[60]}), .I2 ({key_s1[124], key_s0[124]}), .O ({new_AGEMA_signal_1238, \Midori/add_Result_Start [60]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<6>1 ( .I0 ({key_s1[70], key_s0[70]}), .I1 ({input_0_s1[6], input_0_s0[6]}), .I2 ({key_s1[6], key_s0[6]}), .O ({new_AGEMA_signal_1242, \Midori/add_Result_Start [6]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<59>1 ( .I0 ({key_s1[123], key_s0[123]}), .I1 ({input_0_s1[59], input_0_s0[59]}), .I2 ({key_s1[59], key_s0[59]}), .O ({new_AGEMA_signal_1246, \Midori/add_Result_Start [59]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<58>1 ( .I0 ({key_s1[122], key_s0[122]}), .I1 ({input_0_s1[58], input_0_s0[58]}), .I2 ({key_s1[58], key_s0[58]}), .O ({new_AGEMA_signal_1250, \Midori/add_Result_Start [58]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<57>1 ( .I0 ({key_s1[121], key_s0[121]}), .I1 ({input_0_s1[57], input_0_s0[57]}), .I2 ({key_s1[57], key_s0[57]}), .O ({new_AGEMA_signal_1254, \Midori/add_Result_Start [57]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<56>1 ( .I0 ({key_s1[120], key_s0[120]}), .I1 ({input_0_s1[56], input_0_s0[56]}), .I2 ({key_s1[56], key_s0[56]}), .O ({new_AGEMA_signal_1258, \Midori/add_Result_Start [56]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<55>1 ( .I0 ({input_0_s1[55], input_0_s0[55]}), .I1 ({key_s1[55], key_s0[55]}), .I2 ({key_s1[119], key_s0[119]}), .O ({new_AGEMA_signal_1262, \Midori/add_Result_Start [55]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<54>1 ( .I0 ({input_0_s1[54], input_0_s0[54]}), .I1 ({key_s1[54], key_s0[54]}), .I2 ({key_s1[118], key_s0[118]}), .O ({new_AGEMA_signal_1266, \Midori/add_Result_Start [54]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<53>1 ( .I0 ({input_0_s1[53], input_0_s0[53]}), .I1 ({key_s1[53], key_s0[53]}), .I2 ({key_s1[117], key_s0[117]}), .O ({new_AGEMA_signal_1270, \Midori/add_Result_Start [53]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<52>1 ( .I0 ({input_0_s1[52], input_0_s0[52]}), .I1 ({key_s1[52], key_s0[52]}), .I2 ({key_s1[116], key_s0[116]}), .O ({new_AGEMA_signal_1274, \Midori/add_Result_Start [52]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<51>1 ( .I0 ({input_0_s1[51], input_0_s0[51]}), .I1 ({key_s1[51], key_s0[51]}), .I2 ({key_s1[115], key_s0[115]}), .O ({new_AGEMA_signal_1278, \Midori/add_Result_Start [51]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<50>1 ( .I0 ({input_0_s1[50], input_0_s0[50]}), .I1 ({key_s1[50], key_s0[50]}), .I2 ({key_s1[114], key_s0[114]}), .O ({new_AGEMA_signal_1282, \Midori/add_Result_Start [50]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<5>1 ( .I0 ({input_0_s1[5], input_0_s0[5]}), .I1 ({key_s1[5], key_s0[5]}), .I2 ({key_s1[69], key_s0[69]}), .O ({new_AGEMA_signal_1286, \Midori/add_Result_Start [5]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<49>1 ( .I0 ({key_s1[113], key_s0[113]}), .I1 ({input_0_s1[49], input_0_s0[49]}), .I2 ({key_s1[49], key_s0[49]}), .O ({new_AGEMA_signal_1290, \Midori/add_Result_Start [49]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<48>1 ( .I0 ({key_s1[112], key_s0[112]}), .I1 ({input_0_s1[48], input_0_s0[48]}), .I2 ({key_s1[48], key_s0[48]}), .O ({new_AGEMA_signal_1294, \Midori/add_Result_Start [48]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<47>1 ( .I0 ({key_s1[111], key_s0[111]}), .I1 ({input_0_s1[47], input_0_s0[47]}), .I2 ({key_s1[47], key_s0[47]}), .O ({new_AGEMA_signal_1298, \Midori/add_Result_Start [47]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<46>1 ( .I0 ({key_s1[110], key_s0[110]}), .I1 ({input_0_s1[46], input_0_s0[46]}), .I2 ({key_s1[46], key_s0[46]}), .O ({new_AGEMA_signal_1302, \Midori/add_Result_Start [46]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<45>1 ( .I0 ({input_0_s1[45], input_0_s0[45]}), .I1 ({key_s1[45], key_s0[45]}), .I2 ({key_s1[109], key_s0[109]}), .O ({new_AGEMA_signal_1306, \Midori/add_Result_Start [45]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<44>1 ( .I0 ({input_0_s1[44], input_0_s0[44]}), .I1 ({key_s1[44], key_s0[44]}), .I2 ({key_s1[108], key_s0[108]}), .O ({new_AGEMA_signal_1310, \Midori/add_Result_Start [44]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<43>1 ( .I0 ({input_0_s1[43], input_0_s0[43]}), .I1 ({key_s1[43], key_s0[43]}), .I2 ({key_s1[107], key_s0[107]}), .O ({new_AGEMA_signal_1314, \Midori/add_Result_Start [43]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<42>1 ( .I0 ({input_0_s1[42], input_0_s0[42]}), .I1 ({key_s1[42], key_s0[42]}), .I2 ({key_s1[106], key_s0[106]}), .O ({new_AGEMA_signal_1318, \Midori/add_Result_Start [42]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<41>1 ( .I0 ({input_0_s1[41], input_0_s0[41]}), .I1 ({key_s1[41], key_s0[41]}), .I2 ({key_s1[105], key_s0[105]}), .O ({new_AGEMA_signal_1322, \Midori/add_Result_Start [41]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<40>1 ( .I0 ({input_0_s1[40], input_0_s0[40]}), .I1 ({key_s1[40], key_s0[40]}), .I2 ({key_s1[104], key_s0[104]}), .O ({new_AGEMA_signal_1326, \Midori/add_Result_Start [40]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<4>1 ( .I0 ({input_0_s1[4], input_0_s0[4]}), .I1 ({key_s1[4], key_s0[4]}), .I2 ({key_s1[68], key_s0[68]}), .O ({new_AGEMA_signal_1330, \Midori/add_Result_Start [4]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<39>1 ( .I0 ({key_s1[103], key_s0[103]}), .I1 ({input_0_s1[39], input_0_s0[39]}), .I2 ({key_s1[39], key_s0[39]}), .O ({new_AGEMA_signal_1334, \Midori/add_Result_Start [39]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<38>1 ( .I0 ({key_s1[102], key_s0[102]}), .I1 ({input_0_s1[38], input_0_s0[38]}), .I2 ({key_s1[38], key_s0[38]}), .O ({new_AGEMA_signal_1338, \Midori/add_Result_Start [38]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<37>1 ( .I0 ({key_s1[101], key_s0[101]}), .I1 ({input_0_s1[37], input_0_s0[37]}), .I2 ({key_s1[37], key_s0[37]}), .O ({new_AGEMA_signal_1342, \Midori/add_Result_Start [37]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<36>1 ( .I0 ({key_s1[100], key_s0[100]}), .I1 ({input_0_s1[36], input_0_s0[36]}), .I2 ({key_s1[36], key_s0[36]}), .O ({new_AGEMA_signal_1346, \Midori/add_Result_Start [36]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<35>1 ( .I0 ({input_0_s1[35], input_0_s0[35]}), .I1 ({key_s1[35], key_s0[35]}), .I2 ({key_s1[99], key_s0[99]}), .O ({new_AGEMA_signal_1350, \Midori/add_Result_Start [35]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<34>1 ( .I0 ({input_0_s1[34], input_0_s0[34]}), .I1 ({key_s1[34], key_s0[34]}), .I2 ({key_s1[98], key_s0[98]}), .O ({new_AGEMA_signal_1354, \Midori/add_Result_Start [34]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<33>1 ( .I0 ({input_0_s1[33], input_0_s0[33]}), .I1 ({key_s1[33], key_s0[33]}), .I2 ({key_s1[97], key_s0[97]}), .O ({new_AGEMA_signal_1358, \Midori/add_Result_Start [33]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<32>1 ( .I0 ({input_0_s1[32], input_0_s0[32]}), .I1 ({key_s1[32], key_s0[32]}), .I2 ({key_s1[96], key_s0[96]}), .O ({new_AGEMA_signal_1362, \Midori/add_Result_Start [32]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<31>1 ( .I0 ({input_0_s1[31], input_0_s0[31]}), .I1 ({key_s1[31], key_s0[31]}), .I2 ({key_s1[95], key_s0[95]}), .O ({new_AGEMA_signal_1366, \Midori/add_Result_Start [31]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<30>1 ( .I0 ({input_0_s1[30], input_0_s0[30]}), .I1 ({key_s1[30], key_s0[30]}), .I2 ({key_s1[94], key_s0[94]}), .O ({new_AGEMA_signal_1370, \Midori/add_Result_Start [30]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<3>1 ( .I0 ({input_0_s1[3], input_0_s0[3]}), .I1 ({key_s1[3], key_s0[3]}), .I2 ({key_s1[67], key_s0[67]}), .O ({new_AGEMA_signal_1374, \Midori/add_Result_Start [3]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<29>1 ( .I0 ({key_s1[93], key_s0[93]}), .I1 ({input_0_s1[29], input_0_s0[29]}), .I2 ({key_s1[29], key_s0[29]}), .O ({new_AGEMA_signal_1378, \Midori/add_Result_Start [29]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<28>1 ( .I0 ({key_s1[92], key_s0[92]}), .I1 ({input_0_s1[28], input_0_s0[28]}), .I2 ({key_s1[28], key_s0[28]}), .O ({new_AGEMA_signal_1382, \Midori/add_Result_Start [28]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<27>1 ( .I0 ({key_s1[91], key_s0[91]}), .I1 ({input_0_s1[27], input_0_s0[27]}), .I2 ({key_s1[27], key_s0[27]}), .O ({new_AGEMA_signal_1386, \Midori/add_Result_Start [27]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<26>1 ( .I0 ({key_s1[90], key_s0[90]}), .I1 ({input_0_s1[26], input_0_s0[26]}), .I2 ({key_s1[26], key_s0[26]}), .O ({new_AGEMA_signal_1390, \Midori/add_Result_Start [26]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<25>1 ( .I0 ({input_0_s1[25], input_0_s0[25]}), .I1 ({key_s1[25], key_s0[25]}), .I2 ({key_s1[89], key_s0[89]}), .O ({new_AGEMA_signal_1394, \Midori/add_Result_Start [25]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<24>1 ( .I0 ({input_0_s1[24], input_0_s0[24]}), .I1 ({key_s1[24], key_s0[24]}), .I2 ({key_s1[88], key_s0[88]}), .O ({new_AGEMA_signal_1398, \Midori/add_Result_Start [24]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<23>1 ( .I0 ({input_0_s1[23], input_0_s0[23]}), .I1 ({key_s1[23], key_s0[23]}), .I2 ({key_s1[87], key_s0[87]}), .O ({new_AGEMA_signal_1402, \Midori/add_Result_Start [23]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<22>1 ( .I0 ({input_0_s1[22], input_0_s0[22]}), .I1 ({key_s1[22], key_s0[22]}), .I2 ({key_s1[86], key_s0[86]}), .O ({new_AGEMA_signal_1406, \Midori/add_Result_Start [22]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<21>1 ( .I0 ({input_0_s1[21], input_0_s0[21]}), .I1 ({key_s1[21], key_s0[21]}), .I2 ({key_s1[85], key_s0[85]}), .O ({new_AGEMA_signal_1410, \Midori/add_Result_Start [21]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<20>1 ( .I0 ({input_0_s1[20], input_0_s0[20]}), .I1 ({key_s1[20], key_s0[20]}), .I2 ({key_s1[84], key_s0[84]}), .O ({new_AGEMA_signal_1414, \Midori/add_Result_Start [20]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<2>1 ( .I0 ({input_0_s1[2], input_0_s0[2]}), .I1 ({key_s1[2], key_s0[2]}), .I2 ({key_s1[66], key_s0[66]}), .O ({new_AGEMA_signal_1418, \Midori/add_Result_Start [2]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<19>1 ( .I0 ({key_s1[83], key_s0[83]}), .I1 ({input_0_s1[19], input_0_s0[19]}), .I2 ({key_s1[19], key_s0[19]}), .O ({new_AGEMA_signal_1422, \Midori/add_Result_Start [19]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<18>1 ( .I0 ({key_s1[82], key_s0[82]}), .I1 ({input_0_s1[18], input_0_s0[18]}), .I2 ({key_s1[18], key_s0[18]}), .O ({new_AGEMA_signal_1426, \Midori/add_Result_Start [18]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<17>1 ( .I0 ({key_s1[81], key_s0[81]}), .I1 ({input_0_s1[17], input_0_s0[17]}), .I2 ({key_s1[17], key_s0[17]}), .O ({new_AGEMA_signal_1430, \Midori/add_Result_Start [17]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<16>1 ( .I0 ({key_s1[80], key_s0[80]}), .I1 ({input_0_s1[16], input_0_s0[16]}), .I2 ({key_s1[16], key_s0[16]}), .O ({new_AGEMA_signal_1434, \Midori/add_Result_Start [16]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<15>1 ( .I0 ({input_0_s1[15], input_0_s0[15]}), .I1 ({key_s1[15], key_s0[15]}), .I2 ({key_s1[79], key_s0[79]}), .O ({new_AGEMA_signal_1438, \Midori/add_Result_Start [15]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<14>1 ( .I0 ({input_0_s1[14], input_0_s0[14]}), .I1 ({key_s1[14], key_s0[14]}), .I2 ({key_s1[78], key_s0[78]}), .O ({new_AGEMA_signal_1442, \Midori/add_Result_Start [14]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<13>1 ( .I0 ({input_0_s1[13], input_0_s0[13]}), .I1 ({key_s1[13], key_s0[13]}), .I2 ({key_s1[77], key_s0[77]}), .O ({new_AGEMA_signal_1446, \Midori/add_Result_Start [13]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<12>1 ( .I0 ({input_0_s1[12], input_0_s0[12]}), .I1 ({key_s1[12], key_s0[12]}), .I2 ({key_s1[76], key_s0[76]}), .O ({new_AGEMA_signal_1450, \Midori/add_Result_Start [12]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<11>1 ( .I0 ({input_0_s1[11], input_0_s0[11]}), .I1 ({key_s1[11], key_s0[11]}), .I2 ({key_s1[75], key_s0[75]}), .O ({new_AGEMA_signal_1454, \Midori/add_Result_Start [11]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<10>1 ( .I0 ({input_0_s1[10], input_0_s0[10]}), .I1 ({key_s1[10], key_s0[10]}), .I2 ({key_s1[74], key_s0[74]}), .O ({new_AGEMA_signal_1458, \Midori/add_Result_Start [10]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<1>1 ( .I0 ({input_0_s1[1], input_0_s0[1]}), .I1 ({key_s1[1], key_s0[1]}), .I2 ({key_s1[65], key_s0[65]}), .O ({new_AGEMA_signal_1462, \Midori/add_Result_Start [1]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \Midori/add_Result_Start<0>1 ( .I0 ({input_0_s1[0], input_0_s0[0]}), .I1 ({key_s1[0], key_s0[0]}), .I2 ({key_s1[64], key_s0[64]}), .O ({new_AGEMA_signal_1466, \Midori/add_Result_Start [0]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h53AC ) , .MASK ( 4'b1100 ), .INIT2 ( 16'hACAC ) ) \Midori/rounds/Mxor_ProcessedKey<8>_xo<0>1 ( .I0 ({key_s1[8], key_s0[8]}), .I1 ({key_s1[72], key_s0[72]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .I3 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant2 }), .O ({new_AGEMA_signal_1600, \Midori/rounds/ProcessedKey [8]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h53AC ) , .MASK ( 4'b1100 ), .INIT2 ( 16'hACAC ) ) \Midori/rounds/Mxor_ProcessedKey<60>_xo<0>1 ( .I0 ({key_s1[60], key_s0[60]}), .I1 ({key_s1[124], key_s0[124]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .I3 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant15 }), .O ({new_AGEMA_signal_1601, \Midori/rounds/ProcessedKey [60]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h53AC ) , .MASK ( 4'b1100 ), .INIT2 ( 16'hACAC ) ) \Midori/rounds/Mxor_ProcessedKey<4>_xo<0>1 ( .I0 ({key_s1[4], key_s0[4]}), .I1 ({key_s1[68], key_s0[68]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .I3 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant1 }), .O ({new_AGEMA_signal_1602, \Midori/rounds/ProcessedKey [4]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h53AC ) , .MASK ( 4'b1100 ), .INIT2 ( 16'hACAC ) ) \Midori/rounds/Mxor_ProcessedKey<44>_xo<0>1 ( .I0 ({key_s1[44], key_s0[44]}), .I1 ({key_s1[108], key_s0[108]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .I3 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant11 }), .O ({new_AGEMA_signal_1603, \Midori/rounds/ProcessedKey [44]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h53AC ) , .MASK ( 4'b1100 ), .INIT2 ( 16'hACAC ) ) \Midori/rounds/Mxor_ProcessedKey<32>_xo<0>1 ( .I0 ({key_s1[32], key_s0[32]}), .I1 ({key_s1[96], key_s0[96]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .I3 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant8 }), .O ({new_AGEMA_signal_1604, \Midori/rounds/ProcessedKey [32]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h53AC ) , .MASK ( 4'b1100 ), .INIT2 ( 16'hACAC ) ) \Midori/rounds/Mxor_ProcessedKey<28>_xo<0>1 ( .I0 ({key_s1[28], key_s0[28]}), .I1 ({key_s1[92], key_s0[92]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .I3 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant7 }), .O ({new_AGEMA_signal_1605, \Midori/rounds/ProcessedKey [28]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h53AC ) , .MASK ( 4'b1100 ), .INIT2 ( 16'hACAC ) ) \Midori/rounds/Mxor_ProcessedKey<24>_xo<0>1 ( .I0 ({key_s1[24], key_s0[24]}), .I1 ({key_s1[88], key_s0[88]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .I3 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant6 }), .O ({new_AGEMA_signal_1606, \Midori/rounds/ProcessedKey [24]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h53AC ) , .MASK ( 4'b1100 ), .INIT2 ( 16'hACAC ) ) \Midori/rounds/Mxor_ProcessedKey<20>_xo<0>1 ( .I0 ({key_s1[20], key_s0[20]}), .I1 ({key_s1[84], key_s0[84]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .I3 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant5 }), .O ({new_AGEMA_signal_1607, \Midori/rounds/ProcessedKey [20]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h53AC ) , .MASK ( 4'b1100 ), .INIT2 ( 16'hACAC ) ) \Midori/rounds/Mxor_ProcessedKey<12>_xo<0>1 ( .I0 ({key_s1[12], key_s0[12]}), .I1 ({key_s1[76], key_s0[76]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .I3 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant3 }), .O ({new_AGEMA_signal_1608, \Midori/rounds/ProcessedKey [12]}) ) ;
    LUT5 #( .INIT ( 32'h30C34002 ) ) \Midori/rounds/constant_MUX/Mram_roundConstant1111 ( .I0 (enc_dec), .I1 (\controller/roundCounter/count [3]), .I2 (\controller/roundCounter/count [2]), .I3 (\controller/roundCounter/count [1]), .I4 (\controller/roundCounter/count [0]), .O (\Midori/rounds/constant_MUX/Mram_roundConstant11 ) ) ;
    LUT5 #( .INIT ( 32'h005A6186 ) ) \Midori/rounds/constant_MUX/Mram_roundConstant151 ( .I0 (enc_dec), .I1 (\controller/roundCounter/count [3]), .I2 (\controller/roundCounter/count [2]), .I3 (\controller/roundCounter/count [1]), .I4 (\controller/roundCounter/count [0]), .O (\Midori/rounds/constant_MUX/Mram_roundConstant15 ) ) ;
    LUT5 #( .INIT ( 32'h30DB1818 ) ) \Midori/rounds/constant_MUX/Mram_roundConstant61 ( .I0 (enc_dec), .I1 (\controller/roundCounter/count [3]), .I2 (\controller/roundCounter/count [2]), .I3 (\controller/roundCounter/count [1]), .I4 (\controller/roundCounter/count [0]), .O (\Midori/rounds/constant_MUX/Mram_roundConstant6 ) ) ;
    LUT5 #( .INIT ( 32'h003C93C9 ) ) \Midori/rounds/constant_MUX/Mram_roundConstant51 ( .I0 (enc_dec), .I1 (\controller/roundCounter/count [3]), .I2 (\controller/roundCounter/count [2]), .I3 (\controller/roundCounter/count [1]), .I4 (\controller/roundCounter/count [0]), .O (\Midori/rounds/constant_MUX/Mram_roundConstant5 ) ) ;
    LUT5 #( .INIT ( 32'h0F429C39 ) ) \Midori/rounds/constant_MUX/Mram_roundConstant111 ( .I0 (enc_dec), .I1 (\controller/roundCounter/count [3]), .I2 (\controller/roundCounter/count [2]), .I3 (\controller/roundCounter/count [1]), .I4 (\controller/roundCounter/count [0]), .O (\Midori/rounds/constant_MUX/Mram_roundConstant1 ) ) ;
    LUT5 #( .INIT ( 32'h3018C663 ) ) \Midori/rounds/constant_MUX/Mram_roundConstant81 ( .I0 (enc_dec), .I1 (\controller/roundCounter/count [3]), .I2 (\controller/roundCounter/count [2]), .I3 (\controller/roundCounter/count [1]), .I4 (\controller/roundCounter/count [0]), .O (\Midori/rounds/constant_MUX/Mram_roundConstant8 ) ) ;
    LUT5 #( .INIT ( 32'h0C4827E4 ) ) \Midori/rounds/constant_MUX/Mram_roundConstant21 ( .I0 (enc_dec), .I1 (\controller/roundCounter/count [1]), .I2 (\controller/roundCounter/count [3]), .I3 (\controller/roundCounter/count [2]), .I4 (\controller/roundCounter/count [0]), .O (\Midori/rounds/constant_MUX/Mram_roundConstant2 ) ) ;
    LUT5 #( .INIT ( 32'h36E7E427 ) ) \Midori/rounds/constant_MUX/Mram_roundConstant71 ( .I0 (enc_dec), .I1 (\controller/roundCounter/count [3]), .I2 (\controller/roundCounter/count [2]), .I3 (\controller/roundCounter/count [1]), .I4 (\controller/roundCounter/count [0]), .O (\Midori/rounds/constant_MUX/Mram_roundConstant7 ) ) ;
    LUT5 #( .INIT ( 32'h36660810 ) ) \Midori/rounds/constant_MUX/Mram_roundConstant31 ( .I0 (enc_dec), .I1 (\controller/roundCounter/count [3]), .I2 (\controller/roundCounter/count [2]), .I3 (\controller/roundCounter/count [1]), .I4 (\controller/roundCounter/count [0]), .O (\Midori/rounds/constant_MUX/Mram_roundConstant3 ) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[63].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[127], key_s0[127]}), .I2 ({key_s1[63], key_s0[63]}), .O ({new_AGEMA_signal_1467, \Midori/rounds/SelectedKey [63]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[62].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[126], key_s0[126]}), .I2 ({key_s1[62], key_s0[62]}), .O ({new_AGEMA_signal_1468, \Midori/rounds/SelectedKey [62]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[61].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[125], key_s0[125]}), .I2 ({key_s1[61], key_s0[61]}), .O ({new_AGEMA_signal_1469, \Midori/rounds/SelectedKey [61]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[59].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[123], key_s0[123]}), .I2 ({key_s1[59], key_s0[59]}), .O ({new_AGEMA_signal_1470, \Midori/rounds/SelectedKey [59]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[58].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[122], key_s0[122]}), .I2 ({key_s1[58], key_s0[58]}), .O ({new_AGEMA_signal_1471, \Midori/rounds/SelectedKey [58]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[57].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[121], key_s0[121]}), .I2 ({key_s1[57], key_s0[57]}), .O ({new_AGEMA_signal_1472, \Midori/rounds/SelectedKey [57]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[55].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[119], key_s0[119]}), .I2 ({key_s1[55], key_s0[55]}), .O ({new_AGEMA_signal_1473, \Midori/rounds/SelectedKey [55]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[54].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[118], key_s0[118]}), .I2 ({key_s1[54], key_s0[54]}), .O ({new_AGEMA_signal_1474, \Midori/rounds/SelectedKey [54]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[53].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[117], key_s0[117]}), .I2 ({key_s1[53], key_s0[53]}), .O ({new_AGEMA_signal_1475, \Midori/rounds/SelectedKey [53]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[51].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[115], key_s0[115]}), .I2 ({key_s1[51], key_s0[51]}), .O ({new_AGEMA_signal_1476, \Midori/rounds/SelectedKey [51]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[50].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[114], key_s0[114]}), .I2 ({key_s1[50], key_s0[50]}), .O ({new_AGEMA_signal_1477, \Midori/rounds/SelectedKey [50]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[49].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[113], key_s0[113]}), .I2 ({key_s1[49], key_s0[49]}), .O ({new_AGEMA_signal_1478, \Midori/rounds/SelectedKey [49]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[47].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[111], key_s0[111]}), .I2 ({key_s1[47], key_s0[47]}), .O ({new_AGEMA_signal_1479, \Midori/rounds/SelectedKey [47]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[46].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[110], key_s0[110]}), .I2 ({key_s1[46], key_s0[46]}), .O ({new_AGEMA_signal_1480, \Midori/rounds/SelectedKey [46]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[45].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[109], key_s0[109]}), .I2 ({key_s1[45], key_s0[45]}), .O ({new_AGEMA_signal_1481, \Midori/rounds/SelectedKey [45]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[43].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[107], key_s0[107]}), .I2 ({key_s1[43], key_s0[43]}), .O ({new_AGEMA_signal_1482, \Midori/rounds/SelectedKey [43]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[42].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[106], key_s0[106]}), .I2 ({key_s1[42], key_s0[42]}), .O ({new_AGEMA_signal_1483, \Midori/rounds/SelectedKey [42]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[41].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[105], key_s0[105]}), .I2 ({key_s1[41], key_s0[41]}), .O ({new_AGEMA_signal_1484, \Midori/rounds/SelectedKey [41]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[39].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[103], key_s0[103]}), .I2 ({key_s1[39], key_s0[39]}), .O ({new_AGEMA_signal_1485, \Midori/rounds/SelectedKey [39]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[38].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[102], key_s0[102]}), .I2 ({key_s1[38], key_s0[38]}), .O ({new_AGEMA_signal_1486, \Midori/rounds/SelectedKey [38]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[37].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[101], key_s0[101]}), .I2 ({key_s1[37], key_s0[37]}), .O ({new_AGEMA_signal_1487, \Midori/rounds/SelectedKey [37]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[35].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[99], key_s0[99]}), .I2 ({key_s1[35], key_s0[35]}), .O ({new_AGEMA_signal_1488, \Midori/rounds/SelectedKey [35]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[34].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[98], key_s0[98]}), .I2 ({key_s1[34], key_s0[34]}), .O ({new_AGEMA_signal_1489, \Midori/rounds/SelectedKey [34]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[33].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[97], key_s0[97]}), .I2 ({key_s1[33], key_s0[33]}), .O ({new_AGEMA_signal_1490, \Midori/rounds/SelectedKey [33]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[31].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[95], key_s0[95]}), .I2 ({key_s1[31], key_s0[31]}), .O ({new_AGEMA_signal_1491, \Midori/rounds/SelectedKey [31]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[30].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[94], key_s0[94]}), .I2 ({key_s1[30], key_s0[30]}), .O ({new_AGEMA_signal_1492, \Midori/rounds/SelectedKey [30]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[29].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[93], key_s0[93]}), .I2 ({key_s1[29], key_s0[29]}), .O ({new_AGEMA_signal_1493, \Midori/rounds/SelectedKey [29]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[27].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[91], key_s0[91]}), .I2 ({key_s1[27], key_s0[27]}), .O ({new_AGEMA_signal_1494, \Midori/rounds/SelectedKey [27]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[26].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[90], key_s0[90]}), .I2 ({key_s1[26], key_s0[26]}), .O ({new_AGEMA_signal_1495, \Midori/rounds/SelectedKey [26]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[25].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[89], key_s0[89]}), .I2 ({key_s1[25], key_s0[25]}), .O ({new_AGEMA_signal_1496, \Midori/rounds/SelectedKey [25]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[23].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[87], key_s0[87]}), .I2 ({key_s1[23], key_s0[23]}), .O ({new_AGEMA_signal_1497, \Midori/rounds/SelectedKey [23]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[22].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[86], key_s0[86]}), .I2 ({key_s1[22], key_s0[22]}), .O ({new_AGEMA_signal_1498, \Midori/rounds/SelectedKey [22]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[21].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[85], key_s0[85]}), .I2 ({key_s1[21], key_s0[21]}), .O ({new_AGEMA_signal_1499, \Midori/rounds/SelectedKey [21]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[19].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[83], key_s0[83]}), .I2 ({key_s1[19], key_s0[19]}), .O ({new_AGEMA_signal_1500, \Midori/rounds/SelectedKey [19]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[18].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[82], key_s0[82]}), .I2 ({key_s1[18], key_s0[18]}), .O ({new_AGEMA_signal_1501, \Midori/rounds/SelectedKey [18]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[17].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[81], key_s0[81]}), .I2 ({key_s1[17], key_s0[17]}), .O ({new_AGEMA_signal_1502, \Midori/rounds/SelectedKey [17]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[15].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[79], key_s0[79]}), .I2 ({key_s1[15], key_s0[15]}), .O ({new_AGEMA_signal_1503, \Midori/rounds/SelectedKey [15]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[14].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[78], key_s0[78]}), .I2 ({key_s1[14], key_s0[14]}), .O ({new_AGEMA_signal_1504, \Midori/rounds/SelectedKey [14]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[13].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[77], key_s0[77]}), .I2 ({key_s1[13], key_s0[13]}), .O ({new_AGEMA_signal_1505, \Midori/rounds/SelectedKey [13]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[11].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[75], key_s0[75]}), .I2 ({key_s1[11], key_s0[11]}), .O ({new_AGEMA_signal_1506, \Midori/rounds/SelectedKey [11]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[10].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[74], key_s0[74]}), .I2 ({key_s1[10], key_s0[10]}), .O ({new_AGEMA_signal_1507, \Midori/rounds/SelectedKey [10]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[9].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[73], key_s0[73]}), .I2 ({key_s1[9], key_s0[9]}), .O ({new_AGEMA_signal_1508, \Midori/rounds/SelectedKey [9]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[7].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[71], key_s0[71]}), .I2 ({key_s1[7], key_s0[7]}), .O ({new_AGEMA_signal_1509, \Midori/rounds/SelectedKey [7]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[6].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[70], key_s0[70]}), .I2 ({key_s1[6], key_s0[6]}), .O ({new_AGEMA_signal_1510, \Midori/rounds/SelectedKey [6]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[5].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[69], key_s0[69]}), .I2 ({key_s1[5], key_s0[5]}), .O ({new_AGEMA_signal_1511, \Midori/rounds/SelectedKey [5]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[3].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[67], key_s0[67]}), .I2 ({key_s1[3], key_s0[3]}), .O ({new_AGEMA_signal_1512, \Midori/rounds/SelectedKey [3]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[2].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[66], key_s0[66]}), .I2 ({key_s1[2], key_s0[2]}), .O ({new_AGEMA_signal_1513, \Midori/rounds/SelectedKey [2]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \Midori/rounds/MUXInst/gen_mux[1].mux_inst/Mmux_Q11 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[65], key_s0[65]}), .I2 ({key_s1[1], key_s0[1]}), .O ({new_AGEMA_signal_1514, \Midori/rounds/SelectedKey [1]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h9CC6 ) , .MASK ( 4'b1101 ), .INIT2 ( 16'hCCCC ) ) \Midori/rounds/Mxor_ProcessedKey<36>_xo<0>1 ( .I0 ({1'b0, enc_dec}), .I1 ({key_s1[100], key_s0[100]}), .I2 ({1'b0, \controller/roundCounter/count [2]}), .I3 ({1'b0, \controller/roundCounter/count [1]}), .O ({new_AGEMA_signal_1515, \Midori/rounds/Mxor_ProcessedKey<36>_xo<0> }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hDD7D7D7D88282828 ) , .MASK ( 6'b011101 ), .INIT2 ( 64'hDDDDDDDD88888888 ) ) \Midori/rounds/Mxor_ProcessedKey<36>_xo<0>2 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[36], key_s0[36]}), .I2 ({1'b0, \controller/roundCounter/count [1]}), .I3 ({1'b0, \controller/roundCounter/count [2]}), .I4 ({1'b0, \controller/roundCounter/count [3]}), .I5 ({new_AGEMA_signal_1515, \Midori/rounds/Mxor_ProcessedKey<36>_xo<0> }), .O ({new_AGEMA_signal_1609, \Midori/rounds/ProcessedKey [36]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC96C ) , .MASK ( 4'b1101 ), .INIT2 ( 16'hCCCC ) ) \Midori/rounds/Mxor_ProcessedKey<52>_xo<0>1 ( .I0 ({1'b0, enc_dec}), .I1 ({key_s1[116], key_s0[116]}), .I2 ({1'b0, \controller/roundCounter/count [2]}), .I3 ({1'b0, \controller/roundCounter/count [1]}), .O ({new_AGEMA_signal_1516, \Midori/rounds/Mxor_ProcessedKey<52>_xo<0> }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hD7D77DD782822882 ) , .MASK ( 6'b011101 ), .INIT2 ( 64'hDDDDDDDD88888888 ) ) \Midori/rounds/Mxor_ProcessedKey<52>_xo<0>2 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[52], key_s0[52]}), .I2 ({1'b0, \controller/roundCounter/count [2]}), .I3 ({1'b0, \controller/roundCounter/count [3]}), .I4 ({1'b0, \controller/roundCounter/count [1]}), .I5 ({new_AGEMA_signal_1516, \Midori/rounds/Mxor_ProcessedKey<52>_xo<0> }), .O ({new_AGEMA_signal_1610, \Midori/rounds/ProcessedKey [52]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hCCCC3963 ) , .MASK ( 5'b11101 ), .INIT2 ( 32'hCCCCCCCC ) ) \Midori/rounds/Mxor_ProcessedKey<48>_xo<0>1 ( .I0 ({1'b0, enc_dec}), .I1 ({key_s1[48], key_s0[48]}), .I2 ({1'b0, \controller/roundCounter/count [3]}), .I3 ({1'b0, \controller/roundCounter/count [2]}), .I4 ({1'b0, \controller/roundCounter/count [1]}), .O ({new_AGEMA_signal_1517, \Midori/rounds/Mxor_ProcessedKey<48>_xo<0> }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hBEBBBBEB14111141 ) , .MASK ( 6'b011101 ), .INIT2 ( 64'hEEEEEEEE44444444 ) ) \Midori/rounds/Mxor_ProcessedKey<48>_xo<0>2 ( .I0 ({1'b0, \controller/roundCounter/count [0]}), .I1 ({key_s1[112], key_s0[112]}), .I2 ({1'b0, \controller/roundCounter/count [1]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, \controller/roundCounter/count [3]}), .I5 ({new_AGEMA_signal_1517, \Midori/rounds/Mxor_ProcessedKey<48>_xo<0> }), .O ({new_AGEMA_signal_1611, \Midori/rounds/ProcessedKey [48]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h9 ) , .MASK ( 2'b10 ), .INIT2 ( 4'hA ) ) \Midori/rounds/Mxor_ProcessedKey<40>_xo<0>_SW0 ( .I0 ({key_s1[104], key_s0[104]}), .I1 ({1'b0, \controller/roundCounter/count [2]}), .O ({new_AGEMA_signal_1518, N9}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hAAAA033FAAAAFCC0 ) , .MASK ( 6'b011110 ), .INIT2 ( 64'hAAAAFFFFAAAA0000 ) ) \Midori/rounds/Mxor_ProcessedKey<40>_xo<0> ( .I0 ({key_s1[40], key_s0[40]}), .I1 ({1'b0, enc_dec}), .I2 ({1'b0, \controller/roundCounter/count [3]}), .I3 ({1'b0, \controller/roundCounter/count [1]}), .I4 ({1'b0, \controller/roundCounter/count [0]}), .I5 ({new_AGEMA_signal_1518, N9}), .O ({new_AGEMA_signal_1612, \Midori/rounds/ProcessedKey [40]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hA6 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \Midori/rounds/Mxor_ProcessedKey<48>_xo<0>2_SW0 ( .I0 ({key_s1[112], key_s0[112]}), .I1 ({1'b0, \controller/roundCounter/count [3]}), .I2 ({1'b0, \controller/roundCounter/count [1]}), .O ({new_AGEMA_signal_1519, N111}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA569 ) , .MASK ( 4'b1110 ), .INIT2 ( 16'hAAAA ) ) \Midori/rounds/Mxor_ProcessedKey<52>_xo<0>2_SW0 ( .I0 ({key_s1[52], key_s0[52]}), .I1 ({1'b0, \controller/roundCounter/count [3]}), .I2 ({1'b0, \controller/roundCounter/count [2]}), .I3 ({1'b0, \controller/roundCounter/count [1]}), .O ({new_AGEMA_signal_1520, N13}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \Midori/rounds/Mxor_ProcessedKey<44>_xo<0>1_SW0 ( .I0 ({key_s1[44], key_s0[44]}), .I1 ({key_s1[108], key_s0[108]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .O ({new_AGEMA_signal_1521, N15}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA666 ) , .MASK ( 4'b1110 ), .INIT2 ( 16'hAAAA ) ) \Midori/rounds/Mxor_ProcessedKey<36>_xo<0>2_SW0 ( .I0 ({key_s1[36], key_s0[36]}), .I1 ({1'b0, \controller/roundCounter/count_1_1_1069 }), .I2 ({1'b0, \controller/roundCounter/count [3]}), .I3 ({1'b0, \controller/roundCounter/count [2]}), .O ({new_AGEMA_signal_1522, N17}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \Midori/rounds/Mxor_ProcessedKey<32>_xo<0>1_SW0 ( .I0 ({key_s1[32], key_s0[32]}), .I1 ({key_s1[96], key_s0[96]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .O ({new_AGEMA_signal_1523, N19}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \Midori/rounds/Mxor_ProcessedKey<28>_xo<0>1_SW0 ( .I0 ({key_s1[28], key_s0[28]}), .I1 ({key_s1[92], key_s0[92]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .O ({new_AGEMA_signal_1524, N21}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \Midori/rounds/Mxor_ProcessedKey<24>_xo<0>1_SW0 ( .I0 ({key_s1[24], key_s0[24]}), .I1 ({key_s1[88], key_s0[88]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .O ({new_AGEMA_signal_1525, N23}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \Midori/rounds/Mxor_ProcessedKey<20>_xo<0>1_SW0 ( .I0 ({key_s1[20], key_s0[20]}), .I1 ({key_s1[84], key_s0[84]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .O ({new_AGEMA_signal_1526, N25}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \Midori/rounds/Mxor_ProcessedKey<12>_xo<0>1_SW0 ( .I0 ({key_s1[12], key_s0[12]}), .I1 ({key_s1[76], key_s0[76]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .O ({new_AGEMA_signal_1527, N27}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \Midori/rounds/Mxor_ProcessedKey<4>_xo<0>1_SW0 ( .I0 ({key_s1[4], key_s0[4]}), .I1 ({key_s1[68], key_s0[68]}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .O ({new_AGEMA_signal_1528, N29}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA596 ) , .MASK ( 4'b1110 ), .INIT2 ( 16'hAAAA ) ) \Midori/rounds/mul_input_Inst/gen_mux[40].mux_inst/Mmux_Q11_SW0 ( .I0 ({key_s1[104], key_s0[104]}), .I1 ({1'b0, \controller/roundCounter/count_3_2_1071 }), .I2 ({1'b0, \controller/roundCounter/count [2]}), .I3 ({1'b0, \controller/roundCounter/count [1]}), .O ({new_AGEMA_signal_1529, N34}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/Mxor_ProcessedKey<0>_xo<0> ( .s (\controller/roundCounter/count [2]), .b ({new_AGEMA_signal_1530, N36}), .a ({new_AGEMA_signal_1531, N37}), .c ({new_AGEMA_signal_1674, \Midori/rounds/ProcessedKey [0]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h2D88DD2878DD887D ) , .MASK ( 6'b011101 ), .INIT2 ( 64'hDDDDDDDD88888888 ) ) \Midori/rounds/Mxor_ProcessedKey<0>_xo<0>_F ( .I0 ({1'b0, \controller/roundCounter/count_0_1_1068 }), .I1 ({key_s1[0], key_s0[0]}), .I2 ({1'b0, \controller/roundCounter/count_1_1_1069 }), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, \controller/roundCounter/count [3]}), .I5 ({key_s1[64], key_s0[64]}), .O ({new_AGEMA_signal_1530, N36}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hBEBEBEAF14141405 ) , .MASK ( 6'b011011 ), .INIT2 ( 64'hFAFAFAFA50505050 ) ) \Midori/rounds/Mxor_ProcessedKey<0>_xo<0>_G ( .I0 ({1'b0, \controller/roundCounter/count_0_1_1068 }), .I1 ({1'b0, enc_dec}), .I2 ({key_s1[64], key_s0[64]}), .I3 ({1'b0, \controller/roundCounter/count_3_1_1066 }), .I4 ({1'b0, \controller/roundCounter/count_1_2_1072 }), .I5 ({key_s1[0], key_s0[0]}), .O ({new_AGEMA_signal_1531, N37}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/Mxor_ProcessedKey<16>_xo<0> ( .s (\controller/roundCounter/count [3]), .b ({new_AGEMA_signal_1532, N38}), .a ({new_AGEMA_signal_1533, N39}), .c ({new_AGEMA_signal_1675, \Midori/rounds/ProcessedKey [16]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE4C6286CB1937D39 ) , .MASK ( 6'b011011 ), .INIT2 ( 64'hF5F5F5F5A0A0A0A0 ) ) \Midori/rounds/Mxor_ProcessedKey<16>_xo<0>_F ( .I0 ({1'b0, \controller/roundCounter/count_0_1_1068 }), .I1 ({1'b0, \controller/roundCounter/count_2_1_1067 }), .I2 ({key_s1[16], key_s0[16]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, \controller/roundCounter/count_1_2_1072 }), .I5 ({key_s1[80], key_s0[80]}), .O ({new_AGEMA_signal_1532, N38}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9A569A56CF039A56 ) , .MASK ( 6'b110011 ), .INIT2 ( 64'hFC30FC30FC30FC30 ) ) \Midori/rounds/Mxor_ProcessedKey<16>_xo<0>_G ( .I0 ({1'b0, \controller/roundCounter/count_2_1_1067 }), .I1 ({1'b0, \controller/roundCounter/count_0_1_1068 }), .I2 ({key_s1[80], key_s0[80]}), .I3 ({key_s1[16], key_s0[16]}), .I4 ({1'b0, \controller/roundCounter/count_1_2_1072 }), .I5 ({1'b0, enc_dec}), .O ({new_AGEMA_signal_1533, N39}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/Mxor_ProcessedKey<56>_xo<0> ( .s (\controller/roundCounter/count [3]), .b ({new_AGEMA_signal_1534, N40}), .a ({new_AGEMA_signal_1535, N41}), .c ({new_AGEMA_signal_1676, \Midori/rounds/ProcessedKey [56]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hD282D77787D78222 ) , .MASK ( 6'b011101 ), .INIT2 ( 64'hDDDDDDDD88888888 ) ) \Midori/rounds/Mxor_ProcessedKey<56>_xo<0>_F ( .I0 ({1'b0, \controller/roundCounter/count_0_1_1068 }), .I1 ({key_s1[56], key_s0[56]}), .I2 ({1'b0, \controller/roundCounter/count_1_1_1069 }), .I3 ({1'b0, \controller/roundCounter/count_2_2_1070 }), .I4 ({1'b0, enc_dec}), .I5 ({key_s1[120], key_s0[120]}), .O ({new_AGEMA_signal_1534, N40}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hD7825F9382D70AC6 ) , .MASK ( 6'b011011 ), .INIT2 ( 64'hF5F5F5F5A0A0A0A0 ) ) \Midori/rounds/Mxor_ProcessedKey<56>_xo<0>_G ( .I0 ({1'b0, \controller/roundCounter/count_0_1_1068 }), .I1 ({1'b0, \controller/roundCounter/count_1_1_1069 }), .I2 ({key_s1[56], key_s0[56]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, \controller/roundCounter/count [2]}), .I5 ({key_s1[120], key_s0[120]}), .O ({new_AGEMA_signal_1535, N41}) ) ;
    INV \controller/roundCounter/Mcount_count_xor<0>11_INV_0 ( .I (\controller/roundCounter/count [0]), .O (Result[0]) ) ;
    ClockGatingController #(2) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[0].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1786, \Midori/rounds/mul_ResultXORkey [0]}), .I1 ({new_AGEMA_signal_1842, \Midori/rounds/mul_Result [48]}), .I2 ({new_AGEMA_signal_1466, \Midori/add_Result_Start [0]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1860, \Midori/rounds/roundResult_Reg/GEN[0].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[1].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1778, \Midori/rounds/mul_ResultXORkey [1]}), .I1 ({new_AGEMA_signal_1693, \Midori/rounds/mul_Result [49]}), .I2 ({new_AGEMA_signal_1462, \Midori/add_Result_Start [1]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1790, \Midori/rounds/roundResult_Reg/GEN[1].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[2].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1770, \Midori/rounds/mul_ResultXORkey [2]}), .I1 ({new_AGEMA_signal_1685, \Midori/rounds/mul_Result [50]}), .I2 ({new_AGEMA_signal_1418, \Midori/add_Result_Start [2]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1791, \Midori/rounds/roundResult_Reg/GEN[2].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[3].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1762, \Midori/rounds/mul_ResultXORkey [3]}), .I1 ({new_AGEMA_signal_1677, \Midori/rounds/mul_Result [51]}), .I2 ({new_AGEMA_signal_1374, \Midori/add_Result_Start [3]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1792, \Midori/rounds/roundResult_Reg/GEN[3].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[4].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1855, \Midori/rounds/mul_ResultXORkey [4]}), .I1 ({new_AGEMA_signal_1733, \Midori/rounds/mul_Result [44]}), .I2 ({new_AGEMA_signal_1330, \Midori/add_Result_Start [4]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1861, \Midori/rounds/roundResult_Reg/GEN[4].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[5].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1780, \Midori/rounds/mul_ResultXORkey [5]}), .I1 ({new_AGEMA_signal_1725, \Midori/rounds/mul_Result [45]}), .I2 ({new_AGEMA_signal_1286, \Midori/add_Result_Start [5]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1793, \Midori/rounds/roundResult_Reg/GEN[5].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[6].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1772, \Midori/rounds/mul_ResultXORkey [6]}), .I1 ({new_AGEMA_signal_1717, \Midori/rounds/mul_Result [46]}), .I2 ({new_AGEMA_signal_1242, \Midori/add_Result_Start [6]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1794, \Midori/rounds/roundResult_Reg/GEN[6].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[7].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1764, \Midori/rounds/mul_ResultXORkey [7]}), .I1 ({new_AGEMA_signal_1709, \Midori/rounds/mul_Result [47]}), .I2 ({new_AGEMA_signal_1222, \Midori/add_Result_Start [7]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1795, \Midori/rounds/roundResult_Reg/GEN[7].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[8].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1857, \Midori/rounds/mul_ResultXORkey [8]}), .I1 ({new_AGEMA_signal_1856, \Midori/rounds/mul_Result [8]}), .I2 ({new_AGEMA_signal_1218, \Midori/add_Result_Start [8]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1862, \Midori/rounds/roundResult_Reg/GEN[8].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[9].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1782, \Midori/rounds/mul_ResultXORkey [9]}), .I1 ({new_AGEMA_signal_1781, \Midori/rounds/mul_Result [9]}), .I2 ({new_AGEMA_signal_1214, \Midori/add_Result_Start [9]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1796, \Midori/rounds/roundResult_Reg/GEN[9].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[10].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1774, \Midori/rounds/mul_ResultXORkey [10]}), .I1 ({new_AGEMA_signal_1773, \Midori/rounds/mul_Result [10]}), .I2 ({new_AGEMA_signal_1458, \Midori/add_Result_Start [10]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1797, \Midori/rounds/roundResult_Reg/GEN[10].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[11].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1766, \Midori/rounds/mul_ResultXORkey [11]}), .I1 ({new_AGEMA_signal_1765, \Midori/rounds/mul_Result [11]}), .I2 ({new_AGEMA_signal_1454, \Midori/add_Result_Start [11]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1798, \Midori/rounds/roundResult_Reg/GEN[11].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[12].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1859, \Midori/rounds/mul_ResultXORkey [12]}), .I1 ({new_AGEMA_signal_1848, \Midori/rounds/mul_Result [20]}), .I2 ({new_AGEMA_signal_1450, \Midori/add_Result_Start [12]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1863, \Midori/rounds/roundResult_Reg/GEN[12].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[13].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1784, \Midori/rounds/mul_ResultXORkey [13]}), .I1 ({new_AGEMA_signal_1753, \Midori/rounds/mul_Result [21]}), .I2 ({new_AGEMA_signal_1446, \Midori/add_Result_Start [13]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1799, \Midori/rounds/roundResult_Reg/GEN[13].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[14].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1776, \Midori/rounds/mul_ResultXORkey [14]}), .I1 ({new_AGEMA_signal_1745, \Midori/rounds/mul_Result [22]}), .I2 ({new_AGEMA_signal_1442, \Midori/add_Result_Start [14]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1800, \Midori/rounds/roundResult_Reg/GEN[14].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[15].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1768, \Midori/rounds/mul_ResultXORkey [15]}), .I1 ({new_AGEMA_signal_1737, \Midori/rounds/mul_Result [23]}), .I2 ({new_AGEMA_signal_1438, \Midori/add_Result_Start [15]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1801, \Midori/rounds/roundResult_Reg/GEN[15].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[16].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1760, \Midori/rounds/mul_ResultXORkey [16]}), .I1 ({new_AGEMA_signal_1729, \Midori/rounds/mul_Result [36]}), .I2 ({new_AGEMA_signal_1434, \Midori/add_Result_Start [16]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1802, \Midori/rounds/roundResult_Reg/GEN[16].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[17].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1752, \Midori/rounds/mul_ResultXORkey [17]}), .I1 ({new_AGEMA_signal_1721, \Midori/rounds/mul_Result [37]}), .I2 ({new_AGEMA_signal_1430, \Midori/add_Result_Start [17]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1803, \Midori/rounds/roundResult_Reg/GEN[17].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[18].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1744, \Midori/rounds/mul_ResultXORkey [18]}), .I1 ({new_AGEMA_signal_1713, \Midori/rounds/mul_Result [38]}), .I2 ({new_AGEMA_signal_1426, \Midori/add_Result_Start [18]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1804, \Midori/rounds/roundResult_Reg/GEN[18].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[19].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1736, \Midori/rounds/mul_ResultXORkey [19]}), .I1 ({new_AGEMA_signal_1705, \Midori/rounds/mul_Result [39]}), .I2 ({new_AGEMA_signal_1422, \Midori/add_Result_Start [19]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1805, \Midori/rounds/roundResult_Reg/GEN[19].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[20].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1849, \Midori/rounds/mul_ResultXORkey [20]}), .I1 ({new_AGEMA_signal_1701, \Midori/rounds/mul_Result [56]}), .I2 ({new_AGEMA_signal_1414, \Midori/add_Result_Start [20]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1864, \Midori/rounds/roundResult_Reg/GEN[20].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[21].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1754, \Midori/rounds/mul_ResultXORkey [21]}), .I1 ({new_AGEMA_signal_1697, \Midori/rounds/mul_Result [57]}), .I2 ({new_AGEMA_signal_1410, \Midori/add_Result_Start [21]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1806, \Midori/rounds/roundResult_Reg/GEN[21].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[22].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1746, \Midori/rounds/mul_ResultXORkey [22]}), .I1 ({new_AGEMA_signal_1689, \Midori/rounds/mul_Result [58]}), .I2 ({new_AGEMA_signal_1406, \Midori/add_Result_Start [22]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1807, \Midori/rounds/roundResult_Reg/GEN[22].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[23].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1738, \Midori/rounds/mul_ResultXORkey [23]}), .I1 ({new_AGEMA_signal_1681, \Midori/rounds/mul_Result [59]}), .I2 ({new_AGEMA_signal_1402, \Midori/add_Result_Start [23]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1808, \Midori/rounds/roundResult_Reg/GEN[23].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[24].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1851, \Midori/rounds/mul_ResultXORkey [24]}), .I1 ({new_AGEMA_signal_1852, \Midori/rounds/mul_Result [28]}), .I2 ({new_AGEMA_signal_1398, \Midori/add_Result_Start [24]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1865, \Midori/rounds/roundResult_Reg/GEN[24].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[25].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1756, \Midori/rounds/mul_ResultXORkey [25]}), .I1 ({new_AGEMA_signal_1757, \Midori/rounds/mul_Result [29]}), .I2 ({new_AGEMA_signal_1394, \Midori/add_Result_Start [25]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1809, \Midori/rounds/roundResult_Reg/GEN[25].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[26].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1748, \Midori/rounds/mul_ResultXORkey [26]}), .I1 ({new_AGEMA_signal_1749, \Midori/rounds/mul_Result [30]}), .I2 ({new_AGEMA_signal_1390, \Midori/add_Result_Start [26]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1810, \Midori/rounds/roundResult_Reg/GEN[26].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[27].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1740, \Midori/rounds/mul_ResultXORkey [27]}), .I1 ({new_AGEMA_signal_1741, \Midori/rounds/mul_Result [31]}), .I2 ({new_AGEMA_signal_1386, \Midori/add_Result_Start [27]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1811, \Midori/rounds/roundResult_Reg/GEN[27].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[28].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1853, \Midori/rounds/mul_ResultXORkey [28]}), .I1 ({new_AGEMA_signal_1785, \Midori/rounds/mul_Result [0]}), .I2 ({new_AGEMA_signal_1382, \Midori/add_Result_Start [28]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1866, \Midori/rounds/roundResult_Reg/GEN[28].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[29].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1758, \Midori/rounds/mul_ResultXORkey [29]}), .I1 ({new_AGEMA_signal_1777, \Midori/rounds/mul_Result [1]}), .I2 ({new_AGEMA_signal_1378, \Midori/add_Result_Start [29]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1812, \Midori/rounds/roundResult_Reg/GEN[29].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[30].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1750, \Midori/rounds/mul_ResultXORkey [30]}), .I1 ({new_AGEMA_signal_1769, \Midori/rounds/mul_Result [2]}), .I2 ({new_AGEMA_signal_1370, \Midori/add_Result_Start [30]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1813, \Midori/rounds/roundResult_Reg/GEN[30].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[31].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1742, \Midori/rounds/mul_ResultXORkey [31]}), .I1 ({new_AGEMA_signal_1761, \Midori/rounds/mul_Result [3]}), .I2 ({new_AGEMA_signal_1366, \Midori/add_Result_Start [31]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1814, \Midori/rounds/roundResult_Reg/GEN[31].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[32].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1728, \Midori/rounds/mul_ResultXORkey [32]}), .I1 ({new_AGEMA_signal_1858, \Midori/rounds/mul_Result [12]}), .I2 ({new_AGEMA_signal_1362, \Midori/add_Result_Start [32]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1867, \Midori/rounds/roundResult_Reg/GEN[32].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[33].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1720, \Midori/rounds/mul_ResultXORkey [33]}), .I1 ({new_AGEMA_signal_1783, \Midori/rounds/mul_Result [13]}), .I2 ({new_AGEMA_signal_1358, \Midori/add_Result_Start [33]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1815, \Midori/rounds/roundResult_Reg/GEN[33].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[34].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1712, \Midori/rounds/mul_ResultXORkey [34]}), .I1 ({new_AGEMA_signal_1775, \Midori/rounds/mul_Result [14]}), .I2 ({new_AGEMA_signal_1354, \Midori/add_Result_Start [34]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1816, \Midori/rounds/roundResult_Reg/GEN[34].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[35].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1704, \Midori/rounds/mul_ResultXORkey [35]}), .I1 ({new_AGEMA_signal_1767, \Midori/rounds/mul_Result [15]}), .I2 ({new_AGEMA_signal_1350, \Midori/add_Result_Start [35]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1817, \Midori/rounds/roundResult_Reg/GEN[35].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[36].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1730, \Midori/rounds/mul_ResultXORkey [36]}), .I1 ({new_AGEMA_signal_1759, \Midori/rounds/mul_Result [16]}), .I2 ({new_AGEMA_signal_1346, \Midori/add_Result_Start [36]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1818, \Midori/rounds/roundResult_Reg/GEN[36].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[37].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1722, \Midori/rounds/mul_ResultXORkey [37]}), .I1 ({new_AGEMA_signal_1751, \Midori/rounds/mul_Result [17]}), .I2 ({new_AGEMA_signal_1342, \Midori/add_Result_Start [37]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1819, \Midori/rounds/roundResult_Reg/GEN[37].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[38].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1714, \Midori/rounds/mul_ResultXORkey [38]}), .I1 ({new_AGEMA_signal_1743, \Midori/rounds/mul_Result [18]}), .I2 ({new_AGEMA_signal_1338, \Midori/add_Result_Start [38]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1820, \Midori/rounds/roundResult_Reg/GEN[38].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[39].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1706, \Midori/rounds/mul_ResultXORkey [39]}), .I1 ({new_AGEMA_signal_1735, \Midori/rounds/mul_Result [19]}), .I2 ({new_AGEMA_signal_1334, \Midori/add_Result_Start [39]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1821, \Midori/rounds/roundResult_Reg/GEN[39].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[40].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1732, \Midori/rounds/mul_ResultXORkey [40]}), .I1 ({new_AGEMA_signal_1844, \Midori/rounds/mul_Result [52]}), .I2 ({new_AGEMA_signal_1326, \Midori/add_Result_Start [40]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1868, \Midori/rounds/roundResult_Reg/GEN[40].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[41].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1724, \Midori/rounds/mul_ResultXORkey [41]}), .I1 ({new_AGEMA_signal_1695, \Midori/rounds/mul_Result [53]}), .I2 ({new_AGEMA_signal_1322, \Midori/add_Result_Start [41]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1822, \Midori/rounds/roundResult_Reg/GEN[41].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[42].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1716, \Midori/rounds/mul_ResultXORkey [42]}), .I1 ({new_AGEMA_signal_1687, \Midori/rounds/mul_Result [54]}), .I2 ({new_AGEMA_signal_1318, \Midori/add_Result_Start [42]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1823, \Midori/rounds/roundResult_Reg/GEN[42].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[43].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1708, \Midori/rounds/mul_ResultXORkey [43]}), .I1 ({new_AGEMA_signal_1679, \Midori/rounds/mul_Result [55]}), .I2 ({new_AGEMA_signal_1314, \Midori/add_Result_Start [43]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1824, \Midori/rounds/roundResult_Reg/GEN[43].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[44].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1734, \Midori/rounds/mul_ResultXORkey [44]}), .I1 ({new_AGEMA_signal_1731, \Midori/rounds/mul_Result [40]}), .I2 ({new_AGEMA_signal_1310, \Midori/add_Result_Start [44]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1825, \Midori/rounds/roundResult_Reg/GEN[44].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[45].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1726, \Midori/rounds/mul_ResultXORkey [45]}), .I1 ({new_AGEMA_signal_1723, \Midori/rounds/mul_Result [41]}), .I2 ({new_AGEMA_signal_1306, \Midori/add_Result_Start [45]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1826, \Midori/rounds/roundResult_Reg/GEN[45].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[46].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1718, \Midori/rounds/mul_ResultXORkey [46]}), .I1 ({new_AGEMA_signal_1715, \Midori/rounds/mul_Result [42]}), .I2 ({new_AGEMA_signal_1302, \Midori/add_Result_Start [46]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1827, \Midori/rounds/roundResult_Reg/GEN[46].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[47].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1710, \Midori/rounds/mul_ResultXORkey [47]}), .I1 ({new_AGEMA_signal_1707, \Midori/rounds/mul_Result [43]}), .I2 ({new_AGEMA_signal_1298, \Midori/add_Result_Start [47]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1828, \Midori/rounds/roundResult_Reg/GEN[47].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[48].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1843, \Midori/rounds/mul_ResultXORkey [48]}), .I1 ({new_AGEMA_signal_1850, \Midori/rounds/mul_Result [24]}), .I2 ({new_AGEMA_signal_1294, \Midori/add_Result_Start [48]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1869, \Midori/rounds/roundResult_Reg/GEN[48].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[49].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1694, \Midori/rounds/mul_ResultXORkey [49]}), .I1 ({new_AGEMA_signal_1755, \Midori/rounds/mul_Result [25]}), .I2 ({new_AGEMA_signal_1290, \Midori/add_Result_Start [49]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1829, \Midori/rounds/roundResult_Reg/GEN[49].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[50].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1686, \Midori/rounds/mul_ResultXORkey [50]}), .I1 ({new_AGEMA_signal_1747, \Midori/rounds/mul_Result [26]}), .I2 ({new_AGEMA_signal_1282, \Midori/add_Result_Start [50]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1830, \Midori/rounds/roundResult_Reg/GEN[50].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[51].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1678, \Midori/rounds/mul_ResultXORkey [51]}), .I1 ({new_AGEMA_signal_1739, \Midori/rounds/mul_Result [27]}), .I2 ({new_AGEMA_signal_1278, \Midori/add_Result_Start [51]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1831, \Midori/rounds/roundResult_Reg/GEN[51].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[52].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1845, \Midori/rounds/mul_ResultXORkey [52]}), .I1 ({new_AGEMA_signal_1854, \Midori/rounds/mul_Result [4]}), .I2 ({new_AGEMA_signal_1274, \Midori/add_Result_Start [52]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1870, \Midori/rounds/roundResult_Reg/GEN[52].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[53].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1696, \Midori/rounds/mul_ResultXORkey [53]}), .I1 ({new_AGEMA_signal_1779, \Midori/rounds/mul_Result [5]}), .I2 ({new_AGEMA_signal_1270, \Midori/add_Result_Start [53]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1832, \Midori/rounds/roundResult_Reg/GEN[53].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[54].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1688, \Midori/rounds/mul_ResultXORkey [54]}), .I1 ({new_AGEMA_signal_1771, \Midori/rounds/mul_Result [6]}), .I2 ({new_AGEMA_signal_1266, \Midori/add_Result_Start [54]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1833, \Midori/rounds/roundResult_Reg/GEN[54].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[55].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1680, \Midori/rounds/mul_ResultXORkey [55]}), .I1 ({new_AGEMA_signal_1763, \Midori/rounds/mul_Result [7]}), .I2 ({new_AGEMA_signal_1262, \Midori/add_Result_Start [55]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1834, \Midori/rounds/roundResult_Reg/GEN[55].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[56].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1702, \Midori/rounds/mul_ResultXORkey [56]}), .I1 ({new_AGEMA_signal_1727, \Midori/rounds/mul_Result [32]}), .I2 ({new_AGEMA_signal_1258, \Midori/add_Result_Start [56]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1835, \Midori/rounds/roundResult_Reg/GEN[56].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[57].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1698, \Midori/rounds/mul_ResultXORkey [57]}), .I1 ({new_AGEMA_signal_1719, \Midori/rounds/mul_Result [33]}), .I2 ({new_AGEMA_signal_1254, \Midori/add_Result_Start [57]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1836, \Midori/rounds/roundResult_Reg/GEN[57].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[58].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1690, \Midori/rounds/mul_ResultXORkey [58]}), .I1 ({new_AGEMA_signal_1711, \Midori/rounds/mul_Result [34]}), .I2 ({new_AGEMA_signal_1250, \Midori/add_Result_Start [58]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1837, \Midori/rounds/roundResult_Reg/GEN[58].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[59].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1682, \Midori/rounds/mul_ResultXORkey [59]}), .I1 ({new_AGEMA_signal_1703, \Midori/rounds/mul_Result [35]}), .I2 ({new_AGEMA_signal_1246, \Midori/add_Result_Start [59]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1838, \Midori/rounds/roundResult_Reg/GEN[59].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[60].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1847, \Midori/rounds/mul_ResultXORkey [60]}), .I1 ({new_AGEMA_signal_1846, \Midori/rounds/mul_Result [60]}), .I2 ({new_AGEMA_signal_1238, \Midori/add_Result_Start [60]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1871, \Midori/rounds/roundResult_Reg/GEN[60].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[61].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1700, \Midori/rounds/mul_ResultXORkey [61]}), .I1 ({new_AGEMA_signal_1699, \Midori/rounds/mul_Result [61]}), .I2 ({new_AGEMA_signal_1234, \Midori/add_Result_Start [61]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1839, \Midori/rounds/roundResult_Reg/GEN[61].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[62].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1692, \Midori/rounds/mul_ResultXORkey [62]}), .I1 ({new_AGEMA_signal_1691, \Midori/rounds/mul_Result [62]}), .I2 ({new_AGEMA_signal_1230, \Midori/add_Result_Start [62]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1840, \Midori/rounds/roundResult_Reg/GEN[62].SFF/DQ }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \Midori/rounds/roundResult_Reg/GEN[63].SFF/LUTINST ( .I0 ({new_AGEMA_signal_1684, \Midori/rounds/mul_ResultXORkey [63]}), .I1 ({new_AGEMA_signal_1683, \Midori/rounds/mul_Result [63]}), .I2 ({new_AGEMA_signal_1226, \Midori/add_Result_Start [63]}), .I3 ({1'b0, enc_dec}), .I4 ({1'b0, reset}), .O ({new_AGEMA_signal_1841, \Midori/rounds/roundResult_Reg/GEN[63].SFF/DQ }) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[0].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1083, \Midori/rounds/roundResult_Reg/GEN[0].SFF/Q_663 }), .I1 ({new_AGEMA_signal_1084, \Midori/rounds/roundResult_Reg/GEN[1].SFF/Q_664 }), .I2 ({new_AGEMA_signal_1085, \Midori/rounds/roundResult_Reg/GEN[2].SFF/Q_665 }), .I3 ({new_AGEMA_signal_1086, \Midori/rounds/roundResult_Reg/GEN[3].SFF/Q_666 }), .clk (clk), .r ({Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .O ({new_AGEMA_signal_1087, \Midori/rounds_Output [0]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[0].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1083, \Midori/rounds/roundResult_Reg/GEN[0].SFF/Q_663 }), .I1 ({new_AGEMA_signal_1084, \Midori/rounds/roundResult_Reg/GEN[1].SFF/Q_664 }), .I2 ({new_AGEMA_signal_1085, \Midori/rounds/roundResult_Reg/GEN[2].SFF/Q_665 }), .I3 ({new_AGEMA_signal_1086, \Midori/rounds/roundResult_Reg/GEN[3].SFF/Q_666 }), .clk (clk), .r ({Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16]}), .O ({new_AGEMA_signal_1088, \Midori/rounds_Output [1]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[0].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1083, \Midori/rounds/roundResult_Reg/GEN[0].SFF/Q_663 }), .I1 ({new_AGEMA_signal_1084, \Midori/rounds/roundResult_Reg/GEN[1].SFF/Q_664 }), .I2 ({new_AGEMA_signal_1085, \Midori/rounds/roundResult_Reg/GEN[2].SFF/Q_665 }), .I3 ({new_AGEMA_signal_1086, \Midori/rounds/roundResult_Reg/GEN[3].SFF/Q_666 }), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32]}), .O ({new_AGEMA_signal_1089, \Midori/rounds_Output [2]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[0].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1083, \Midori/rounds/roundResult_Reg/GEN[0].SFF/Q_663 }), .I1 ({new_AGEMA_signal_1084, \Midori/rounds/roundResult_Reg/GEN[1].SFF/Q_664 }), .I2 ({new_AGEMA_signal_1085, \Midori/rounds/roundResult_Reg/GEN[2].SFF/Q_665 }), .I3 ({new_AGEMA_signal_1086, \Midori/rounds/roundResult_Reg/GEN[3].SFF/Q_666 }), .clk (clk), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .O ({new_AGEMA_signal_1090, \Midori/rounds_Output [3]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[1].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1091, \Midori/rounds/roundResult_Reg/GEN[4].SFF/Q_667 }), .I1 ({new_AGEMA_signal_1092, \Midori/rounds/roundResult_Reg/GEN[5].SFF/Q_668 }), .I2 ({new_AGEMA_signal_1093, \Midori/rounds/roundResult_Reg/GEN[6].SFF/Q_669 }), .I3 ({new_AGEMA_signal_1094, \Midori/rounds/roundResult_Reg/GEN[7].SFF/Q_670 }), .clk (clk), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64]}), .O ({new_AGEMA_signal_1095, \Midori/rounds_Output [4]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[1].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1091, \Midori/rounds/roundResult_Reg/GEN[4].SFF/Q_667 }), .I1 ({new_AGEMA_signal_1092, \Midori/rounds/roundResult_Reg/GEN[5].SFF/Q_668 }), .I2 ({new_AGEMA_signal_1093, \Midori/rounds/roundResult_Reg/GEN[6].SFF/Q_669 }), .I3 ({new_AGEMA_signal_1094, \Midori/rounds/roundResult_Reg/GEN[7].SFF/Q_670 }), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .O ({new_AGEMA_signal_1096, \Midori/rounds_Output [5]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[1].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1091, \Midori/rounds/roundResult_Reg/GEN[4].SFF/Q_667 }), .I1 ({new_AGEMA_signal_1092, \Midori/rounds/roundResult_Reg/GEN[5].SFF/Q_668 }), .I2 ({new_AGEMA_signal_1093, \Midori/rounds/roundResult_Reg/GEN[6].SFF/Q_669 }), .I3 ({new_AGEMA_signal_1094, \Midori/rounds/roundResult_Reg/GEN[7].SFF/Q_670 }), .clk (clk), .r ({Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .O ({new_AGEMA_signal_1097, \Midori/rounds_Output [6]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[1].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1091, \Midori/rounds/roundResult_Reg/GEN[4].SFF/Q_667 }), .I1 ({new_AGEMA_signal_1092, \Midori/rounds/roundResult_Reg/GEN[5].SFF/Q_668 }), .I2 ({new_AGEMA_signal_1093, \Midori/rounds/roundResult_Reg/GEN[6].SFF/Q_669 }), .I3 ({new_AGEMA_signal_1094, \Midori/rounds/roundResult_Reg/GEN[7].SFF/Q_670 }), .clk (clk), .r ({Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112]}), .O ({new_AGEMA_signal_1098, \Midori/rounds_Output [7]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[2].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1099, \Midori/rounds/roundResult_Reg/GEN[8].SFF/Q_671 }), .I1 ({new_AGEMA_signal_1100, \Midori/rounds/roundResult_Reg/GEN[9].SFF/Q_672 }), .I2 ({new_AGEMA_signal_1101, \Midori/rounds/roundResult_Reg/GEN[10].SFF/Q_673 }), .I3 ({new_AGEMA_signal_1102, \Midori/rounds/roundResult_Reg/GEN[11].SFF/Q_674 }), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128]}), .O ({new_AGEMA_signal_1103, \Midori/rounds_Output [8]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[2].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1099, \Midori/rounds/roundResult_Reg/GEN[8].SFF/Q_671 }), .I1 ({new_AGEMA_signal_1100, \Midori/rounds/roundResult_Reg/GEN[9].SFF/Q_672 }), .I2 ({new_AGEMA_signal_1101, \Midori/rounds/roundResult_Reg/GEN[10].SFF/Q_673 }), .I3 ({new_AGEMA_signal_1102, \Midori/rounds/roundResult_Reg/GEN[11].SFF/Q_674 }), .clk (clk), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .O ({new_AGEMA_signal_1104, \Midori/rounds_Output [9]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[2].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1099, \Midori/rounds/roundResult_Reg/GEN[8].SFF/Q_671 }), .I1 ({new_AGEMA_signal_1100, \Midori/rounds/roundResult_Reg/GEN[9].SFF/Q_672 }), .I2 ({new_AGEMA_signal_1101, \Midori/rounds/roundResult_Reg/GEN[10].SFF/Q_673 }), .I3 ({new_AGEMA_signal_1102, \Midori/rounds/roundResult_Reg/GEN[11].SFF/Q_674 }), .clk (clk), .r ({Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .O ({new_AGEMA_signal_1105, \Midori/rounds_Output [10]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[2].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1099, \Midori/rounds/roundResult_Reg/GEN[8].SFF/Q_671 }), .I1 ({new_AGEMA_signal_1100, \Midori/rounds/roundResult_Reg/GEN[9].SFF/Q_672 }), .I2 ({new_AGEMA_signal_1101, \Midori/rounds/roundResult_Reg/GEN[10].SFF/Q_673 }), .I3 ({new_AGEMA_signal_1102, \Midori/rounds/roundResult_Reg/GEN[11].SFF/Q_674 }), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180], Fresh[179], Fresh[178], Fresh[177], Fresh[176]}), .O ({new_AGEMA_signal_1106, \Midori/rounds_Output [11]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[3].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1107, \Midori/rounds/roundResult_Reg/GEN[12].SFF/Q_675 }), .I1 ({new_AGEMA_signal_1108, \Midori/rounds/roundResult_Reg/GEN[13].SFF/Q_676 }), .I2 ({new_AGEMA_signal_1109, \Midori/rounds/roundResult_Reg/GEN[14].SFF/Q_677 }), .I3 ({new_AGEMA_signal_1110, \Midori/rounds/roundResult_Reg/GEN[15].SFF/Q_678 }), .clk (clk), .r ({Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .O ({new_AGEMA_signal_1111, \Midori/rounds_Output [12]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[3].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1107, \Midori/rounds/roundResult_Reg/GEN[12].SFF/Q_675 }), .I1 ({new_AGEMA_signal_1108, \Midori/rounds/roundResult_Reg/GEN[13].SFF/Q_676 }), .I2 ({new_AGEMA_signal_1109, \Midori/rounds/roundResult_Reg/GEN[14].SFF/Q_677 }), .I3 ({new_AGEMA_signal_1110, \Midori/rounds/roundResult_Reg/GEN[15].SFF/Q_678 }), .clk (clk), .r ({Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208]}), .O ({new_AGEMA_signal_1112, \Midori/rounds_Output [13]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[3].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1107, \Midori/rounds/roundResult_Reg/GEN[12].SFF/Q_675 }), .I1 ({new_AGEMA_signal_1108, \Midori/rounds/roundResult_Reg/GEN[13].SFF/Q_676 }), .I2 ({new_AGEMA_signal_1109, \Midori/rounds/roundResult_Reg/GEN[14].SFF/Q_677 }), .I3 ({new_AGEMA_signal_1110, \Midori/rounds/roundResult_Reg/GEN[15].SFF/Q_678 }), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224]}), .O ({new_AGEMA_signal_1113, \Midori/rounds_Output [14]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[3].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1107, \Midori/rounds/roundResult_Reg/GEN[12].SFF/Q_675 }), .I1 ({new_AGEMA_signal_1108, \Midori/rounds/roundResult_Reg/GEN[13].SFF/Q_676 }), .I2 ({new_AGEMA_signal_1109, \Midori/rounds/roundResult_Reg/GEN[14].SFF/Q_677 }), .I3 ({new_AGEMA_signal_1110, \Midori/rounds/roundResult_Reg/GEN[15].SFF/Q_678 }), .clk (clk), .r ({Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .O ({new_AGEMA_signal_1114, \Midori/rounds_Output [15]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[4].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1115, \Midori/rounds/roundResult_Reg/GEN[16].SFF/Q_679 }), .I1 ({new_AGEMA_signal_1116, \Midori/rounds/roundResult_Reg/GEN[17].SFF/Q_680 }), .I2 ({new_AGEMA_signal_1117, \Midori/rounds/roundResult_Reg/GEN[18].SFF/Q_681 }), .I3 ({new_AGEMA_signal_1118, \Midori/rounds/roundResult_Reg/GEN[19].SFF/Q_682 }), .clk (clk), .r ({Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256]}), .O ({new_AGEMA_signal_1119, \Midori/rounds_Output [16]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[4].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1115, \Midori/rounds/roundResult_Reg/GEN[16].SFF/Q_679 }), .I1 ({new_AGEMA_signal_1116, \Midori/rounds/roundResult_Reg/GEN[17].SFF/Q_680 }), .I2 ({new_AGEMA_signal_1117, \Midori/rounds/roundResult_Reg/GEN[18].SFF/Q_681 }), .I3 ({new_AGEMA_signal_1118, \Midori/rounds/roundResult_Reg/GEN[19].SFF/Q_682 }), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272]}), .O ({new_AGEMA_signal_1120, \Midori/rounds_Output [17]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[4].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1115, \Midori/rounds/roundResult_Reg/GEN[16].SFF/Q_679 }), .I1 ({new_AGEMA_signal_1116, \Midori/rounds/roundResult_Reg/GEN[17].SFF/Q_680 }), .I2 ({new_AGEMA_signal_1117, \Midori/rounds/roundResult_Reg/GEN[18].SFF/Q_681 }), .I3 ({new_AGEMA_signal_1118, \Midori/rounds/roundResult_Reg/GEN[19].SFF/Q_682 }), .clk (clk), .r ({Fresh[303], Fresh[302], Fresh[301], Fresh[300], Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .O ({new_AGEMA_signal_1121, \Midori/rounds_Output [18]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[4].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1115, \Midori/rounds/roundResult_Reg/GEN[16].SFF/Q_679 }), .I1 ({new_AGEMA_signal_1116, \Midori/rounds/roundResult_Reg/GEN[17].SFF/Q_680 }), .I2 ({new_AGEMA_signal_1117, \Midori/rounds/roundResult_Reg/GEN[18].SFF/Q_681 }), .I3 ({new_AGEMA_signal_1118, \Midori/rounds/roundResult_Reg/GEN[19].SFF/Q_682 }), .clk (clk), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304]}), .O ({new_AGEMA_signal_1122, \Midori/rounds_Output [19]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[5].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1123, \Midori/rounds/roundResult_Reg/GEN[20].SFF/Q_683 }), .I1 ({new_AGEMA_signal_1124, \Midori/rounds/roundResult_Reg/GEN[21].SFF/Q_684 }), .I2 ({new_AGEMA_signal_1125, \Midori/rounds/roundResult_Reg/GEN[22].SFF/Q_685 }), .I3 ({new_AGEMA_signal_1126, \Midori/rounds/roundResult_Reg/GEN[23].SFF/Q_686 }), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .O ({new_AGEMA_signal_1127, \Midori/rounds_Output [20]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[5].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1123, \Midori/rounds/roundResult_Reg/GEN[20].SFF/Q_683 }), .I1 ({new_AGEMA_signal_1124, \Midori/rounds/roundResult_Reg/GEN[21].SFF/Q_684 }), .I2 ({new_AGEMA_signal_1125, \Midori/rounds/roundResult_Reg/GEN[22].SFF/Q_685 }), .I3 ({new_AGEMA_signal_1126, \Midori/rounds/roundResult_Reg/GEN[23].SFF/Q_686 }), .clk (clk), .r ({Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .O ({new_AGEMA_signal_1128, \Midori/rounds_Output [21]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[5].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1123, \Midori/rounds/roundResult_Reg/GEN[20].SFF/Q_683 }), .I1 ({new_AGEMA_signal_1124, \Midori/rounds/roundResult_Reg/GEN[21].SFF/Q_684 }), .I2 ({new_AGEMA_signal_1125, \Midori/rounds/roundResult_Reg/GEN[22].SFF/Q_685 }), .I3 ({new_AGEMA_signal_1126, \Midori/rounds/roundResult_Reg/GEN[23].SFF/Q_686 }), .clk (clk), .r ({Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360], Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352]}), .O ({new_AGEMA_signal_1129, \Midori/rounds_Output [22]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[5].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1123, \Midori/rounds/roundResult_Reg/GEN[20].SFF/Q_683 }), .I1 ({new_AGEMA_signal_1124, \Midori/rounds/roundResult_Reg/GEN[21].SFF/Q_684 }), .I2 ({new_AGEMA_signal_1125, \Midori/rounds/roundResult_Reg/GEN[22].SFF/Q_685 }), .I3 ({new_AGEMA_signal_1126, \Midori/rounds/roundResult_Reg/GEN[23].SFF/Q_686 }), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368]}), .O ({new_AGEMA_signal_1130, \Midori/rounds_Output [23]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[6].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1131, \Midori/rounds/roundResult_Reg/GEN[24].SFF/Q_687 }), .I1 ({new_AGEMA_signal_1132, \Midori/rounds/roundResult_Reg/GEN[25].SFF/Q_688 }), .I2 ({new_AGEMA_signal_1133, \Midori/rounds/roundResult_Reg/GEN[26].SFF/Q_689 }), .I3 ({new_AGEMA_signal_1134, \Midori/rounds/roundResult_Reg/GEN[27].SFF/Q_690 }), .clk (clk), .r ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .O ({new_AGEMA_signal_1135, \Midori/rounds_Output [24]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[6].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1131, \Midori/rounds/roundResult_Reg/GEN[24].SFF/Q_687 }), .I1 ({new_AGEMA_signal_1132, \Midori/rounds/roundResult_Reg/GEN[25].SFF/Q_688 }), .I2 ({new_AGEMA_signal_1133, \Midori/rounds/roundResult_Reg/GEN[26].SFF/Q_689 }), .I3 ({new_AGEMA_signal_1134, \Midori/rounds/roundResult_Reg/GEN[27].SFF/Q_690 }), .clk (clk), .r ({Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .O ({new_AGEMA_signal_1136, \Midori/rounds_Output [25]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[6].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1131, \Midori/rounds/roundResult_Reg/GEN[24].SFF/Q_687 }), .I1 ({new_AGEMA_signal_1132, \Midori/rounds/roundResult_Reg/GEN[25].SFF/Q_688 }), .I2 ({new_AGEMA_signal_1133, \Midori/rounds/roundResult_Reg/GEN[26].SFF/Q_689 }), .I3 ({new_AGEMA_signal_1134, \Midori/rounds/roundResult_Reg/GEN[27].SFF/Q_690 }), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420], Fresh[419], Fresh[418], Fresh[417], Fresh[416]}), .O ({new_AGEMA_signal_1137, \Midori/rounds_Output [26]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[6].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1131, \Midori/rounds/roundResult_Reg/GEN[24].SFF/Q_687 }), .I1 ({new_AGEMA_signal_1132, \Midori/rounds/roundResult_Reg/GEN[25].SFF/Q_688 }), .I2 ({new_AGEMA_signal_1133, \Midori/rounds/roundResult_Reg/GEN[26].SFF/Q_689 }), .I3 ({new_AGEMA_signal_1134, \Midori/rounds/roundResult_Reg/GEN[27].SFF/Q_690 }), .clk (clk), .r ({Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .O ({new_AGEMA_signal_1138, \Midori/rounds_Output [27]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[7].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1139, \Midori/rounds/roundResult_Reg/GEN[28].SFF/Q_691 }), .I1 ({new_AGEMA_signal_1140, \Midori/rounds/roundResult_Reg/GEN[29].SFF/Q_692 }), .I2 ({new_AGEMA_signal_1141, \Midori/rounds/roundResult_Reg/GEN[30].SFF/Q_693 }), .I3 ({new_AGEMA_signal_1142, \Midori/rounds/roundResult_Reg/GEN[31].SFF/Q_694 }), .clk (clk), .r ({Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448]}), .O ({new_AGEMA_signal_1143, \Midori/rounds_Output [28]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[7].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1139, \Midori/rounds/roundResult_Reg/GEN[28].SFF/Q_691 }), .I1 ({new_AGEMA_signal_1140, \Midori/rounds/roundResult_Reg/GEN[29].SFF/Q_692 }), .I2 ({new_AGEMA_signal_1141, \Midori/rounds/roundResult_Reg/GEN[30].SFF/Q_693 }), .I3 ({new_AGEMA_signal_1142, \Midori/rounds/roundResult_Reg/GEN[31].SFF/Q_694 }), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464]}), .O ({new_AGEMA_signal_1144, \Midori/rounds_Output [29]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[7].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1139, \Midori/rounds/roundResult_Reg/GEN[28].SFF/Q_691 }), .I1 ({new_AGEMA_signal_1140, \Midori/rounds/roundResult_Reg/GEN[29].SFF/Q_692 }), .I2 ({new_AGEMA_signal_1141, \Midori/rounds/roundResult_Reg/GEN[30].SFF/Q_693 }), .I3 ({new_AGEMA_signal_1142, \Midori/rounds/roundResult_Reg/GEN[31].SFF/Q_694 }), .clk (clk), .r ({Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .O ({new_AGEMA_signal_1145, \Midori/rounds_Output [30]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[7].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1139, \Midori/rounds/roundResult_Reg/GEN[28].SFF/Q_691 }), .I1 ({new_AGEMA_signal_1140, \Midori/rounds/roundResult_Reg/GEN[29].SFF/Q_692 }), .I2 ({new_AGEMA_signal_1141, \Midori/rounds/roundResult_Reg/GEN[30].SFF/Q_693 }), .I3 ({new_AGEMA_signal_1142, \Midori/rounds/roundResult_Reg/GEN[31].SFF/Q_694 }), .clk (clk), .r ({Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496]}), .O ({new_AGEMA_signal_1146, \Midori/rounds_Output [31]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[8].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1147, \Midori/rounds/roundResult_Reg/GEN[32].SFF/Q_695 }), .I1 ({new_AGEMA_signal_1148, \Midori/rounds/roundResult_Reg/GEN[33].SFF/Q_696 }), .I2 ({new_AGEMA_signal_1149, \Midori/rounds/roundResult_Reg/GEN[34].SFF/Q_697 }), .I3 ({new_AGEMA_signal_1150, \Midori/rounds/roundResult_Reg/GEN[35].SFF/Q_698 }), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512]}), .O ({new_AGEMA_signal_1151, \Midori/rounds_Output [32]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[8].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1147, \Midori/rounds/roundResult_Reg/GEN[32].SFF/Q_695 }), .I1 ({new_AGEMA_signal_1148, \Midori/rounds/roundResult_Reg/GEN[33].SFF/Q_696 }), .I2 ({new_AGEMA_signal_1149, \Midori/rounds/roundResult_Reg/GEN[34].SFF/Q_697 }), .I3 ({new_AGEMA_signal_1150, \Midori/rounds/roundResult_Reg/GEN[35].SFF/Q_698 }), .clk (clk), .r ({Fresh[543], Fresh[542], Fresh[541], Fresh[540], Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .O ({new_AGEMA_signal_1152, \Midori/rounds_Output [33]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[8].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1147, \Midori/rounds/roundResult_Reg/GEN[32].SFF/Q_695 }), .I1 ({new_AGEMA_signal_1148, \Midori/rounds/roundResult_Reg/GEN[33].SFF/Q_696 }), .I2 ({new_AGEMA_signal_1149, \Midori/rounds/roundResult_Reg/GEN[34].SFF/Q_697 }), .I3 ({new_AGEMA_signal_1150, \Midori/rounds/roundResult_Reg/GEN[35].SFF/Q_698 }), .clk (clk), .r ({Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544]}), .O ({new_AGEMA_signal_1153, \Midori/rounds_Output [34]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[8].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1147, \Midori/rounds/roundResult_Reg/GEN[32].SFF/Q_695 }), .I1 ({new_AGEMA_signal_1148, \Midori/rounds/roundResult_Reg/GEN[33].SFF/Q_696 }), .I2 ({new_AGEMA_signal_1149, \Midori/rounds/roundResult_Reg/GEN[34].SFF/Q_697 }), .I3 ({new_AGEMA_signal_1150, \Midori/rounds/roundResult_Reg/GEN[35].SFF/Q_698 }), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .O ({new_AGEMA_signal_1154, \Midori/rounds_Output [35]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[9].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1155, \Midori/rounds/roundResult_Reg/GEN[36].SFF/Q_699 }), .I1 ({new_AGEMA_signal_1156, \Midori/rounds/roundResult_Reg/GEN[37].SFF/Q_700 }), .I2 ({new_AGEMA_signal_1157, \Midori/rounds/roundResult_Reg/GEN[38].SFF/Q_701 }), .I3 ({new_AGEMA_signal_1158, \Midori/rounds/roundResult_Reg/GEN[39].SFF/Q_702 }), .clk (clk), .r ({Fresh[591], Fresh[590], Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .O ({new_AGEMA_signal_1159, \Midori/rounds_Output [36]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[9].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1155, \Midori/rounds/roundResult_Reg/GEN[36].SFF/Q_699 }), .I1 ({new_AGEMA_signal_1156, \Midori/rounds/roundResult_Reg/GEN[37].SFF/Q_700 }), .I2 ({new_AGEMA_signal_1157, \Midori/rounds/roundResult_Reg/GEN[38].SFF/Q_701 }), .I3 ({new_AGEMA_signal_1158, \Midori/rounds/roundResult_Reg/GEN[39].SFF/Q_702 }), .clk (clk), .r ({Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600], Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592]}), .O ({new_AGEMA_signal_1160, \Midori/rounds_Output [37]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[9].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1155, \Midori/rounds/roundResult_Reg/GEN[36].SFF/Q_699 }), .I1 ({new_AGEMA_signal_1156, \Midori/rounds/roundResult_Reg/GEN[37].SFF/Q_700 }), .I2 ({new_AGEMA_signal_1157, \Midori/rounds/roundResult_Reg/GEN[38].SFF/Q_701 }), .I3 ({new_AGEMA_signal_1158, \Midori/rounds/roundResult_Reg/GEN[39].SFF/Q_702 }), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610], Fresh[609], Fresh[608]}), .O ({new_AGEMA_signal_1161, \Midori/rounds_Output [38]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[9].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1155, \Midori/rounds/roundResult_Reg/GEN[36].SFF/Q_699 }), .I1 ({new_AGEMA_signal_1156, \Midori/rounds/roundResult_Reg/GEN[37].SFF/Q_700 }), .I2 ({new_AGEMA_signal_1157, \Midori/rounds/roundResult_Reg/GEN[38].SFF/Q_701 }), .I3 ({new_AGEMA_signal_1158, \Midori/rounds/roundResult_Reg/GEN[39].SFF/Q_702 }), .clk (clk), .r ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .O ({new_AGEMA_signal_1162, \Midori/rounds_Output [39]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[10].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1163, \Midori/rounds/roundResult_Reg/GEN[40].SFF/Q_703 }), .I1 ({new_AGEMA_signal_1164, \Midori/rounds/roundResult_Reg/GEN[41].SFF/Q_704 }), .I2 ({new_AGEMA_signal_1165, \Midori/rounds/roundResult_Reg/GEN[42].SFF/Q_705 }), .I3 ({new_AGEMA_signal_1166, \Midori/rounds/roundResult_Reg/GEN[43].SFF/Q_706 }), .clk (clk), .r ({Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .O ({new_AGEMA_signal_1167, \Midori/rounds_Output [40]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[10].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1163, \Midori/rounds/roundResult_Reg/GEN[40].SFF/Q_703 }), .I1 ({new_AGEMA_signal_1164, \Midori/rounds/roundResult_Reg/GEN[41].SFF/Q_704 }), .I2 ({new_AGEMA_signal_1165, \Midori/rounds/roundResult_Reg/GEN[42].SFF/Q_705 }), .I3 ({new_AGEMA_signal_1166, \Midori/rounds/roundResult_Reg/GEN[43].SFF/Q_706 }), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660], Fresh[659], Fresh[658], Fresh[657], Fresh[656]}), .O ({new_AGEMA_signal_1168, \Midori/rounds_Output [41]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[10].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1163, \Midori/rounds/roundResult_Reg/GEN[40].SFF/Q_703 }), .I1 ({new_AGEMA_signal_1164, \Midori/rounds/roundResult_Reg/GEN[41].SFF/Q_704 }), .I2 ({new_AGEMA_signal_1165, \Midori/rounds/roundResult_Reg/GEN[42].SFF/Q_705 }), .I3 ({new_AGEMA_signal_1166, \Midori/rounds/roundResult_Reg/GEN[43].SFF/Q_706 }), .clk (clk), .r ({Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .O ({new_AGEMA_signal_1169, \Midori/rounds_Output [42]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[10].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1163, \Midori/rounds/roundResult_Reg/GEN[40].SFF/Q_703 }), .I1 ({new_AGEMA_signal_1164, \Midori/rounds/roundResult_Reg/GEN[41].SFF/Q_704 }), .I2 ({new_AGEMA_signal_1165, \Midori/rounds/roundResult_Reg/GEN[42].SFF/Q_705 }), .I3 ({new_AGEMA_signal_1166, \Midori/rounds/roundResult_Reg/GEN[43].SFF/Q_706 }), .clk (clk), .r ({Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688]}), .O ({new_AGEMA_signal_1170, \Midori/rounds_Output [43]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[11].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1171, \Midori/rounds/roundResult_Reg/GEN[44].SFF/Q_707 }), .I1 ({new_AGEMA_signal_1172, \Midori/rounds/roundResult_Reg/GEN[45].SFF/Q_708 }), .I2 ({new_AGEMA_signal_1173, \Midori/rounds/roundResult_Reg/GEN[46].SFF/Q_709 }), .I3 ({new_AGEMA_signal_1174, \Midori/rounds/roundResult_Reg/GEN[47].SFF/Q_710 }), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704]}), .O ({new_AGEMA_signal_1175, \Midori/rounds_Output [44]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[11].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1171, \Midori/rounds/roundResult_Reg/GEN[44].SFF/Q_707 }), .I1 ({new_AGEMA_signal_1172, \Midori/rounds/roundResult_Reg/GEN[45].SFF/Q_708 }), .I2 ({new_AGEMA_signal_1173, \Midori/rounds/roundResult_Reg/GEN[46].SFF/Q_709 }), .I3 ({new_AGEMA_signal_1174, \Midori/rounds/roundResult_Reg/GEN[47].SFF/Q_710 }), .clk (clk), .r ({Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .O ({new_AGEMA_signal_1176, \Midori/rounds_Output [45]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[11].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1171, \Midori/rounds/roundResult_Reg/GEN[44].SFF/Q_707 }), .I1 ({new_AGEMA_signal_1172, \Midori/rounds/roundResult_Reg/GEN[45].SFF/Q_708 }), .I2 ({new_AGEMA_signal_1173, \Midori/rounds/roundResult_Reg/GEN[46].SFF/Q_709 }), .I3 ({new_AGEMA_signal_1174, \Midori/rounds/roundResult_Reg/GEN[47].SFF/Q_710 }), .clk (clk), .r ({Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736]}), .O ({new_AGEMA_signal_1177, \Midori/rounds_Output [46]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[11].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1171, \Midori/rounds/roundResult_Reg/GEN[44].SFF/Q_707 }), .I1 ({new_AGEMA_signal_1172, \Midori/rounds/roundResult_Reg/GEN[45].SFF/Q_708 }), .I2 ({new_AGEMA_signal_1173, \Midori/rounds/roundResult_Reg/GEN[46].SFF/Q_709 }), .I3 ({new_AGEMA_signal_1174, \Midori/rounds/roundResult_Reg/GEN[47].SFF/Q_710 }), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752]}), .O ({new_AGEMA_signal_1178, \Midori/rounds_Output [47]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[12].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1179, \Midori/rounds/roundResult_Reg/GEN[48].SFF/Q_711 }), .I1 ({new_AGEMA_signal_1180, \Midori/rounds/roundResult_Reg/GEN[49].SFF/Q_712 }), .I2 ({new_AGEMA_signal_1181, \Midori/rounds/roundResult_Reg/GEN[50].SFF/Q_713 }), .I3 ({new_AGEMA_signal_1182, \Midori/rounds/roundResult_Reg/GEN[51].SFF/Q_714 }), .clk (clk), .r ({Fresh[783], Fresh[782], Fresh[781], Fresh[780], Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .O ({new_AGEMA_signal_1183, \Midori/rounds_Output [48]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[12].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1179, \Midori/rounds/roundResult_Reg/GEN[48].SFF/Q_711 }), .I1 ({new_AGEMA_signal_1180, \Midori/rounds/roundResult_Reg/GEN[49].SFF/Q_712 }), .I2 ({new_AGEMA_signal_1181, \Midori/rounds/roundResult_Reg/GEN[50].SFF/Q_713 }), .I3 ({new_AGEMA_signal_1182, \Midori/rounds/roundResult_Reg/GEN[51].SFF/Q_714 }), .clk (clk), .r ({Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784]}), .O ({new_AGEMA_signal_1184, \Midori/rounds_Output [49]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[12].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1179, \Midori/rounds/roundResult_Reg/GEN[48].SFF/Q_711 }), .I1 ({new_AGEMA_signal_1180, \Midori/rounds/roundResult_Reg/GEN[49].SFF/Q_712 }), .I2 ({new_AGEMA_signal_1181, \Midori/rounds/roundResult_Reg/GEN[50].SFF/Q_713 }), .I3 ({new_AGEMA_signal_1182, \Midori/rounds/roundResult_Reg/GEN[51].SFF/Q_714 }), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .O ({new_AGEMA_signal_1185, \Midori/rounds_Output [50]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[12].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1179, \Midori/rounds/roundResult_Reg/GEN[48].SFF/Q_711 }), .I1 ({new_AGEMA_signal_1180, \Midori/rounds/roundResult_Reg/GEN[49].SFF/Q_712 }), .I2 ({new_AGEMA_signal_1181, \Midori/rounds/roundResult_Reg/GEN[50].SFF/Q_713 }), .I3 ({new_AGEMA_signal_1182, \Midori/rounds/roundResult_Reg/GEN[51].SFF/Q_714 }), .clk (clk), .r ({Fresh[831], Fresh[830], Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .O ({new_AGEMA_signal_1186, \Midori/rounds_Output [51]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[13].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1187, \Midori/rounds/roundResult_Reg/GEN[52].SFF/Q_715 }), .I1 ({new_AGEMA_signal_1188, \Midori/rounds/roundResult_Reg/GEN[53].SFF/Q_716 }), .I2 ({new_AGEMA_signal_1189, \Midori/rounds/roundResult_Reg/GEN[54].SFF/Q_717 }), .I3 ({new_AGEMA_signal_1190, \Midori/rounds/roundResult_Reg/GEN[55].SFF/Q_718 }), .clk (clk), .r ({Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840], Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832]}), .O ({new_AGEMA_signal_1191, \Midori/rounds_Output [52]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[13].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1187, \Midori/rounds/roundResult_Reg/GEN[52].SFF/Q_715 }), .I1 ({new_AGEMA_signal_1188, \Midori/rounds/roundResult_Reg/GEN[53].SFF/Q_716 }), .I2 ({new_AGEMA_signal_1189, \Midori/rounds/roundResult_Reg/GEN[54].SFF/Q_717 }), .I3 ({new_AGEMA_signal_1190, \Midori/rounds/roundResult_Reg/GEN[55].SFF/Q_718 }), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850], Fresh[849], Fresh[848]}), .O ({new_AGEMA_signal_1192, \Midori/rounds_Output [53]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[13].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1187, \Midori/rounds/roundResult_Reg/GEN[52].SFF/Q_715 }), .I1 ({new_AGEMA_signal_1188, \Midori/rounds/roundResult_Reg/GEN[53].SFF/Q_716 }), .I2 ({new_AGEMA_signal_1189, \Midori/rounds/roundResult_Reg/GEN[54].SFF/Q_717 }), .I3 ({new_AGEMA_signal_1190, \Midori/rounds/roundResult_Reg/GEN[55].SFF/Q_718 }), .clk (clk), .r ({Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .O ({new_AGEMA_signal_1193, \Midori/rounds_Output [54]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[13].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1187, \Midori/rounds/roundResult_Reg/GEN[52].SFF/Q_715 }), .I1 ({new_AGEMA_signal_1188, \Midori/rounds/roundResult_Reg/GEN[53].SFF/Q_716 }), .I2 ({new_AGEMA_signal_1189, \Midori/rounds/roundResult_Reg/GEN[54].SFF/Q_717 }), .I3 ({new_AGEMA_signal_1190, \Midori/rounds/roundResult_Reg/GEN[55].SFF/Q_718 }), .clk (clk), .r ({Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880]}), .O ({new_AGEMA_signal_1194, \Midori/rounds_Output [55]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[14].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1195, \Midori/rounds/roundResult_Reg/GEN[56].SFF/Q_719 }), .I1 ({new_AGEMA_signal_1196, \Midori/rounds/roundResult_Reg/GEN[57].SFF/Q_720 }), .I2 ({new_AGEMA_signal_1197, \Midori/rounds/roundResult_Reg/GEN[58].SFF/Q_721 }), .I3 ({new_AGEMA_signal_1198, \Midori/rounds/roundResult_Reg/GEN[59].SFF/Q_722 }), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900], Fresh[899], Fresh[898], Fresh[897], Fresh[896]}), .O ({new_AGEMA_signal_1199, \Midori/rounds_Output [56]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[14].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1195, \Midori/rounds/roundResult_Reg/GEN[56].SFF/Q_719 }), .I1 ({new_AGEMA_signal_1196, \Midori/rounds/roundResult_Reg/GEN[57].SFF/Q_720 }), .I2 ({new_AGEMA_signal_1197, \Midori/rounds/roundResult_Reg/GEN[58].SFF/Q_721 }), .I3 ({new_AGEMA_signal_1198, \Midori/rounds/roundResult_Reg/GEN[59].SFF/Q_722 }), .clk (clk), .r ({Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .O ({new_AGEMA_signal_1200, \Midori/rounds_Output [57]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[14].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1195, \Midori/rounds/roundResult_Reg/GEN[56].SFF/Q_719 }), .I1 ({new_AGEMA_signal_1196, \Midori/rounds/roundResult_Reg/GEN[57].SFF/Q_720 }), .I2 ({new_AGEMA_signal_1197, \Midori/rounds/roundResult_Reg/GEN[58].SFF/Q_721 }), .I3 ({new_AGEMA_signal_1198, \Midori/rounds/roundResult_Reg/GEN[59].SFF/Q_722 }), .clk (clk), .r ({Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928]}), .O ({new_AGEMA_signal_1201, \Midori/rounds_Output [58]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[14].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1195, \Midori/rounds/roundResult_Reg/GEN[56].SFF/Q_719 }), .I1 ({new_AGEMA_signal_1196, \Midori/rounds/roundResult_Reg/GEN[57].SFF/Q_720 }), .I2 ({new_AGEMA_signal_1197, \Midori/rounds/roundResult_Reg/GEN[58].SFF/Q_721 }), .I3 ({new_AGEMA_signal_1198, \Midori/rounds/roundResult_Reg/GEN[59].SFF/Q_722 }), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944]}), .O ({new_AGEMA_signal_1202, \Midori/rounds_Output [59]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0EEC ) ) \Midori/rounds/sub/substition_PRINCE[15].sBox_PRINCE/y_0 ( .I0 ({new_AGEMA_signal_1203, \Midori/rounds/roundResult_Reg/GEN[60].SFF/Q_723 }), .I1 ({new_AGEMA_signal_1204, \Midori/rounds/roundResult_Reg/GEN[61].SFF/Q_724 }), .I2 ({new_AGEMA_signal_1205, \Midori/rounds/roundResult_Reg/GEN[62].SFF/Q_725 }), .I3 ({new_AGEMA_signal_1206, \Midori/rounds/roundResult_Reg/GEN[63].SFF/Q_726 }), .clk (clk), .r ({Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .O ({new_AGEMA_signal_1207, \Midori/rounds_Output [60]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA0FA ) ) \Midori/rounds/sub/substition_PRINCE[15].sBox_PRINCE/y_1 ( .I0 ({new_AGEMA_signal_1203, \Midori/rounds/roundResult_Reg/GEN[60].SFF/Q_723 }), .I1 ({new_AGEMA_signal_1204, \Midori/rounds/roundResult_Reg/GEN[61].SFF/Q_724 }), .I2 ({new_AGEMA_signal_1205, \Midori/rounds/roundResult_Reg/GEN[62].SFF/Q_725 }), .I3 ({new_AGEMA_signal_1206, \Midori/rounds/roundResult_Reg/GEN[63].SFF/Q_726 }), .clk (clk), .r ({Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976]}), .O ({new_AGEMA_signal_1208, \Midori/rounds_Output [61]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \Midori/rounds/sub/substition_PRINCE[15].sBox_PRINCE/y_2 ( .I0 ({new_AGEMA_signal_1203, \Midori/rounds/roundResult_Reg/GEN[60].SFF/Q_723 }), .I1 ({new_AGEMA_signal_1204, \Midori/rounds/roundResult_Reg/GEN[61].SFF/Q_724 }), .I2 ({new_AGEMA_signal_1205, \Midori/rounds/roundResult_Reg/GEN[62].SFF/Q_725 }), .I3 ({new_AGEMA_signal_1206, \Midori/rounds/roundResult_Reg/GEN[63].SFF/Q_726 }), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992]}), .O ({new_AGEMA_signal_1209, \Midori/rounds_Output [62]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0377 ) ) \Midori/rounds/sub/substition_PRINCE[15].sBox_PRINCE/y_3 ( .I0 ({new_AGEMA_signal_1203, \Midori/rounds/roundResult_Reg/GEN[60].SFF/Q_723 }), .I1 ({new_AGEMA_signal_1204, \Midori/rounds/roundResult_Reg/GEN[61].SFF/Q_724 }), .I2 ({new_AGEMA_signal_1205, \Midori/rounds/roundResult_Reg/GEN[62].SFF/Q_725 }), .I3 ({new_AGEMA_signal_1206, \Midori/rounds/roundResult_Reg/GEN[63].SFF/Q_726 }), .clk (clk), .r ({Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020], Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .O ({new_AGEMA_signal_1210, \Midori/rounds_Output [63]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[3].INST3 ( .I0 ({new_AGEMA_signal_1635, \Midori/rounds/mul_input [55]}), .I1 ({new_AGEMA_signal_1632, \Midori/rounds/mul_input [59]}), .I2 ({new_AGEMA_signal_1626, \Midori/rounds/mul_input [63]}), .I3 ({new_AGEMA_signal_1476, \Midori/rounds/SelectedKey [51]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1677, \Midori/rounds/mul_Result [51]}), .O6 ({new_AGEMA_signal_1678, \Midori/rounds/mul_ResultXORkey [51]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[3].INST2 ( .I0 ({new_AGEMA_signal_1638, \Midori/rounds/mul_input [51]}), .I1 ({new_AGEMA_signal_1632, \Midori/rounds/mul_input [59]}), .I2 ({new_AGEMA_signal_1626, \Midori/rounds/mul_input [63]}), .I3 ({new_AGEMA_signal_1473, \Midori/rounds/SelectedKey [55]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1679, \Midori/rounds/mul_Result [55]}), .O6 ({new_AGEMA_signal_1680, \Midori/rounds/mul_ResultXORkey [55]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[3].INST1 ( .I0 ({new_AGEMA_signal_1638, \Midori/rounds/mul_input [51]}), .I1 ({new_AGEMA_signal_1635, \Midori/rounds/mul_input [55]}), .I2 ({new_AGEMA_signal_1626, \Midori/rounds/mul_input [63]}), .I3 ({new_AGEMA_signal_1470, \Midori/rounds/SelectedKey [59]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1681, \Midori/rounds/mul_Result [59]}), .O6 ({new_AGEMA_signal_1682, \Midori/rounds/mul_ResultXORkey [59]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[3].INST0 ( .I0 ({new_AGEMA_signal_1638, \Midori/rounds/mul_input [51]}), .I1 ({new_AGEMA_signal_1635, \Midori/rounds/mul_input [55]}), .I2 ({new_AGEMA_signal_1632, \Midori/rounds/mul_input [59]}), .I3 ({new_AGEMA_signal_1467, \Midori/rounds/SelectedKey [63]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1683, \Midori/rounds/mul_Result [63]}), .O6 ({new_AGEMA_signal_1684, \Midori/rounds/mul_ResultXORkey [63]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[2].INST3 ( .I0 ({new_AGEMA_signal_1636, \Midori/rounds/mul_input [54]}), .I1 ({new_AGEMA_signal_1633, \Midori/rounds/mul_input [58]}), .I2 ({new_AGEMA_signal_1627, \Midori/rounds/mul_input [62]}), .I3 ({new_AGEMA_signal_1477, \Midori/rounds/SelectedKey [50]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1685, \Midori/rounds/mul_Result [50]}), .O6 ({new_AGEMA_signal_1686, \Midori/rounds/mul_ResultXORkey [50]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[2].INST2 ( .I0 ({new_AGEMA_signal_1639, \Midori/rounds/mul_input [50]}), .I1 ({new_AGEMA_signal_1633, \Midori/rounds/mul_input [58]}), .I2 ({new_AGEMA_signal_1627, \Midori/rounds/mul_input [62]}), .I3 ({new_AGEMA_signal_1474, \Midori/rounds/SelectedKey [54]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1687, \Midori/rounds/mul_Result [54]}), .O6 ({new_AGEMA_signal_1688, \Midori/rounds/mul_ResultXORkey [54]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[2].INST1 ( .I0 ({new_AGEMA_signal_1639, \Midori/rounds/mul_input [50]}), .I1 ({new_AGEMA_signal_1636, \Midori/rounds/mul_input [54]}), .I2 ({new_AGEMA_signal_1627, \Midori/rounds/mul_input [62]}), .I3 ({new_AGEMA_signal_1471, \Midori/rounds/SelectedKey [58]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1689, \Midori/rounds/mul_Result [58]}), .O6 ({new_AGEMA_signal_1690, \Midori/rounds/mul_ResultXORkey [58]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[2].INST0 ( .I0 ({new_AGEMA_signal_1639, \Midori/rounds/mul_input [50]}), .I1 ({new_AGEMA_signal_1636, \Midori/rounds/mul_input [54]}), .I2 ({new_AGEMA_signal_1633, \Midori/rounds/mul_input [58]}), .I3 ({new_AGEMA_signal_1468, \Midori/rounds/SelectedKey [62]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1691, \Midori/rounds/mul_Result [62]}), .O6 ({new_AGEMA_signal_1692, \Midori/rounds/mul_ResultXORkey [62]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[1].INST3 ( .I0 ({new_AGEMA_signal_1637, \Midori/rounds/mul_input [53]}), .I1 ({new_AGEMA_signal_1634, \Midori/rounds/mul_input [57]}), .I2 ({new_AGEMA_signal_1628, \Midori/rounds/mul_input [61]}), .I3 ({new_AGEMA_signal_1478, \Midori/rounds/SelectedKey [49]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1693, \Midori/rounds/mul_Result [49]}), .O6 ({new_AGEMA_signal_1694, \Midori/rounds/mul_ResultXORkey [49]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[1].INST2 ( .I0 ({new_AGEMA_signal_1640, \Midori/rounds/mul_input [49]}), .I1 ({new_AGEMA_signal_1634, \Midori/rounds/mul_input [57]}), .I2 ({new_AGEMA_signal_1628, \Midori/rounds/mul_input [61]}), .I3 ({new_AGEMA_signal_1475, \Midori/rounds/SelectedKey [53]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1695, \Midori/rounds/mul_Result [53]}), .O6 ({new_AGEMA_signal_1696, \Midori/rounds/mul_ResultXORkey [53]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[1].INST1 ( .I0 ({new_AGEMA_signal_1640, \Midori/rounds/mul_input [49]}), .I1 ({new_AGEMA_signal_1637, \Midori/rounds/mul_input [53]}), .I2 ({new_AGEMA_signal_1628, \Midori/rounds/mul_input [61]}), .I3 ({new_AGEMA_signal_1472, \Midori/rounds/SelectedKey [57]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1697, \Midori/rounds/mul_Result [57]}), .O6 ({new_AGEMA_signal_1698, \Midori/rounds/mul_ResultXORkey [57]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[1].INST0 ( .I0 ({new_AGEMA_signal_1640, \Midori/rounds/mul_input [49]}), .I1 ({new_AGEMA_signal_1637, \Midori/rounds/mul_input [53]}), .I2 ({new_AGEMA_signal_1634, \Midori/rounds/mul_input [57]}), .I3 ({new_AGEMA_signal_1469, \Midori/rounds/SelectedKey [61]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1699, \Midori/rounds/mul_Result [61]}), .O6 ({new_AGEMA_signal_1700, \Midori/rounds/mul_ResultXORkey [61]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[0].INST3 ( .I0 ({new_AGEMA_signal_1616, \Midori/rounds/mul_input [52]}), .I1 ({new_AGEMA_signal_1787, \Midori/rounds/mul_input [56]}), .I2 ({new_AGEMA_signal_1613, \Midori/rounds/mul_input [60]}), .I3 ({new_AGEMA_signal_1611, \Midori/rounds/ProcessedKey [48]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1842, \Midori/rounds/mul_Result [48]}), .O6 ({new_AGEMA_signal_1843, \Midori/rounds/mul_ResultXORkey [48]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[0].INST2 ( .I0 ({new_AGEMA_signal_1615, \Midori/rounds/mul_input [48]}), .I1 ({new_AGEMA_signal_1787, \Midori/rounds/mul_input [56]}), .I2 ({new_AGEMA_signal_1613, \Midori/rounds/mul_input [60]}), .I3 ({new_AGEMA_signal_1610, \Midori/rounds/ProcessedKey [52]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1844, \Midori/rounds/mul_Result [52]}), .O6 ({new_AGEMA_signal_1845, \Midori/rounds/mul_ResultXORkey [52]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[0].INST1 ( .I0 ({new_AGEMA_signal_1615, \Midori/rounds/mul_input [48]}), .I1 ({new_AGEMA_signal_1616, \Midori/rounds/mul_input [52]}), .I2 ({new_AGEMA_signal_1613, \Midori/rounds/mul_input [60]}), .I3 ({new_AGEMA_signal_1676, \Midori/rounds/ProcessedKey [56]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1701, \Midori/rounds/mul_Result [56]}), .O6 ({new_AGEMA_signal_1702, \Midori/rounds/mul_ResultXORkey [56]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC1/LoopGen[0].INST0 ( .I0 ({new_AGEMA_signal_1615, \Midori/rounds/mul_input [48]}), .I1 ({new_AGEMA_signal_1616, \Midori/rounds/mul_input [52]}), .I2 ({new_AGEMA_signal_1787, \Midori/rounds/mul_input [56]}), .I3 ({new_AGEMA_signal_1601, \Midori/rounds/ProcessedKey [60]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1846, \Midori/rounds/mul_Result [60]}), .O6 ({new_AGEMA_signal_1847, \Midori/rounds/mul_ResultXORkey [60]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[3].INST3 ( .I0 ({new_AGEMA_signal_1647, \Midori/rounds/mul_input [39]}), .I1 ({new_AGEMA_signal_1644, \Midori/rounds/mul_input [43]}), .I2 ({new_AGEMA_signal_1641, \Midori/rounds/mul_input [47]}), .I3 ({new_AGEMA_signal_1488, \Midori/rounds/SelectedKey [35]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1703, \Midori/rounds/mul_Result [35]}), .O6 ({new_AGEMA_signal_1704, \Midori/rounds/mul_ResultXORkey [35]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[3].INST2 ( .I0 ({new_AGEMA_signal_1650, \Midori/rounds/mul_input [35]}), .I1 ({new_AGEMA_signal_1644, \Midori/rounds/mul_input [43]}), .I2 ({new_AGEMA_signal_1641, \Midori/rounds/mul_input [47]}), .I3 ({new_AGEMA_signal_1485, \Midori/rounds/SelectedKey [39]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1705, \Midori/rounds/mul_Result [39]}), .O6 ({new_AGEMA_signal_1706, \Midori/rounds/mul_ResultXORkey [39]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[3].INST1 ( .I0 ({new_AGEMA_signal_1650, \Midori/rounds/mul_input [35]}), .I1 ({new_AGEMA_signal_1647, \Midori/rounds/mul_input [39]}), .I2 ({new_AGEMA_signal_1641, \Midori/rounds/mul_input [47]}), .I3 ({new_AGEMA_signal_1482, \Midori/rounds/SelectedKey [43]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1707, \Midori/rounds/mul_Result [43]}), .O6 ({new_AGEMA_signal_1708, \Midori/rounds/mul_ResultXORkey [43]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[3].INST0 ( .I0 ({new_AGEMA_signal_1650, \Midori/rounds/mul_input [35]}), .I1 ({new_AGEMA_signal_1647, \Midori/rounds/mul_input [39]}), .I2 ({new_AGEMA_signal_1644, \Midori/rounds/mul_input [43]}), .I3 ({new_AGEMA_signal_1479, \Midori/rounds/SelectedKey [47]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1709, \Midori/rounds/mul_Result [47]}), .O6 ({new_AGEMA_signal_1710, \Midori/rounds/mul_ResultXORkey [47]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[2].INST3 ( .I0 ({new_AGEMA_signal_1648, \Midori/rounds/mul_input [38]}), .I1 ({new_AGEMA_signal_1645, \Midori/rounds/mul_input [42]}), .I2 ({new_AGEMA_signal_1642, \Midori/rounds/mul_input [46]}), .I3 ({new_AGEMA_signal_1489, \Midori/rounds/SelectedKey [34]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1711, \Midori/rounds/mul_Result [34]}), .O6 ({new_AGEMA_signal_1712, \Midori/rounds/mul_ResultXORkey [34]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[2].INST2 ( .I0 ({new_AGEMA_signal_1651, \Midori/rounds/mul_input [34]}), .I1 ({new_AGEMA_signal_1645, \Midori/rounds/mul_input [42]}), .I2 ({new_AGEMA_signal_1642, \Midori/rounds/mul_input [46]}), .I3 ({new_AGEMA_signal_1486, \Midori/rounds/SelectedKey [38]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1713, \Midori/rounds/mul_Result [38]}), .O6 ({new_AGEMA_signal_1714, \Midori/rounds/mul_ResultXORkey [38]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[2].INST1 ( .I0 ({new_AGEMA_signal_1651, \Midori/rounds/mul_input [34]}), .I1 ({new_AGEMA_signal_1648, \Midori/rounds/mul_input [38]}), .I2 ({new_AGEMA_signal_1642, \Midori/rounds/mul_input [46]}), .I3 ({new_AGEMA_signal_1483, \Midori/rounds/SelectedKey [42]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1715, \Midori/rounds/mul_Result [42]}), .O6 ({new_AGEMA_signal_1716, \Midori/rounds/mul_ResultXORkey [42]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[2].INST0 ( .I0 ({new_AGEMA_signal_1651, \Midori/rounds/mul_input [34]}), .I1 ({new_AGEMA_signal_1648, \Midori/rounds/mul_input [38]}), .I2 ({new_AGEMA_signal_1645, \Midori/rounds/mul_input [42]}), .I3 ({new_AGEMA_signal_1480, \Midori/rounds/SelectedKey [46]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1717, \Midori/rounds/mul_Result [46]}), .O6 ({new_AGEMA_signal_1718, \Midori/rounds/mul_ResultXORkey [46]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[1].INST3 ( .I0 ({new_AGEMA_signal_1649, \Midori/rounds/mul_input [37]}), .I1 ({new_AGEMA_signal_1646, \Midori/rounds/mul_input [41]}), .I2 ({new_AGEMA_signal_1643, \Midori/rounds/mul_input [45]}), .I3 ({new_AGEMA_signal_1490, \Midori/rounds/SelectedKey [33]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1719, \Midori/rounds/mul_Result [33]}), .O6 ({new_AGEMA_signal_1720, \Midori/rounds/mul_ResultXORkey [33]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[1].INST2 ( .I0 ({new_AGEMA_signal_1652, \Midori/rounds/mul_input [33]}), .I1 ({new_AGEMA_signal_1646, \Midori/rounds/mul_input [41]}), .I2 ({new_AGEMA_signal_1643, \Midori/rounds/mul_input [45]}), .I3 ({new_AGEMA_signal_1487, \Midori/rounds/SelectedKey [37]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1721, \Midori/rounds/mul_Result [37]}), .O6 ({new_AGEMA_signal_1722, \Midori/rounds/mul_ResultXORkey [37]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[1].INST1 ( .I0 ({new_AGEMA_signal_1652, \Midori/rounds/mul_input [33]}), .I1 ({new_AGEMA_signal_1649, \Midori/rounds/mul_input [37]}), .I2 ({new_AGEMA_signal_1643, \Midori/rounds/mul_input [45]}), .I3 ({new_AGEMA_signal_1484, \Midori/rounds/SelectedKey [41]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1723, \Midori/rounds/mul_Result [41]}), .O6 ({new_AGEMA_signal_1724, \Midori/rounds/mul_ResultXORkey [41]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[1].INST0 ( .I0 ({new_AGEMA_signal_1652, \Midori/rounds/mul_input [33]}), .I1 ({new_AGEMA_signal_1649, \Midori/rounds/mul_input [37]}), .I2 ({new_AGEMA_signal_1646, \Midori/rounds/mul_input [41]}), .I3 ({new_AGEMA_signal_1481, \Midori/rounds/SelectedKey [45]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1725, \Midori/rounds/mul_Result [45]}), .O6 ({new_AGEMA_signal_1726, \Midori/rounds/mul_ResultXORkey [45]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[0].INST3 ( .I0 ({new_AGEMA_signal_1618, \Midori/rounds/mul_input [36]}), .I1 ({new_AGEMA_signal_1625, \Midori/rounds/mul_input [40]}), .I2 ({new_AGEMA_signal_1617, \Midori/rounds/mul_input [44]}), .I3 ({new_AGEMA_signal_1604, \Midori/rounds/ProcessedKey [32]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1727, \Midori/rounds/mul_Result [32]}), .O6 ({new_AGEMA_signal_1728, \Midori/rounds/mul_ResultXORkey [32]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[0].INST2 ( .I0 ({new_AGEMA_signal_1619, \Midori/rounds/mul_input [32]}), .I1 ({new_AGEMA_signal_1625, \Midori/rounds/mul_input [40]}), .I2 ({new_AGEMA_signal_1617, \Midori/rounds/mul_input [44]}), .I3 ({new_AGEMA_signal_1609, \Midori/rounds/ProcessedKey [36]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1729, \Midori/rounds/mul_Result [36]}), .O6 ({new_AGEMA_signal_1730, \Midori/rounds/mul_ResultXORkey [36]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[0].INST1 ( .I0 ({new_AGEMA_signal_1619, \Midori/rounds/mul_input [32]}), .I1 ({new_AGEMA_signal_1618, \Midori/rounds/mul_input [36]}), .I2 ({new_AGEMA_signal_1617, \Midori/rounds/mul_input [44]}), .I3 ({new_AGEMA_signal_1612, \Midori/rounds/ProcessedKey [40]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1731, \Midori/rounds/mul_Result [40]}), .O6 ({new_AGEMA_signal_1732, \Midori/rounds/mul_ResultXORkey [40]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC2/LoopGen[0].INST0 ( .I0 ({new_AGEMA_signal_1619, \Midori/rounds/mul_input [32]}), .I1 ({new_AGEMA_signal_1618, \Midori/rounds/mul_input [36]}), .I2 ({new_AGEMA_signal_1625, \Midori/rounds/mul_input [40]}), .I3 ({new_AGEMA_signal_1603, \Midori/rounds/ProcessedKey [44]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1733, \Midori/rounds/mul_Result [44]}), .O6 ({new_AGEMA_signal_1734, \Midori/rounds/mul_ResultXORkey [44]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[3].INST3 ( .I0 ({new_AGEMA_signal_1659, \Midori/rounds/mul_input [23]}), .I1 ({new_AGEMA_signal_1656, \Midori/rounds/mul_input [27]}), .I2 ({new_AGEMA_signal_1653, \Midori/rounds/mul_input [31]}), .I3 ({new_AGEMA_signal_1500, \Midori/rounds/SelectedKey [19]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1735, \Midori/rounds/mul_Result [19]}), .O6 ({new_AGEMA_signal_1736, \Midori/rounds/mul_ResultXORkey [19]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[3].INST2 ( .I0 ({new_AGEMA_signal_1662, \Midori/rounds/mul_input [19]}), .I1 ({new_AGEMA_signal_1656, \Midori/rounds/mul_input [27]}), .I2 ({new_AGEMA_signal_1653, \Midori/rounds/mul_input [31]}), .I3 ({new_AGEMA_signal_1497, \Midori/rounds/SelectedKey [23]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1737, \Midori/rounds/mul_Result [23]}), .O6 ({new_AGEMA_signal_1738, \Midori/rounds/mul_ResultXORkey [23]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[3].INST1 ( .I0 ({new_AGEMA_signal_1662, \Midori/rounds/mul_input [19]}), .I1 ({new_AGEMA_signal_1659, \Midori/rounds/mul_input [23]}), .I2 ({new_AGEMA_signal_1653, \Midori/rounds/mul_input [31]}), .I3 ({new_AGEMA_signal_1494, \Midori/rounds/SelectedKey [27]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1739, \Midori/rounds/mul_Result [27]}), .O6 ({new_AGEMA_signal_1740, \Midori/rounds/mul_ResultXORkey [27]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[3].INST0 ( .I0 ({new_AGEMA_signal_1662, \Midori/rounds/mul_input [19]}), .I1 ({new_AGEMA_signal_1659, \Midori/rounds/mul_input [23]}), .I2 ({new_AGEMA_signal_1656, \Midori/rounds/mul_input [27]}), .I3 ({new_AGEMA_signal_1491, \Midori/rounds/SelectedKey [31]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1741, \Midori/rounds/mul_Result [31]}), .O6 ({new_AGEMA_signal_1742, \Midori/rounds/mul_ResultXORkey [31]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[2].INST3 ( .I0 ({new_AGEMA_signal_1660, \Midori/rounds/mul_input [22]}), .I1 ({new_AGEMA_signal_1657, \Midori/rounds/mul_input [26]}), .I2 ({new_AGEMA_signal_1654, \Midori/rounds/mul_input [30]}), .I3 ({new_AGEMA_signal_1501, \Midori/rounds/SelectedKey [18]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1743, \Midori/rounds/mul_Result [18]}), .O6 ({new_AGEMA_signal_1744, \Midori/rounds/mul_ResultXORkey [18]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[2].INST2 ( .I0 ({new_AGEMA_signal_1663, \Midori/rounds/mul_input [18]}), .I1 ({new_AGEMA_signal_1657, \Midori/rounds/mul_input [26]}), .I2 ({new_AGEMA_signal_1654, \Midori/rounds/mul_input [30]}), .I3 ({new_AGEMA_signal_1498, \Midori/rounds/SelectedKey [22]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1745, \Midori/rounds/mul_Result [22]}), .O6 ({new_AGEMA_signal_1746, \Midori/rounds/mul_ResultXORkey [22]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[2].INST1 ( .I0 ({new_AGEMA_signal_1663, \Midori/rounds/mul_input [18]}), .I1 ({new_AGEMA_signal_1660, \Midori/rounds/mul_input [22]}), .I2 ({new_AGEMA_signal_1654, \Midori/rounds/mul_input [30]}), .I3 ({new_AGEMA_signal_1495, \Midori/rounds/SelectedKey [26]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1747, \Midori/rounds/mul_Result [26]}), .O6 ({new_AGEMA_signal_1748, \Midori/rounds/mul_ResultXORkey [26]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[2].INST0 ( .I0 ({new_AGEMA_signal_1663, \Midori/rounds/mul_input [18]}), .I1 ({new_AGEMA_signal_1660, \Midori/rounds/mul_input [22]}), .I2 ({new_AGEMA_signal_1657, \Midori/rounds/mul_input [26]}), .I3 ({new_AGEMA_signal_1492, \Midori/rounds/SelectedKey [30]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1749, \Midori/rounds/mul_Result [30]}), .O6 ({new_AGEMA_signal_1750, \Midori/rounds/mul_ResultXORkey [30]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[1].INST3 ( .I0 ({new_AGEMA_signal_1661, \Midori/rounds/mul_input [21]}), .I1 ({new_AGEMA_signal_1658, \Midori/rounds/mul_input [25]}), .I2 ({new_AGEMA_signal_1655, \Midori/rounds/mul_input [29]}), .I3 ({new_AGEMA_signal_1502, \Midori/rounds/SelectedKey [17]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1751, \Midori/rounds/mul_Result [17]}), .O6 ({new_AGEMA_signal_1752, \Midori/rounds/mul_ResultXORkey [17]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[1].INST2 ( .I0 ({new_AGEMA_signal_1664, \Midori/rounds/mul_input [17]}), .I1 ({new_AGEMA_signal_1658, \Midori/rounds/mul_input [25]}), .I2 ({new_AGEMA_signal_1655, \Midori/rounds/mul_input [29]}), .I3 ({new_AGEMA_signal_1499, \Midori/rounds/SelectedKey [21]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1753, \Midori/rounds/mul_Result [21]}), .O6 ({new_AGEMA_signal_1754, \Midori/rounds/mul_ResultXORkey [21]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[1].INST1 ( .I0 ({new_AGEMA_signal_1664, \Midori/rounds/mul_input [17]}), .I1 ({new_AGEMA_signal_1661, \Midori/rounds/mul_input [21]}), .I2 ({new_AGEMA_signal_1655, \Midori/rounds/mul_input [29]}), .I3 ({new_AGEMA_signal_1496, \Midori/rounds/SelectedKey [25]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1755, \Midori/rounds/mul_Result [25]}), .O6 ({new_AGEMA_signal_1756, \Midori/rounds/mul_ResultXORkey [25]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[1].INST0 ( .I0 ({new_AGEMA_signal_1664, \Midori/rounds/mul_input [17]}), .I1 ({new_AGEMA_signal_1661, \Midori/rounds/mul_input [21]}), .I2 ({new_AGEMA_signal_1658, \Midori/rounds/mul_input [25]}), .I3 ({new_AGEMA_signal_1493, \Midori/rounds/SelectedKey [29]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1757, \Midori/rounds/mul_Result [29]}), .O6 ({new_AGEMA_signal_1758, \Midori/rounds/mul_ResultXORkey [29]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[0].INST3 ( .I0 ({new_AGEMA_signal_1622, \Midori/rounds/mul_input [20]}), .I1 ({new_AGEMA_signal_1621, \Midori/rounds/mul_input [24]}), .I2 ({new_AGEMA_signal_1620, \Midori/rounds/mul_input [28]}), .I3 ({new_AGEMA_signal_1675, \Midori/rounds/ProcessedKey [16]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1759, \Midori/rounds/mul_Result [16]}), .O6 ({new_AGEMA_signal_1760, \Midori/rounds/mul_ResultXORkey [16]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[0].INST2 ( .I0 ({new_AGEMA_signal_1788, \Midori/rounds/mul_input [16]}), .I1 ({new_AGEMA_signal_1621, \Midori/rounds/mul_input [24]}), .I2 ({new_AGEMA_signal_1620, \Midori/rounds/mul_input [28]}), .I3 ({new_AGEMA_signal_1607, \Midori/rounds/ProcessedKey [20]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1848, \Midori/rounds/mul_Result [20]}), .O6 ({new_AGEMA_signal_1849, \Midori/rounds/mul_ResultXORkey [20]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[0].INST1 ( .I0 ({new_AGEMA_signal_1788, \Midori/rounds/mul_input [16]}), .I1 ({new_AGEMA_signal_1622, \Midori/rounds/mul_input [20]}), .I2 ({new_AGEMA_signal_1620, \Midori/rounds/mul_input [28]}), .I3 ({new_AGEMA_signal_1606, \Midori/rounds/ProcessedKey [24]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1850, \Midori/rounds/mul_Result [24]}), .O6 ({new_AGEMA_signal_1851, \Midori/rounds/mul_ResultXORkey [24]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC3/LoopGen[0].INST0 ( .I0 ({new_AGEMA_signal_1788, \Midori/rounds/mul_input [16]}), .I1 ({new_AGEMA_signal_1622, \Midori/rounds/mul_input [20]}), .I2 ({new_AGEMA_signal_1621, \Midori/rounds/mul_input [24]}), .I3 ({new_AGEMA_signal_1605, \Midori/rounds/ProcessedKey [28]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1852, \Midori/rounds/mul_Result [28]}), .O6 ({new_AGEMA_signal_1853, \Midori/rounds/mul_ResultXORkey [28]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[3].INST3 ( .I0 ({new_AGEMA_signal_1668, \Midori/rounds/mul_input [7]}), .I1 ({new_AGEMA_signal_1629, \Midori/rounds/mul_input [11]}), .I2 ({new_AGEMA_signal_1665, \Midori/rounds/mul_input [15]}), .I3 ({new_AGEMA_signal_1512, \Midori/rounds/SelectedKey [3]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1761, \Midori/rounds/mul_Result [3]}), .O6 ({new_AGEMA_signal_1762, \Midori/rounds/mul_ResultXORkey [3]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[3].INST2 ( .I0 ({new_AGEMA_signal_1671, \Midori/rounds/mul_input [3]}), .I1 ({new_AGEMA_signal_1629, \Midori/rounds/mul_input [11]}), .I2 ({new_AGEMA_signal_1665, \Midori/rounds/mul_input [15]}), .I3 ({new_AGEMA_signal_1509, \Midori/rounds/SelectedKey [7]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1763, \Midori/rounds/mul_Result [7]}), .O6 ({new_AGEMA_signal_1764, \Midori/rounds/mul_ResultXORkey [7]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[3].INST1 ( .I0 ({new_AGEMA_signal_1671, \Midori/rounds/mul_input [3]}), .I1 ({new_AGEMA_signal_1668, \Midori/rounds/mul_input [7]}), .I2 ({new_AGEMA_signal_1665, \Midori/rounds/mul_input [15]}), .I3 ({new_AGEMA_signal_1506, \Midori/rounds/SelectedKey [11]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1765, \Midori/rounds/mul_Result [11]}), .O6 ({new_AGEMA_signal_1766, \Midori/rounds/mul_ResultXORkey [11]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[3].INST0 ( .I0 ({new_AGEMA_signal_1671, \Midori/rounds/mul_input [3]}), .I1 ({new_AGEMA_signal_1668, \Midori/rounds/mul_input [7]}), .I2 ({new_AGEMA_signal_1629, \Midori/rounds/mul_input [11]}), .I3 ({new_AGEMA_signal_1503, \Midori/rounds/SelectedKey [15]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1767, \Midori/rounds/mul_Result [15]}), .O6 ({new_AGEMA_signal_1768, \Midori/rounds/mul_ResultXORkey [15]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[2].INST3 ( .I0 ({new_AGEMA_signal_1669, \Midori/rounds/mul_input [6]}), .I1 ({new_AGEMA_signal_1630, \Midori/rounds/mul_input [10]}), .I2 ({new_AGEMA_signal_1666, \Midori/rounds/mul_input [14]}), .I3 ({new_AGEMA_signal_1513, \Midori/rounds/SelectedKey [2]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1769, \Midori/rounds/mul_Result [2]}), .O6 ({new_AGEMA_signal_1770, \Midori/rounds/mul_ResultXORkey [2]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[2].INST2 ( .I0 ({new_AGEMA_signal_1672, \Midori/rounds/mul_input [2]}), .I1 ({new_AGEMA_signal_1630, \Midori/rounds/mul_input [10]}), .I2 ({new_AGEMA_signal_1666, \Midori/rounds/mul_input [14]}), .I3 ({new_AGEMA_signal_1510, \Midori/rounds/SelectedKey [6]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1771, \Midori/rounds/mul_Result [6]}), .O6 ({new_AGEMA_signal_1772, \Midori/rounds/mul_ResultXORkey [6]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[2].INST1 ( .I0 ({new_AGEMA_signal_1672, \Midori/rounds/mul_input [2]}), .I1 ({new_AGEMA_signal_1669, \Midori/rounds/mul_input [6]}), .I2 ({new_AGEMA_signal_1666, \Midori/rounds/mul_input [14]}), .I3 ({new_AGEMA_signal_1507, \Midori/rounds/SelectedKey [10]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1773, \Midori/rounds/mul_Result [10]}), .O6 ({new_AGEMA_signal_1774, \Midori/rounds/mul_ResultXORkey [10]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[2].INST0 ( .I0 ({new_AGEMA_signal_1672, \Midori/rounds/mul_input [2]}), .I1 ({new_AGEMA_signal_1669, \Midori/rounds/mul_input [6]}), .I2 ({new_AGEMA_signal_1630, \Midori/rounds/mul_input [10]}), .I3 ({new_AGEMA_signal_1504, \Midori/rounds/SelectedKey [14]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1775, \Midori/rounds/mul_Result [14]}), .O6 ({new_AGEMA_signal_1776, \Midori/rounds/mul_ResultXORkey [14]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[1].INST3 ( .I0 ({new_AGEMA_signal_1670, \Midori/rounds/mul_input [5]}), .I1 ({new_AGEMA_signal_1631, \Midori/rounds/mul_input [9]}), .I2 ({new_AGEMA_signal_1667, \Midori/rounds/mul_input [13]}), .I3 ({new_AGEMA_signal_1514, \Midori/rounds/SelectedKey [1]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1777, \Midori/rounds/mul_Result [1]}), .O6 ({new_AGEMA_signal_1778, \Midori/rounds/mul_ResultXORkey [1]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[1].INST2 ( .I0 ({new_AGEMA_signal_1673, \Midori/rounds/mul_input [1]}), .I1 ({new_AGEMA_signal_1631, \Midori/rounds/mul_input [9]}), .I2 ({new_AGEMA_signal_1667, \Midori/rounds/mul_input [13]}), .I3 ({new_AGEMA_signal_1511, \Midori/rounds/SelectedKey [5]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1779, \Midori/rounds/mul_Result [5]}), .O6 ({new_AGEMA_signal_1780, \Midori/rounds/mul_ResultXORkey [5]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[1].INST1 ( .I0 ({new_AGEMA_signal_1673, \Midori/rounds/mul_input [1]}), .I1 ({new_AGEMA_signal_1670, \Midori/rounds/mul_input [5]}), .I2 ({new_AGEMA_signal_1667, \Midori/rounds/mul_input [13]}), .I3 ({new_AGEMA_signal_1508, \Midori/rounds/SelectedKey [9]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1781, \Midori/rounds/mul_Result [9]}), .O6 ({new_AGEMA_signal_1782, \Midori/rounds/mul_ResultXORkey [9]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[1].INST0 ( .I0 ({new_AGEMA_signal_1673, \Midori/rounds/mul_input [1]}), .I1 ({new_AGEMA_signal_1670, \Midori/rounds/mul_input [5]}), .I2 ({new_AGEMA_signal_1631, \Midori/rounds/mul_input [9]}), .I3 ({new_AGEMA_signal_1505, \Midori/rounds/SelectedKey [13]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1783, \Midori/rounds/mul_Result [13]}), .O6 ({new_AGEMA_signal_1784, \Midori/rounds/mul_ResultXORkey [13]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[0].INST3 ( .I0 ({new_AGEMA_signal_1624, \Midori/rounds/mul_input [4]}), .I1 ({new_AGEMA_signal_1614, \Midori/rounds/mul_input [8]}), .I2 ({new_AGEMA_signal_1623, \Midori/rounds/mul_input [12]}), .I3 ({new_AGEMA_signal_1674, \Midori/rounds/ProcessedKey [0]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1785, \Midori/rounds/mul_Result [0]}), .O6 ({new_AGEMA_signal_1786, \Midori/rounds/mul_ResultXORkey [0]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[0].INST2 ( .I0 ({new_AGEMA_signal_1789, \Midori/rounds/mul_input [0]}), .I1 ({new_AGEMA_signal_1614, \Midori/rounds/mul_input [8]}), .I2 ({new_AGEMA_signal_1623, \Midori/rounds/mul_input [12]}), .I3 ({new_AGEMA_signal_1602, \Midori/rounds/ProcessedKey [4]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1854, \Midori/rounds/mul_Result [4]}), .O6 ({new_AGEMA_signal_1855, \Midori/rounds/mul_ResultXORkey [4]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[0].INST1 ( .I0 ({new_AGEMA_signal_1789, \Midori/rounds/mul_input [0]}), .I1 ({new_AGEMA_signal_1624, \Midori/rounds/mul_input [4]}), .I2 ({new_AGEMA_signal_1623, \Midori/rounds/mul_input [12]}), .I3 ({new_AGEMA_signal_1600, \Midori/rounds/ProcessedKey [8]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1856, \Midori/rounds/mul_Result [8]}), .O6 ({new_AGEMA_signal_1857, \Midori/rounds/mul_ResultXORkey [8]}) ) ;
    LUT6_2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h0000699600009696 ) , .MASK ( 6'b110000 ), .INIT2 ( 64'h0000699600009696 ) ) \Midori/rounds/mul/MC4/LoopGen[0].INST0 ( .I0 ({new_AGEMA_signal_1789, \Midori/rounds/mul_input [0]}), .I1 ({new_AGEMA_signal_1624, \Midori/rounds/mul_input [4]}), .I2 ({new_AGEMA_signal_1614, \Midori/rounds/mul_input [8]}), .I3 ({new_AGEMA_signal_1608, \Midori/rounds/ProcessedKey [12]}), .I4 ({1'b0, 1'b0}), .I5 (1'b1), .O5 ({new_AGEMA_signal_1858, \Midori/rounds/mul_Result [12]}), .O6 ({new_AGEMA_signal_1859, \Midori/rounds/mul_ResultXORkey [12]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<9>1 ( .I0 ({key_s1[73], key_s0[73]}), .I1 ({new_AGEMA_signal_1104, \Midori/rounds_Output [9]}), .I2 ({key_s1[9], key_s0[9]}), .O ({output_1_s1[9], output_1_s0[9]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<8>1 ( .I0 ({key_s1[72], key_s0[72]}), .I1 ({new_AGEMA_signal_1103, \Midori/rounds_Output [8]}), .I2 ({key_s1[8], key_s0[8]}), .O ({output_1_s1[8], output_1_s0[8]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<7>1 ( .I0 ({key_s1[71], key_s0[71]}), .I1 ({new_AGEMA_signal_1098, \Midori/rounds_Output [7]}), .I2 ({key_s1[7], key_s0[7]}), .O ({output_1_s1[7], output_1_s0[7]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<63>1 ( .I0 ({new_AGEMA_signal_1210, \Midori/rounds_Output [63]}), .I1 ({key_s1[63], key_s0[63]}), .I2 ({key_s1[127], key_s0[127]}), .O ({output_1_s1[63], output_1_s0[63]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<62>1 ( .I0 ({new_AGEMA_signal_1209, \Midori/rounds_Output [62]}), .I1 ({key_s1[62], key_s0[62]}), .I2 ({key_s1[126], key_s0[126]}), .O ({output_1_s1[62], output_1_s0[62]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<61>1 ( .I0 ({new_AGEMA_signal_1208, \Midori/rounds_Output [61]}), .I1 ({key_s1[61], key_s0[61]}), .I2 ({key_s1[125], key_s0[125]}), .O ({output_1_s1[61], output_1_s0[61]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<60>1 ( .I0 ({new_AGEMA_signal_1207, \Midori/rounds_Output [60]}), .I1 ({key_s1[60], key_s0[60]}), .I2 ({key_s1[124], key_s0[124]}), .O ({output_1_s1[60], output_1_s0[60]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<6>1 ( .I0 ({key_s1[70], key_s0[70]}), .I1 ({new_AGEMA_signal_1097, \Midori/rounds_Output [6]}), .I2 ({key_s1[6], key_s0[6]}), .O ({output_1_s1[6], output_1_s0[6]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<59>1 ( .I0 ({key_s1[123], key_s0[123]}), .I1 ({new_AGEMA_signal_1202, \Midori/rounds_Output [59]}), .I2 ({key_s1[59], key_s0[59]}), .O ({output_1_s1[59], output_1_s0[59]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<58>1 ( .I0 ({key_s1[122], key_s0[122]}), .I1 ({new_AGEMA_signal_1201, \Midori/rounds_Output [58]}), .I2 ({key_s1[58], key_s0[58]}), .O ({output_1_s1[58], output_1_s0[58]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<57>1 ( .I0 ({key_s1[121], key_s0[121]}), .I1 ({new_AGEMA_signal_1200, \Midori/rounds_Output [57]}), .I2 ({key_s1[57], key_s0[57]}), .O ({output_1_s1[57], output_1_s0[57]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<56>1 ( .I0 ({key_s1[120], key_s0[120]}), .I1 ({new_AGEMA_signal_1199, \Midori/rounds_Output [56]}), .I2 ({key_s1[56], key_s0[56]}), .O ({output_1_s1[56], output_1_s0[56]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<55>1 ( .I0 ({new_AGEMA_signal_1194, \Midori/rounds_Output [55]}), .I1 ({key_s1[55], key_s0[55]}), .I2 ({key_s1[119], key_s0[119]}), .O ({output_1_s1[55], output_1_s0[55]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<54>1 ( .I0 ({new_AGEMA_signal_1193, \Midori/rounds_Output [54]}), .I1 ({key_s1[54], key_s0[54]}), .I2 ({key_s1[118], key_s0[118]}), .O ({output_1_s1[54], output_1_s0[54]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<53>1 ( .I0 ({new_AGEMA_signal_1192, \Midori/rounds_Output [53]}), .I1 ({key_s1[53], key_s0[53]}), .I2 ({key_s1[117], key_s0[117]}), .O ({output_1_s1[53], output_1_s0[53]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<52>1 ( .I0 ({new_AGEMA_signal_1191, \Midori/rounds_Output [52]}), .I1 ({key_s1[52], key_s0[52]}), .I2 ({key_s1[116], key_s0[116]}), .O ({output_1_s1[52], output_1_s0[52]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<51>1 ( .I0 ({new_AGEMA_signal_1186, \Midori/rounds_Output [51]}), .I1 ({key_s1[51], key_s0[51]}), .I2 ({key_s1[115], key_s0[115]}), .O ({output_1_s1[51], output_1_s0[51]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<50>1 ( .I0 ({new_AGEMA_signal_1185, \Midori/rounds_Output [50]}), .I1 ({key_s1[50], key_s0[50]}), .I2 ({key_s1[114], key_s0[114]}), .O ({output_1_s1[50], output_1_s0[50]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<5>1 ( .I0 ({new_AGEMA_signal_1096, \Midori/rounds_Output [5]}), .I1 ({key_s1[5], key_s0[5]}), .I2 ({key_s1[69], key_s0[69]}), .O ({output_1_s1[5], output_1_s0[5]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<49>1 ( .I0 ({key_s1[113], key_s0[113]}), .I1 ({new_AGEMA_signal_1184, \Midori/rounds_Output [49]}), .I2 ({key_s1[49], key_s0[49]}), .O ({output_1_s1[49], output_1_s0[49]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<48>1 ( .I0 ({key_s1[112], key_s0[112]}), .I1 ({new_AGEMA_signal_1183, \Midori/rounds_Output [48]}), .I2 ({key_s1[48], key_s0[48]}), .O ({output_1_s1[48], output_1_s0[48]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<47>1 ( .I0 ({key_s1[111], key_s0[111]}), .I1 ({new_AGEMA_signal_1178, \Midori/rounds_Output [47]}), .I2 ({key_s1[47], key_s0[47]}), .O ({output_1_s1[47], output_1_s0[47]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<46>1 ( .I0 ({key_s1[110], key_s0[110]}), .I1 ({new_AGEMA_signal_1177, \Midori/rounds_Output [46]}), .I2 ({key_s1[46], key_s0[46]}), .O ({output_1_s1[46], output_1_s0[46]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<45>1 ( .I0 ({new_AGEMA_signal_1176, \Midori/rounds_Output [45]}), .I1 ({key_s1[45], key_s0[45]}), .I2 ({key_s1[109], key_s0[109]}), .O ({output_1_s1[45], output_1_s0[45]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<44>1 ( .I0 ({new_AGEMA_signal_1175, \Midori/rounds_Output [44]}), .I1 ({key_s1[44], key_s0[44]}), .I2 ({key_s1[108], key_s0[108]}), .O ({output_1_s1[44], output_1_s0[44]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<43>1 ( .I0 ({new_AGEMA_signal_1170, \Midori/rounds_Output [43]}), .I1 ({key_s1[43], key_s0[43]}), .I2 ({key_s1[107], key_s0[107]}), .O ({output_1_s1[43], output_1_s0[43]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<42>1 ( .I0 ({new_AGEMA_signal_1169, \Midori/rounds_Output [42]}), .I1 ({key_s1[42], key_s0[42]}), .I2 ({key_s1[106], key_s0[106]}), .O ({output_1_s1[42], output_1_s0[42]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<41>1 ( .I0 ({new_AGEMA_signal_1168, \Midori/rounds_Output [41]}), .I1 ({key_s1[41], key_s0[41]}), .I2 ({key_s1[105], key_s0[105]}), .O ({output_1_s1[41], output_1_s0[41]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<40>1 ( .I0 ({new_AGEMA_signal_1167, \Midori/rounds_Output [40]}), .I1 ({key_s1[40], key_s0[40]}), .I2 ({key_s1[104], key_s0[104]}), .O ({output_1_s1[40], output_1_s0[40]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<4>1 ( .I0 ({new_AGEMA_signal_1095, \Midori/rounds_Output [4]}), .I1 ({key_s1[4], key_s0[4]}), .I2 ({key_s1[68], key_s0[68]}), .O ({output_1_s1[4], output_1_s0[4]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<39>1 ( .I0 ({key_s1[103], key_s0[103]}), .I1 ({new_AGEMA_signal_1162, \Midori/rounds_Output [39]}), .I2 ({key_s1[39], key_s0[39]}), .O ({output_1_s1[39], output_1_s0[39]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<38>1 ( .I0 ({key_s1[102], key_s0[102]}), .I1 ({new_AGEMA_signal_1161, \Midori/rounds_Output [38]}), .I2 ({key_s1[38], key_s0[38]}), .O ({output_1_s1[38], output_1_s0[38]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<37>1 ( .I0 ({key_s1[101], key_s0[101]}), .I1 ({new_AGEMA_signal_1160, \Midori/rounds_Output [37]}), .I2 ({key_s1[37], key_s0[37]}), .O ({output_1_s1[37], output_1_s0[37]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<36>1 ( .I0 ({key_s1[100], key_s0[100]}), .I1 ({new_AGEMA_signal_1159, \Midori/rounds_Output [36]}), .I2 ({key_s1[36], key_s0[36]}), .O ({output_1_s1[36], output_1_s0[36]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<35>1 ( .I0 ({new_AGEMA_signal_1154, \Midori/rounds_Output [35]}), .I1 ({key_s1[35], key_s0[35]}), .I2 ({key_s1[99], key_s0[99]}), .O ({output_1_s1[35], output_1_s0[35]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<34>1 ( .I0 ({new_AGEMA_signal_1153, \Midori/rounds_Output [34]}), .I1 ({key_s1[34], key_s0[34]}), .I2 ({key_s1[98], key_s0[98]}), .O ({output_1_s1[34], output_1_s0[34]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<33>1 ( .I0 ({new_AGEMA_signal_1152, \Midori/rounds_Output [33]}), .I1 ({key_s1[33], key_s0[33]}), .I2 ({key_s1[97], key_s0[97]}), .O ({output_1_s1[33], output_1_s0[33]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<32>1 ( .I0 ({new_AGEMA_signal_1151, \Midori/rounds_Output [32]}), .I1 ({key_s1[32], key_s0[32]}), .I2 ({key_s1[96], key_s0[96]}), .O ({output_1_s1[32], output_1_s0[32]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<31>1 ( .I0 ({new_AGEMA_signal_1146, \Midori/rounds_Output [31]}), .I1 ({key_s1[31], key_s0[31]}), .I2 ({key_s1[95], key_s0[95]}), .O ({output_1_s1[31], output_1_s0[31]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<30>1 ( .I0 ({new_AGEMA_signal_1145, \Midori/rounds_Output [30]}), .I1 ({key_s1[30], key_s0[30]}), .I2 ({key_s1[94], key_s0[94]}), .O ({output_1_s1[30], output_1_s0[30]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<3>1 ( .I0 ({new_AGEMA_signal_1090, \Midori/rounds_Output [3]}), .I1 ({key_s1[3], key_s0[3]}), .I2 ({key_s1[67], key_s0[67]}), .O ({output_1_s1[3], output_1_s0[3]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<29>1 ( .I0 ({key_s1[93], key_s0[93]}), .I1 ({new_AGEMA_signal_1144, \Midori/rounds_Output [29]}), .I2 ({key_s1[29], key_s0[29]}), .O ({output_1_s1[29], output_1_s0[29]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<28>1 ( .I0 ({key_s1[92], key_s0[92]}), .I1 ({new_AGEMA_signal_1143, \Midori/rounds_Output [28]}), .I2 ({key_s1[28], key_s0[28]}), .O ({output_1_s1[28], output_1_s0[28]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<27>1 ( .I0 ({key_s1[91], key_s0[91]}), .I1 ({new_AGEMA_signal_1138, \Midori/rounds_Output [27]}), .I2 ({key_s1[27], key_s0[27]}), .O ({output_1_s1[27], output_1_s0[27]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<26>1 ( .I0 ({key_s1[90], key_s0[90]}), .I1 ({new_AGEMA_signal_1137, \Midori/rounds_Output [26]}), .I2 ({key_s1[26], key_s0[26]}), .O ({output_1_s1[26], output_1_s0[26]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<25>1 ( .I0 ({new_AGEMA_signal_1136, \Midori/rounds_Output [25]}), .I1 ({key_s1[25], key_s0[25]}), .I2 ({key_s1[89], key_s0[89]}), .O ({output_1_s1[25], output_1_s0[25]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<24>1 ( .I0 ({new_AGEMA_signal_1135, \Midori/rounds_Output [24]}), .I1 ({key_s1[24], key_s0[24]}), .I2 ({key_s1[88], key_s0[88]}), .O ({output_1_s1[24], output_1_s0[24]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<23>1 ( .I0 ({new_AGEMA_signal_1130, \Midori/rounds_Output [23]}), .I1 ({key_s1[23], key_s0[23]}), .I2 ({key_s1[87], key_s0[87]}), .O ({output_1_s1[23], output_1_s0[23]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<22>1 ( .I0 ({new_AGEMA_signal_1129, \Midori/rounds_Output [22]}), .I1 ({key_s1[22], key_s0[22]}), .I2 ({key_s1[86], key_s0[86]}), .O ({output_1_s1[22], output_1_s0[22]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<21>1 ( .I0 ({new_AGEMA_signal_1128, \Midori/rounds_Output [21]}), .I1 ({key_s1[21], key_s0[21]}), .I2 ({key_s1[85], key_s0[85]}), .O ({output_1_s1[21], output_1_s0[21]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<20>1 ( .I0 ({new_AGEMA_signal_1127, \Midori/rounds_Output [20]}), .I1 ({key_s1[20], key_s0[20]}), .I2 ({key_s1[84], key_s0[84]}), .O ({output_1_s1[20], output_1_s0[20]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<2>1 ( .I0 ({new_AGEMA_signal_1089, \Midori/rounds_Output [2]}), .I1 ({key_s1[2], key_s0[2]}), .I2 ({key_s1[66], key_s0[66]}), .O ({output_1_s1[2], output_1_s0[2]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<19>1 ( .I0 ({key_s1[83], key_s0[83]}), .I1 ({new_AGEMA_signal_1122, \Midori/rounds_Output [19]}), .I2 ({key_s1[19], key_s0[19]}), .O ({output_1_s1[19], output_1_s0[19]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<18>1 ( .I0 ({key_s1[82], key_s0[82]}), .I1 ({new_AGEMA_signal_1121, \Midori/rounds_Output [18]}), .I2 ({key_s1[18], key_s0[18]}), .O ({output_1_s1[18], output_1_s0[18]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<17>1 ( .I0 ({key_s1[81], key_s0[81]}), .I1 ({new_AGEMA_signal_1120, \Midori/rounds_Output [17]}), .I2 ({key_s1[17], key_s0[17]}), .O ({output_1_s1[17], output_1_s0[17]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<16>1 ( .I0 ({key_s1[80], key_s0[80]}), .I1 ({new_AGEMA_signal_1119, \Midori/rounds_Output [16]}), .I2 ({key_s1[16], key_s0[16]}), .O ({output_1_s1[16], output_1_s0[16]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<15>1 ( .I0 ({new_AGEMA_signal_1114, \Midori/rounds_Output [15]}), .I1 ({key_s1[15], key_s0[15]}), .I2 ({key_s1[79], key_s0[79]}), .O ({output_1_s1[15], output_1_s0[15]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<14>1 ( .I0 ({new_AGEMA_signal_1113, \Midori/rounds_Output [14]}), .I1 ({key_s1[14], key_s0[14]}), .I2 ({key_s1[78], key_s0[78]}), .O ({output_1_s1[14], output_1_s0[14]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<13>1 ( .I0 ({new_AGEMA_signal_1112, \Midori/rounds_Output [13]}), .I1 ({key_s1[13], key_s0[13]}), .I2 ({key_s1[77], key_s0[77]}), .O ({output_1_s1[13], output_1_s0[13]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<12>1 ( .I0 ({new_AGEMA_signal_1111, \Midori/rounds_Output [12]}), .I1 ({key_s1[12], key_s0[12]}), .I2 ({key_s1[76], key_s0[76]}), .O ({output_1_s1[12], output_1_s0[12]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<11>1 ( .I0 ({new_AGEMA_signal_1106, \Midori/rounds_Output [11]}), .I1 ({key_s1[11], key_s0[11]}), .I2 ({key_s1[75], key_s0[75]}), .O ({output_1_s1[11], output_1_s0[11]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<10>1 ( .I0 ({new_AGEMA_signal_1105, \Midori/rounds_Output [10]}), .I1 ({key_s1[10], key_s0[10]}), .I2 ({key_s1[74], key_s0[74]}), .O ({output_1_s1[10], output_1_s0[10]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<1>1 ( .I0 ({new_AGEMA_signal_1088, \Midori/rounds_Output [1]}), .I1 ({key_s1[1], key_s0[1]}), .I2 ({key_s1[65], key_s0[65]}), .O ({output_1_s1[1], output_1_s0[1]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \output<0>1 ( .I0 ({new_AGEMA_signal_1087, \Midori/rounds_Output [0]}), .I1 ({key_s1[0], key_s0[0]}), .I2 ({key_s1[64], key_s0[64]}), .O ({output_1_s1[0], output_1_s0[0]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h4EE4 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h4EE4 ) ) \Midori/rounds/mul_input_Inst/gen_mux[56].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({new_AGEMA_signal_1127, \Midori/rounds_Output [20]}), .I2 ({new_AGEMA_signal_1199, \Midori/rounds_Output [56]}), .I3 ({new_AGEMA_signal_1676, \Midori/rounds/ProcessedKey [56]}), .O ({new_AGEMA_signal_1787, \Midori/rounds/mul_input [56]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h4EE4 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h4EE4 ) ) \Midori/rounds/mul_input_Inst/gen_mux[16].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({new_AGEMA_signal_1159, \Midori/rounds_Output [36]}), .I2 ({new_AGEMA_signal_1119, \Midori/rounds_Output [16]}), .I3 ({new_AGEMA_signal_1675, \Midori/rounds/ProcessedKey [16]}), .O ({new_AGEMA_signal_1788, \Midori/rounds/mul_input [16]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h4EE4 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h4EE4 ) ) \Midori/rounds/mul_input_Inst/gen_mux[0].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({new_AGEMA_signal_1143, \Midori/rounds_Output [28]}), .I2 ({new_AGEMA_signal_1087, \Midori/rounds_Output [0]}), .I3 ({new_AGEMA_signal_1674, \Midori/rounds/ProcessedKey [0]}), .O ({new_AGEMA_signal_1789, \Midori/rounds/mul_input [0]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hAFCF50305F3FA0C0 ) , .MASK ( 6'b101100 ), .INIT2 ( 64'h5F3FA0C05F3FA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[60].mux_inst/Mmux_Q11 ( .I0 ({key_s1[60], key_s0[60]}), .I1 ({key_s1[124], key_s0[124]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1207, \Midori/rounds_Output [60]}), .I5 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant15 }), .O ({new_AGEMA_signal_1613, \Midori/rounds/mul_input [60]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hAFCF50305F3FA0C0 ) , .MASK ( 6'b101100 ), .INIT2 ( 64'h5F3FA0C05F3FA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[8].mux_inst/Mmux_Q11 ( .I0 ({key_s1[8], key_s0[8]}), .I1 ({key_s1[72], key_s0[72]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1103, \Midori/rounds_Output [8]}), .I5 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant2 }), .O ({new_AGEMA_signal_1614, \Midori/rounds/mul_input [8]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h75FD20A8DF578A02 ) , .MASK ( 6'b000011 ), .INIT2 ( 64'h57DF028AFD75A820 ) ) \Midori/rounds/mul_input_Inst/gen_mux[48].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({1'b0, \controller/roundCounter/count [0]}), .I2 ({new_AGEMA_signal_1519, N111}), .I3 ({new_AGEMA_signal_1517, \Midori/rounds/Mxor_ProcessedKey<48>_xo<0> }), .I4 ({new_AGEMA_signal_1087, \Midori/rounds_Output [0]}), .I5 ({new_AGEMA_signal_1183, \Midori/rounds_Output [48]}), .O ({new_AGEMA_signal_1615, \Midori/rounds/mul_input [48]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h57DF028AFD75A820 ) , .MASK ( 6'b000011 ), .INIT2 ( 64'h57DF028AFD75A820 ) ) \Midori/rounds/mul_input_Inst/gen_mux[52].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({1'b0, \controller/roundCounter/count [0]}), .I2 ({new_AGEMA_signal_1516, \Midori/rounds/Mxor_ProcessedKey<52>_xo<0> }), .I3 ({new_AGEMA_signal_1520, N13}), .I4 ({new_AGEMA_signal_1167, \Midori/rounds_Output [40]}), .I5 ({new_AGEMA_signal_1191, \Midori/rounds_Output [52]}), .O ({new_AGEMA_signal_1616, \Midori/rounds/mul_input [52]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD87272D8 ) , .MASK ( 5'b10001 ), .INIT2 ( 32'h72D872D8 ) ) \Midori/rounds/mul_input_Inst/gen_mux[44].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({new_AGEMA_signal_1521, N15}), .I2 ({new_AGEMA_signal_1095, \Midori/rounds_Output [4]}), .I3 ({new_AGEMA_signal_1175, \Midori/rounds_Output [44]}), .I4 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant11 }), .O ({new_AGEMA_signal_1617, \Midori/rounds/mul_input [44]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h57DF028AFD75A820 ) , .MASK ( 6'b000011 ), .INIT2 ( 64'h57DF028AFD75A820 ) ) \Midori/rounds/mul_input_Inst/gen_mux[36].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({1'b0, \controller/roundCounter/count [0]}), .I2 ({new_AGEMA_signal_1515, \Midori/rounds/Mxor_ProcessedKey<36>_xo<0> }), .I3 ({new_AGEMA_signal_1522, N17}), .I4 ({new_AGEMA_signal_1119, \Midori/rounds_Output [16]}), .I5 ({new_AGEMA_signal_1159, \Midori/rounds_Output [36]}), .O ({new_AGEMA_signal_1618, \Midori/rounds/mul_input [36]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD87272D8 ) , .MASK ( 5'b10001 ), .INIT2 ( 32'h72D872D8 ) ) \Midori/rounds/mul_input_Inst/gen_mux[32].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({new_AGEMA_signal_1523, N19}), .I2 ({new_AGEMA_signal_1199, \Midori/rounds_Output [56]}), .I3 ({new_AGEMA_signal_1151, \Midori/rounds_Output [32]}), .I4 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant8 }), .O ({new_AGEMA_signal_1619, \Midori/rounds/mul_input [32]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD87272D8 ) , .MASK ( 5'b10001 ), .INIT2 ( 32'h72D872D8 ) ) \Midori/rounds/mul_input_Inst/gen_mux[28].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({new_AGEMA_signal_1524, N21}), .I2 ({new_AGEMA_signal_1135, \Midori/rounds_Output [24]}), .I3 ({new_AGEMA_signal_1143, \Midori/rounds_Output [28]}), .I4 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant7 }), .O ({new_AGEMA_signal_1620, \Midori/rounds/mul_input [28]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD87272D8 ) , .MASK ( 5'b10001 ), .INIT2 ( 32'h72D872D8 ) ) \Midori/rounds/mul_input_Inst/gen_mux[24].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({new_AGEMA_signal_1525, N23}), .I2 ({new_AGEMA_signal_1183, \Midori/rounds_Output [48]}), .I3 ({new_AGEMA_signal_1135, \Midori/rounds_Output [24]}), .I4 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant6 }), .O ({new_AGEMA_signal_1621, \Midori/rounds/mul_input [24]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD87272D8 ) , .MASK ( 5'b10001 ), .INIT2 ( 32'h72D872D8 ) ) \Midori/rounds/mul_input_Inst/gen_mux[20].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({new_AGEMA_signal_1526, N25}), .I2 ({new_AGEMA_signal_1111, \Midori/rounds_Output [12]}), .I3 ({new_AGEMA_signal_1127, \Midori/rounds_Output [20]}), .I4 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant5 }), .O ({new_AGEMA_signal_1622, \Midori/rounds/mul_input [20]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD87272D8 ) , .MASK ( 5'b10001 ), .INIT2 ( 32'h72D872D8 ) ) \Midori/rounds/mul_input_Inst/gen_mux[12].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({new_AGEMA_signal_1527, N27}), .I2 ({new_AGEMA_signal_1151, \Midori/rounds_Output [32]}), .I3 ({new_AGEMA_signal_1111, \Midori/rounds_Output [12]}), .I4 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant3 }), .O ({new_AGEMA_signal_1623, \Midori/rounds/mul_input [12]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD87272D8 ) , .MASK ( 5'b10001 ), .INIT2 ( 32'h72D872D8 ) ) \Midori/rounds/mul_input_Inst/gen_mux[4].mux_inst/Mmux_Q11 ( .I0 ({1'b0, enc_dec}), .I1 ({new_AGEMA_signal_1528, N29}), .I2 ({new_AGEMA_signal_1191, \Midori/rounds_Output [52]}), .I3 ({new_AGEMA_signal_1095, \Midori/rounds_Output [4]}), .I4 ({1'b0, \Midori/rounds/constant_MUX/Mram_roundConstant1 }), .O ({new_AGEMA_signal_1624, \Midori/rounds/mul_input [4]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h7F734C40B3BF808C ) , .MASK ( 6'b000110 ), .INIT2 ( 64'h737F404CBFB38C80 ) ) \Midori/rounds/mul_input_Inst/gen_mux[40].mux_inst/Mmux_Q11 ( .I0 ({key_s1[40], key_s0[40]}), .I1 ({1'b0, enc_dec}), .I2 ({1'b0, \controller/roundCounter/count [0]}), .I3 ({new_AGEMA_signal_1529, N34}), .I4 ({new_AGEMA_signal_1175, \Midori/rounds_Output [44]}), .I5 ({new_AGEMA_signal_1167, \Midori/rounds_Output [40]}), .O ({new_AGEMA_signal_1625, \Midori/rounds/mul_input [40]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h5F3FA0C0 ) , .MASK ( 5'b01100 ), .INIT2 ( 32'h5F3FA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[63].mux_inst/Mmux_Q11 ( .I0 ({key_s1[63], key_s0[63]}), .I1 ({key_s1[127], key_s0[127]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1210, \Midori/rounds_Output [63]}), .O ({new_AGEMA_signal_1626, \Midori/rounds/mul_input [63]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h5F3FA0C0 ) , .MASK ( 5'b01100 ), .INIT2 ( 32'h5F3FA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[62].mux_inst/Mmux_Q11 ( .I0 ({key_s1[62], key_s0[62]}), .I1 ({key_s1[126], key_s0[126]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1209, \Midori/rounds_Output [62]}), .O ({new_AGEMA_signal_1627, \Midori/rounds/mul_input [62]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h5F3FA0C0 ) , .MASK ( 5'b01100 ), .INIT2 ( 32'h5F3FA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[61].mux_inst/Mmux_Q11 ( .I0 ({key_s1[61], key_s0[61]}), .I1 ({key_s1[125], key_s0[125]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1208, \Midori/rounds_Output [61]}), .O ({new_AGEMA_signal_1628, \Midori/rounds/mul_input [61]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h5F3FA0C0 ) , .MASK ( 5'b01100 ), .INIT2 ( 32'h5F3FA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[11].mux_inst/Mmux_Q11 ( .I0 ({key_s1[11], key_s0[11]}), .I1 ({key_s1[75], key_s0[75]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1106, \Midori/rounds_Output [11]}), .O ({new_AGEMA_signal_1629, \Midori/rounds/mul_input [11]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h5F3FA0C0 ) , .MASK ( 5'b01100 ), .INIT2 ( 32'h5F3FA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[10].mux_inst/Mmux_Q11 ( .I0 ({key_s1[10], key_s0[10]}), .I1 ({key_s1[74], key_s0[74]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1105, \Midori/rounds_Output [10]}), .O ({new_AGEMA_signal_1630, \Midori/rounds/mul_input [10]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h5F3FA0C0 ) , .MASK ( 5'b01100 ), .INIT2 ( 32'h5F3FA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[9].mux_inst/Mmux_Q11 ( .I0 ({key_s1[9], key_s0[9]}), .I1 ({key_s1[73], key_s0[73]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1104, \Midori/rounds_Output [9]}), .O ({new_AGEMA_signal_1631, \Midori/rounds/mul_input [9]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[59].mux_inst/Mmux_Q11 ( .I0 ({key_s1[59], key_s0[59]}), .I1 ({key_s1[123], key_s0[123]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1130, \Midori/rounds_Output [23]}), .I5 ({new_AGEMA_signal_1202, \Midori/rounds_Output [59]}), .O ({new_AGEMA_signal_1632, \Midori/rounds/mul_input [59]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[58].mux_inst/Mmux_Q11 ( .I0 ({key_s1[58], key_s0[58]}), .I1 ({key_s1[122], key_s0[122]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1129, \Midori/rounds_Output [22]}), .I5 ({new_AGEMA_signal_1201, \Midori/rounds_Output [58]}), .O ({new_AGEMA_signal_1633, \Midori/rounds/mul_input [58]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[57].mux_inst/Mmux_Q11 ( .I0 ({key_s1[57], key_s0[57]}), .I1 ({key_s1[121], key_s0[121]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1128, \Midori/rounds_Output [21]}), .I5 ({new_AGEMA_signal_1200, \Midori/rounds_Output [57]}), .O ({new_AGEMA_signal_1634, \Midori/rounds/mul_input [57]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[55].mux_inst/Mmux_Q11 ( .I0 ({key_s1[55], key_s0[55]}), .I1 ({key_s1[119], key_s0[119]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1170, \Midori/rounds_Output [43]}), .I5 ({new_AGEMA_signal_1194, \Midori/rounds_Output [55]}), .O ({new_AGEMA_signal_1635, \Midori/rounds/mul_input [55]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[54].mux_inst/Mmux_Q11 ( .I0 ({key_s1[54], key_s0[54]}), .I1 ({key_s1[118], key_s0[118]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1169, \Midori/rounds_Output [42]}), .I5 ({new_AGEMA_signal_1193, \Midori/rounds_Output [54]}), .O ({new_AGEMA_signal_1636, \Midori/rounds/mul_input [54]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[53].mux_inst/Mmux_Q11 ( .I0 ({key_s1[53], key_s0[53]}), .I1 ({key_s1[117], key_s0[117]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1168, \Midori/rounds_Output [41]}), .I5 ({new_AGEMA_signal_1192, \Midori/rounds_Output [53]}), .O ({new_AGEMA_signal_1637, \Midori/rounds/mul_input [53]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[51].mux_inst/Mmux_Q11 ( .I0 ({key_s1[51], key_s0[51]}), .I1 ({key_s1[115], key_s0[115]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1090, \Midori/rounds_Output [3]}), .I5 ({new_AGEMA_signal_1186, \Midori/rounds_Output [51]}), .O ({new_AGEMA_signal_1638, \Midori/rounds/mul_input [51]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[50].mux_inst/Mmux_Q11 ( .I0 ({key_s1[50], key_s0[50]}), .I1 ({key_s1[114], key_s0[114]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1089, \Midori/rounds_Output [2]}), .I5 ({new_AGEMA_signal_1185, \Midori/rounds_Output [50]}), .O ({new_AGEMA_signal_1639, \Midori/rounds/mul_input [50]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[49].mux_inst/Mmux_Q11 ( .I0 ({key_s1[49], key_s0[49]}), .I1 ({key_s1[113], key_s0[113]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1088, \Midori/rounds_Output [1]}), .I5 ({new_AGEMA_signal_1184, \Midori/rounds_Output [49]}), .O ({new_AGEMA_signal_1640, \Midori/rounds/mul_input [49]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[47].mux_inst/Mmux_Q11 ( .I0 ({key_s1[47], key_s0[47]}), .I1 ({key_s1[111], key_s0[111]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1098, \Midori/rounds_Output [7]}), .I5 ({new_AGEMA_signal_1178, \Midori/rounds_Output [47]}), .O ({new_AGEMA_signal_1641, \Midori/rounds/mul_input [47]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[46].mux_inst/Mmux_Q11 ( .I0 ({key_s1[46], key_s0[46]}), .I1 ({key_s1[110], key_s0[110]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1097, \Midori/rounds_Output [6]}), .I5 ({new_AGEMA_signal_1177, \Midori/rounds_Output [46]}), .O ({new_AGEMA_signal_1642, \Midori/rounds/mul_input [46]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[45].mux_inst/Mmux_Q11 ( .I0 ({key_s1[45], key_s0[45]}), .I1 ({key_s1[109], key_s0[109]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1096, \Midori/rounds_Output [5]}), .I5 ({new_AGEMA_signal_1176, \Midori/rounds_Output [45]}), .O ({new_AGEMA_signal_1643, \Midori/rounds/mul_input [45]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[43].mux_inst/Mmux_Q11 ( .I0 ({key_s1[43], key_s0[43]}), .I1 ({key_s1[107], key_s0[107]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1178, \Midori/rounds_Output [47]}), .I5 ({new_AGEMA_signal_1170, \Midori/rounds_Output [43]}), .O ({new_AGEMA_signal_1644, \Midori/rounds/mul_input [43]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[42].mux_inst/Mmux_Q11 ( .I0 ({key_s1[42], key_s0[42]}), .I1 ({key_s1[106], key_s0[106]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1177, \Midori/rounds_Output [46]}), .I5 ({new_AGEMA_signal_1169, \Midori/rounds_Output [42]}), .O ({new_AGEMA_signal_1645, \Midori/rounds/mul_input [42]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[41].mux_inst/Mmux_Q11 ( .I0 ({key_s1[41], key_s0[41]}), .I1 ({key_s1[105], key_s0[105]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1176, \Midori/rounds_Output [45]}), .I5 ({new_AGEMA_signal_1168, \Midori/rounds_Output [41]}), .O ({new_AGEMA_signal_1646, \Midori/rounds/mul_input [41]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[39].mux_inst/Mmux_Q11 ( .I0 ({key_s1[39], key_s0[39]}), .I1 ({key_s1[103], key_s0[103]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1122, \Midori/rounds_Output [19]}), .I5 ({new_AGEMA_signal_1162, \Midori/rounds_Output [39]}), .O ({new_AGEMA_signal_1647, \Midori/rounds/mul_input [39]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[38].mux_inst/Mmux_Q11 ( .I0 ({key_s1[38], key_s0[38]}), .I1 ({key_s1[102], key_s0[102]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1121, \Midori/rounds_Output [18]}), .I5 ({new_AGEMA_signal_1161, \Midori/rounds_Output [38]}), .O ({new_AGEMA_signal_1648, \Midori/rounds/mul_input [38]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[37].mux_inst/Mmux_Q11 ( .I0 ({key_s1[37], key_s0[37]}), .I1 ({key_s1[101], key_s0[101]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1120, \Midori/rounds_Output [17]}), .I5 ({new_AGEMA_signal_1160, \Midori/rounds_Output [37]}), .O ({new_AGEMA_signal_1649, \Midori/rounds/mul_input [37]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[35].mux_inst/Mmux_Q11 ( .I0 ({key_s1[35], key_s0[35]}), .I1 ({key_s1[99], key_s0[99]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1202, \Midori/rounds_Output [59]}), .I5 ({new_AGEMA_signal_1154, \Midori/rounds_Output [35]}), .O ({new_AGEMA_signal_1650, \Midori/rounds/mul_input [35]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[34].mux_inst/Mmux_Q11 ( .I0 ({key_s1[34], key_s0[34]}), .I1 ({key_s1[98], key_s0[98]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1201, \Midori/rounds_Output [58]}), .I5 ({new_AGEMA_signal_1153, \Midori/rounds_Output [34]}), .O ({new_AGEMA_signal_1651, \Midori/rounds/mul_input [34]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[33].mux_inst/Mmux_Q11 ( .I0 ({key_s1[33], key_s0[33]}), .I1 ({key_s1[97], key_s0[97]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1200, \Midori/rounds_Output [57]}), .I5 ({new_AGEMA_signal_1152, \Midori/rounds_Output [33]}), .O ({new_AGEMA_signal_1652, \Midori/rounds/mul_input [33]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[31].mux_inst/Mmux_Q11 ( .I0 ({key_s1[31], key_s0[31]}), .I1 ({key_s1[95], key_s0[95]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1138, \Midori/rounds_Output [27]}), .I5 ({new_AGEMA_signal_1146, \Midori/rounds_Output [31]}), .O ({new_AGEMA_signal_1653, \Midori/rounds/mul_input [31]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[30].mux_inst/Mmux_Q11 ( .I0 ({key_s1[30], key_s0[30]}), .I1 ({key_s1[94], key_s0[94]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1137, \Midori/rounds_Output [26]}), .I5 ({new_AGEMA_signal_1145, \Midori/rounds_Output [30]}), .O ({new_AGEMA_signal_1654, \Midori/rounds/mul_input [30]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[29].mux_inst/Mmux_Q11 ( .I0 ({key_s1[29], key_s0[29]}), .I1 ({key_s1[93], key_s0[93]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1136, \Midori/rounds_Output [25]}), .I5 ({new_AGEMA_signal_1144, \Midori/rounds_Output [29]}), .O ({new_AGEMA_signal_1655, \Midori/rounds/mul_input [29]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[27].mux_inst/Mmux_Q11 ( .I0 ({key_s1[27], key_s0[27]}), .I1 ({key_s1[91], key_s0[91]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1186, \Midori/rounds_Output [51]}), .I5 ({new_AGEMA_signal_1138, \Midori/rounds_Output [27]}), .O ({new_AGEMA_signal_1656, \Midori/rounds/mul_input [27]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[26].mux_inst/Mmux_Q11 ( .I0 ({key_s1[26], key_s0[26]}), .I1 ({key_s1[90], key_s0[90]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1185, \Midori/rounds_Output [50]}), .I5 ({new_AGEMA_signal_1137, \Midori/rounds_Output [26]}), .O ({new_AGEMA_signal_1657, \Midori/rounds/mul_input [26]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[25].mux_inst/Mmux_Q11 ( .I0 ({key_s1[25], key_s0[25]}), .I1 ({key_s1[89], key_s0[89]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1184, \Midori/rounds_Output [49]}), .I5 ({new_AGEMA_signal_1136, \Midori/rounds_Output [25]}), .O ({new_AGEMA_signal_1658, \Midori/rounds/mul_input [25]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[23].mux_inst/Mmux_Q11 ( .I0 ({key_s1[23], key_s0[23]}), .I1 ({key_s1[87], key_s0[87]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1114, \Midori/rounds_Output [15]}), .I5 ({new_AGEMA_signal_1130, \Midori/rounds_Output [23]}), .O ({new_AGEMA_signal_1659, \Midori/rounds/mul_input [23]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[22].mux_inst/Mmux_Q11 ( .I0 ({key_s1[22], key_s0[22]}), .I1 ({key_s1[86], key_s0[86]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1113, \Midori/rounds_Output [14]}), .I5 ({new_AGEMA_signal_1129, \Midori/rounds_Output [22]}), .O ({new_AGEMA_signal_1660, \Midori/rounds/mul_input [22]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[21].mux_inst/Mmux_Q11 ( .I0 ({key_s1[21], key_s0[21]}), .I1 ({key_s1[85], key_s0[85]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1112, \Midori/rounds_Output [13]}), .I5 ({new_AGEMA_signal_1128, \Midori/rounds_Output [21]}), .O ({new_AGEMA_signal_1661, \Midori/rounds/mul_input [21]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[19].mux_inst/Mmux_Q11 ( .I0 ({key_s1[19], key_s0[19]}), .I1 ({key_s1[83], key_s0[83]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1162, \Midori/rounds_Output [39]}), .I5 ({new_AGEMA_signal_1122, \Midori/rounds_Output [19]}), .O ({new_AGEMA_signal_1662, \Midori/rounds/mul_input [19]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[18].mux_inst/Mmux_Q11 ( .I0 ({key_s1[18], key_s0[18]}), .I1 ({key_s1[82], key_s0[82]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1161, \Midori/rounds_Output [38]}), .I5 ({new_AGEMA_signal_1121, \Midori/rounds_Output [18]}), .O ({new_AGEMA_signal_1663, \Midori/rounds/mul_input [18]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[17].mux_inst/Mmux_Q11 ( .I0 ({key_s1[17], key_s0[17]}), .I1 ({key_s1[81], key_s0[81]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1160, \Midori/rounds_Output [37]}), .I5 ({new_AGEMA_signal_1120, \Midori/rounds_Output [17]}), .O ({new_AGEMA_signal_1664, \Midori/rounds/mul_input [17]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[15].mux_inst/Mmux_Q11 ( .I0 ({key_s1[15], key_s0[15]}), .I1 ({key_s1[79], key_s0[79]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1154, \Midori/rounds_Output [35]}), .I5 ({new_AGEMA_signal_1114, \Midori/rounds_Output [15]}), .O ({new_AGEMA_signal_1665, \Midori/rounds/mul_input [15]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[14].mux_inst/Mmux_Q11 ( .I0 ({key_s1[14], key_s0[14]}), .I1 ({key_s1[78], key_s0[78]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1153, \Midori/rounds_Output [34]}), .I5 ({new_AGEMA_signal_1113, \Midori/rounds_Output [14]}), .O ({new_AGEMA_signal_1666, \Midori/rounds/mul_input [14]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[13].mux_inst/Mmux_Q11 ( .I0 ({key_s1[13], key_s0[13]}), .I1 ({key_s1[77], key_s0[77]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1152, \Midori/rounds_Output [33]}), .I5 ({new_AGEMA_signal_1112, \Midori/rounds_Output [13]}), .O ({new_AGEMA_signal_1667, \Midori/rounds/mul_input [13]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[7].mux_inst/Mmux_Q11 ( .I0 ({key_s1[7], key_s0[7]}), .I1 ({key_s1[71], key_s0[71]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1194, \Midori/rounds_Output [55]}), .I5 ({new_AGEMA_signal_1098, \Midori/rounds_Output [7]}), .O ({new_AGEMA_signal_1668, \Midori/rounds/mul_input [7]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[6].mux_inst/Mmux_Q11 ( .I0 ({key_s1[6], key_s0[6]}), .I1 ({key_s1[70], key_s0[70]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1193, \Midori/rounds_Output [54]}), .I5 ({new_AGEMA_signal_1097, \Midori/rounds_Output [6]}), .O ({new_AGEMA_signal_1669, \Midori/rounds/mul_input [6]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[5].mux_inst/Mmux_Q11 ( .I0 ({key_s1[5], key_s0[5]}), .I1 ({key_s1[69], key_s0[69]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1192, \Midori/rounds_Output [53]}), .I5 ({new_AGEMA_signal_1096, \Midori/rounds_Output [5]}), .O ({new_AGEMA_signal_1670, \Midori/rounds/mul_input [5]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[3].mux_inst/Mmux_Q11 ( .I0 ({key_s1[3], key_s0[3]}), .I1 ({key_s1[67], key_s0[67]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1146, \Midori/rounds_Output [31]}), .I5 ({new_AGEMA_signal_1090, \Midori/rounds_Output [3]}), .O ({new_AGEMA_signal_1671, \Midori/rounds/mul_input [3]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[2].mux_inst/Mmux_Q11 ( .I0 ({key_s1[2], key_s0[2]}), .I1 ({key_s1[66], key_s0[66]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1145, \Midori/rounds_Output [30]}), .I5 ({new_AGEMA_signal_1089, \Midori/rounds_Output [2]}), .O ({new_AGEMA_signal_1672, \Midori/rounds/mul_input [2]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5F3F5030AFCFA0C0 ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h5F3F5030AFCFA0C0 ) ) \Midori/rounds/mul_input_Inst/gen_mux[1].mux_inst/Mmux_Q11 ( .I0 ({key_s1[1], key_s0[1]}), .I1 ({key_s1[65], key_s0[65]}), .I2 ({1'b0, enc_dec}), .I3 ({1'b0, \controller/roundCounter/count [0]}), .I4 ({new_AGEMA_signal_1144, \Midori/rounds_Output [29]}), .I5 ({new_AGEMA_signal_1088, \Midori/rounds_Output [1]}), .O ({new_AGEMA_signal_1673, \Midori/rounds/mul_input [1]}) ) ;

    /* register cells */
    FDR \controller/roundCounter/count_0 ( .D (Result[0]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count [0]) ) ;
    FDR \controller/roundCounter/count_1 ( .D (Result[1]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count [1]) ) ;
    FDR \controller/roundCounter/count_2 ( .D (Result[2]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count [2]) ) ;
    FDR \controller/roundCounter/count_3 ( .D (Result[3]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count [3]) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1860, \Midori/rounds/roundResult_Reg/GEN[0].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1083, \Midori/rounds/roundResult_Reg/GEN[0].SFF/Q_663 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1790, \Midori/rounds/roundResult_Reg/GEN[1].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1084, \Midori/rounds/roundResult_Reg/GEN[1].SFF/Q_664 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1791, \Midori/rounds/roundResult_Reg/GEN[2].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1085, \Midori/rounds/roundResult_Reg/GEN[2].SFF/Q_665 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1792, \Midori/rounds/roundResult_Reg/GEN[3].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1086, \Midori/rounds/roundResult_Reg/GEN[3].SFF/Q_666 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1861, \Midori/rounds/roundResult_Reg/GEN[4].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1091, \Midori/rounds/roundResult_Reg/GEN[4].SFF/Q_667 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1793, \Midori/rounds/roundResult_Reg/GEN[5].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1092, \Midori/rounds/roundResult_Reg/GEN[5].SFF/Q_668 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1794, \Midori/rounds/roundResult_Reg/GEN[6].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1093, \Midori/rounds/roundResult_Reg/GEN[6].SFF/Q_669 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1795, \Midori/rounds/roundResult_Reg/GEN[7].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1094, \Midori/rounds/roundResult_Reg/GEN[7].SFF/Q_670 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[8].SFF/Q ( .D ({new_AGEMA_signal_1862, \Midori/rounds/roundResult_Reg/GEN[8].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1099, \Midori/rounds/roundResult_Reg/GEN[8].SFF/Q_671 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[9].SFF/Q ( .D ({new_AGEMA_signal_1796, \Midori/rounds/roundResult_Reg/GEN[9].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1100, \Midori/rounds/roundResult_Reg/GEN[9].SFF/Q_672 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[10].SFF/Q ( .D ({new_AGEMA_signal_1797, \Midori/rounds/roundResult_Reg/GEN[10].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1101, \Midori/rounds/roundResult_Reg/GEN[10].SFF/Q_673 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[11].SFF/Q ( .D ({new_AGEMA_signal_1798, \Midori/rounds/roundResult_Reg/GEN[11].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1102, \Midori/rounds/roundResult_Reg/GEN[11].SFF/Q_674 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[12].SFF/Q ( .D ({new_AGEMA_signal_1863, \Midori/rounds/roundResult_Reg/GEN[12].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1107, \Midori/rounds/roundResult_Reg/GEN[12].SFF/Q_675 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[13].SFF/Q ( .D ({new_AGEMA_signal_1799, \Midori/rounds/roundResult_Reg/GEN[13].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1108, \Midori/rounds/roundResult_Reg/GEN[13].SFF/Q_676 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[14].SFF/Q ( .D ({new_AGEMA_signal_1800, \Midori/rounds/roundResult_Reg/GEN[14].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1109, \Midori/rounds/roundResult_Reg/GEN[14].SFF/Q_677 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[15].SFF/Q ( .D ({new_AGEMA_signal_1801, \Midori/rounds/roundResult_Reg/GEN[15].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1110, \Midori/rounds/roundResult_Reg/GEN[15].SFF/Q_678 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[16].SFF/Q ( .D ({new_AGEMA_signal_1802, \Midori/rounds/roundResult_Reg/GEN[16].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1115, \Midori/rounds/roundResult_Reg/GEN[16].SFF/Q_679 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[17].SFF/Q ( .D ({new_AGEMA_signal_1803, \Midori/rounds/roundResult_Reg/GEN[17].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1116, \Midori/rounds/roundResult_Reg/GEN[17].SFF/Q_680 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[18].SFF/Q ( .D ({new_AGEMA_signal_1804, \Midori/rounds/roundResult_Reg/GEN[18].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1117, \Midori/rounds/roundResult_Reg/GEN[18].SFF/Q_681 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[19].SFF/Q ( .D ({new_AGEMA_signal_1805, \Midori/rounds/roundResult_Reg/GEN[19].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1118, \Midori/rounds/roundResult_Reg/GEN[19].SFF/Q_682 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[20].SFF/Q ( .D ({new_AGEMA_signal_1864, \Midori/rounds/roundResult_Reg/GEN[20].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1123, \Midori/rounds/roundResult_Reg/GEN[20].SFF/Q_683 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[21].SFF/Q ( .D ({new_AGEMA_signal_1806, \Midori/rounds/roundResult_Reg/GEN[21].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1124, \Midori/rounds/roundResult_Reg/GEN[21].SFF/Q_684 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[22].SFF/Q ( .D ({new_AGEMA_signal_1807, \Midori/rounds/roundResult_Reg/GEN[22].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1125, \Midori/rounds/roundResult_Reg/GEN[22].SFF/Q_685 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[23].SFF/Q ( .D ({new_AGEMA_signal_1808, \Midori/rounds/roundResult_Reg/GEN[23].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1126, \Midori/rounds/roundResult_Reg/GEN[23].SFF/Q_686 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[24].SFF/Q ( .D ({new_AGEMA_signal_1865, \Midori/rounds/roundResult_Reg/GEN[24].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1131, \Midori/rounds/roundResult_Reg/GEN[24].SFF/Q_687 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[25].SFF/Q ( .D ({new_AGEMA_signal_1809, \Midori/rounds/roundResult_Reg/GEN[25].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1132, \Midori/rounds/roundResult_Reg/GEN[25].SFF/Q_688 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[26].SFF/Q ( .D ({new_AGEMA_signal_1810, \Midori/rounds/roundResult_Reg/GEN[26].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1133, \Midori/rounds/roundResult_Reg/GEN[26].SFF/Q_689 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[27].SFF/Q ( .D ({new_AGEMA_signal_1811, \Midori/rounds/roundResult_Reg/GEN[27].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1134, \Midori/rounds/roundResult_Reg/GEN[27].SFF/Q_690 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[28].SFF/Q ( .D ({new_AGEMA_signal_1866, \Midori/rounds/roundResult_Reg/GEN[28].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1139, \Midori/rounds/roundResult_Reg/GEN[28].SFF/Q_691 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[29].SFF/Q ( .D ({new_AGEMA_signal_1812, \Midori/rounds/roundResult_Reg/GEN[29].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1140, \Midori/rounds/roundResult_Reg/GEN[29].SFF/Q_692 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[30].SFF/Q ( .D ({new_AGEMA_signal_1813, \Midori/rounds/roundResult_Reg/GEN[30].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1141, \Midori/rounds/roundResult_Reg/GEN[30].SFF/Q_693 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[31].SFF/Q ( .D ({new_AGEMA_signal_1814, \Midori/rounds/roundResult_Reg/GEN[31].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1142, \Midori/rounds/roundResult_Reg/GEN[31].SFF/Q_694 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[32].SFF/Q ( .D ({new_AGEMA_signal_1867, \Midori/rounds/roundResult_Reg/GEN[32].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1147, \Midori/rounds/roundResult_Reg/GEN[32].SFF/Q_695 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[33].SFF/Q ( .D ({new_AGEMA_signal_1815, \Midori/rounds/roundResult_Reg/GEN[33].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1148, \Midori/rounds/roundResult_Reg/GEN[33].SFF/Q_696 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[34].SFF/Q ( .D ({new_AGEMA_signal_1816, \Midori/rounds/roundResult_Reg/GEN[34].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1149, \Midori/rounds/roundResult_Reg/GEN[34].SFF/Q_697 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[35].SFF/Q ( .D ({new_AGEMA_signal_1817, \Midori/rounds/roundResult_Reg/GEN[35].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1150, \Midori/rounds/roundResult_Reg/GEN[35].SFF/Q_698 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[36].SFF/Q ( .D ({new_AGEMA_signal_1818, \Midori/rounds/roundResult_Reg/GEN[36].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1155, \Midori/rounds/roundResult_Reg/GEN[36].SFF/Q_699 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[37].SFF/Q ( .D ({new_AGEMA_signal_1819, \Midori/rounds/roundResult_Reg/GEN[37].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1156, \Midori/rounds/roundResult_Reg/GEN[37].SFF/Q_700 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[38].SFF/Q ( .D ({new_AGEMA_signal_1820, \Midori/rounds/roundResult_Reg/GEN[38].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1157, \Midori/rounds/roundResult_Reg/GEN[38].SFF/Q_701 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[39].SFF/Q ( .D ({new_AGEMA_signal_1821, \Midori/rounds/roundResult_Reg/GEN[39].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1158, \Midori/rounds/roundResult_Reg/GEN[39].SFF/Q_702 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[40].SFF/Q ( .D ({new_AGEMA_signal_1868, \Midori/rounds/roundResult_Reg/GEN[40].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1163, \Midori/rounds/roundResult_Reg/GEN[40].SFF/Q_703 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[41].SFF/Q ( .D ({new_AGEMA_signal_1822, \Midori/rounds/roundResult_Reg/GEN[41].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1164, \Midori/rounds/roundResult_Reg/GEN[41].SFF/Q_704 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[42].SFF/Q ( .D ({new_AGEMA_signal_1823, \Midori/rounds/roundResult_Reg/GEN[42].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1165, \Midori/rounds/roundResult_Reg/GEN[42].SFF/Q_705 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[43].SFF/Q ( .D ({new_AGEMA_signal_1824, \Midori/rounds/roundResult_Reg/GEN[43].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1166, \Midori/rounds/roundResult_Reg/GEN[43].SFF/Q_706 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[44].SFF/Q ( .D ({new_AGEMA_signal_1825, \Midori/rounds/roundResult_Reg/GEN[44].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1171, \Midori/rounds/roundResult_Reg/GEN[44].SFF/Q_707 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[45].SFF/Q ( .D ({new_AGEMA_signal_1826, \Midori/rounds/roundResult_Reg/GEN[45].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1172, \Midori/rounds/roundResult_Reg/GEN[45].SFF/Q_708 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[46].SFF/Q ( .D ({new_AGEMA_signal_1827, \Midori/rounds/roundResult_Reg/GEN[46].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1173, \Midori/rounds/roundResult_Reg/GEN[46].SFF/Q_709 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[47].SFF/Q ( .D ({new_AGEMA_signal_1828, \Midori/rounds/roundResult_Reg/GEN[47].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1174, \Midori/rounds/roundResult_Reg/GEN[47].SFF/Q_710 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[48].SFF/Q ( .D ({new_AGEMA_signal_1869, \Midori/rounds/roundResult_Reg/GEN[48].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1179, \Midori/rounds/roundResult_Reg/GEN[48].SFF/Q_711 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[49].SFF/Q ( .D ({new_AGEMA_signal_1829, \Midori/rounds/roundResult_Reg/GEN[49].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1180, \Midori/rounds/roundResult_Reg/GEN[49].SFF/Q_712 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[50].SFF/Q ( .D ({new_AGEMA_signal_1830, \Midori/rounds/roundResult_Reg/GEN[50].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1181, \Midori/rounds/roundResult_Reg/GEN[50].SFF/Q_713 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[51].SFF/Q ( .D ({new_AGEMA_signal_1831, \Midori/rounds/roundResult_Reg/GEN[51].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1182, \Midori/rounds/roundResult_Reg/GEN[51].SFF/Q_714 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[52].SFF/Q ( .D ({new_AGEMA_signal_1870, \Midori/rounds/roundResult_Reg/GEN[52].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1187, \Midori/rounds/roundResult_Reg/GEN[52].SFF/Q_715 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[53].SFF/Q ( .D ({new_AGEMA_signal_1832, \Midori/rounds/roundResult_Reg/GEN[53].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1188, \Midori/rounds/roundResult_Reg/GEN[53].SFF/Q_716 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[54].SFF/Q ( .D ({new_AGEMA_signal_1833, \Midori/rounds/roundResult_Reg/GEN[54].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1189, \Midori/rounds/roundResult_Reg/GEN[54].SFF/Q_717 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[55].SFF/Q ( .D ({new_AGEMA_signal_1834, \Midori/rounds/roundResult_Reg/GEN[55].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1190, \Midori/rounds/roundResult_Reg/GEN[55].SFF/Q_718 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[56].SFF/Q ( .D ({new_AGEMA_signal_1835, \Midori/rounds/roundResult_Reg/GEN[56].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1195, \Midori/rounds/roundResult_Reg/GEN[56].SFF/Q_719 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[57].SFF/Q ( .D ({new_AGEMA_signal_1836, \Midori/rounds/roundResult_Reg/GEN[57].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1196, \Midori/rounds/roundResult_Reg/GEN[57].SFF/Q_720 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[58].SFF/Q ( .D ({new_AGEMA_signal_1837, \Midori/rounds/roundResult_Reg/GEN[58].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1197, \Midori/rounds/roundResult_Reg/GEN[58].SFF/Q_721 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[59].SFF/Q ( .D ({new_AGEMA_signal_1838, \Midori/rounds/roundResult_Reg/GEN[59].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1198, \Midori/rounds/roundResult_Reg/GEN[59].SFF/Q_722 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[60].SFF/Q ( .D ({new_AGEMA_signal_1871, \Midori/rounds/roundResult_Reg/GEN[60].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1203, \Midori/rounds/roundResult_Reg/GEN[60].SFF/Q_723 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[61].SFF/Q ( .D ({new_AGEMA_signal_1839, \Midori/rounds/roundResult_Reg/GEN[61].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1204, \Midori/rounds/roundResult_Reg/GEN[61].SFF/Q_724 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[62].SFF/Q ( .D ({new_AGEMA_signal_1840, \Midori/rounds/roundResult_Reg/GEN[62].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1205, \Midori/rounds/roundResult_Reg/GEN[62].SFF/Q_725 }) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \Midori/rounds/roundResult_Reg/GEN[63].SFF/Q ( .D ({new_AGEMA_signal_1841, \Midori/rounds/roundResult_Reg/GEN[63].SFF/DQ }), .clk (clk_gated), .Q ({new_AGEMA_signal_1206, \Midori/rounds/roundResult_Reg/GEN[63].SFF/Q_726 }) ) ;
    FDR \controller/roundCounter/count_3_1 ( .D (Result[3]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count_3_1_1066 ) ) ;
    FDR \controller/roundCounter/count_2_1 ( .D (Result[2]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count_2_1_1067 ) ) ;
    FDR \controller/roundCounter/count_0_1 ( .D (Result[0]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count_0_1_1068 ) ) ;
    FDR \controller/roundCounter/count_1_1 ( .D (Result[1]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count_1_1_1069 ) ) ;
    FDR \controller/roundCounter/count_2_2 ( .D (Result[2]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count_2_2_1070 ) ) ;
    FDR \controller/roundCounter/count_3_2 ( .D (Result[3]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count_3_2_1071 ) ) ;
    FDR \controller/roundCounter/count_1_2 ( .D (Result[1]), .C (clk_gated), .R (reset), .Q (\controller/roundCounter/count_1_2_1072 ) ) ;
endmodule
